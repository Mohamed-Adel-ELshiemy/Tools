
module instr_mem ( pc, instruction );
  input [15:0] pc;
  output [15:0] instruction;

  assign instruction[0] = 1'b0;
  assign instruction[1] = 1'b0;
  assign instruction[2] = 1'b0;
  assign instruction[3] = 1'b0;
  assign instruction[4] = 1'b0;
  assign instruction[5] = 1'b0;
  assign instruction[6] = 1'b0;
  assign instruction[7] = 1'b0;
  assign instruction[8] = 1'b0;
  assign instruction[9] = 1'b0;
  assign instruction[10] = 1'b0;
  assign instruction[11] = 1'b0;
  assign instruction[12] = 1'b0;
  assign instruction[13] = 1'b0;
  assign instruction[14] = 1'b0;
  assign instruction[15] = 1'b0;

endmodule


module control ( opcode, reset, reg_dst, mem_to_reg, alu_op, jump, branch, 
        mem_read, mem_write, alu_src, reg_write, sign_or_zero );
  input [2:0] opcode;
  output [1:0] reg_dst;
  output [1:0] mem_to_reg;
  output [1:0] alu_op;
  input reset;
  output jump, branch, mem_read, mem_write, alu_src, reg_write, sign_or_zero;
  wire   n7, n8, n9, n10, n11, n12, n13, n1, n2, n4, n5, n6;
  assign mem_to_reg[1] = reg_dst[1];
  assign alu_src = alu_op[1];
  assign mem_read = mem_to_reg[0];

  NOR4_X2 U8 ( .A1(n2), .A2(n4), .A3(opcode[2]), .A4(reset), .ZN(reg_dst[1])
         );
  NOR2_X1 U3 ( .A1(n12), .A2(reset), .ZN(alu_op[1]) );
  NOR4_X4 U4 ( .A1(n2), .A2(n5), .A3(opcode[1]), .A4(reset), .ZN(mem_write) );
  INV_X1 U5 ( .A(n9), .ZN(mem_to_reg[0]) );
  AND2_X1 U6 ( .A1(n2), .A2(n7), .ZN(reg_dst[0]) );
  OR3_X1 U7 ( .A1(mem_to_reg[0]), .A2(mem_write), .A3(branch), .ZN(alu_op[0])
         );
  AND2_X1 U9 ( .A1(n5), .A2(n11), .ZN(jump) );
  NAND2_X1 U10 ( .A1(opcode[0]), .A2(n7), .ZN(sign_or_zero) );
  NOR3_X1 U11 ( .A1(n4), .A2(n5), .A3(n2), .ZN(n10) );
  OAI211_X1 U12 ( .C1(reset), .C2(n8), .A(n9), .B(n1), .ZN(reg_write) );
  AOI21_X1 U13 ( .B1(n4), .B2(n5), .A(n10), .ZN(n8) );
  INV_X1 U14 ( .A(reg_dst[1]), .ZN(n1) );
  AOI211_X1 U15 ( .C1(n4), .C2(opcode[0]), .A(n13), .B(n10), .ZN(n12) );
  NOR3_X1 U16 ( .A1(opcode[2]), .A2(reset), .A3(opcode[1]), .ZN(n7) );
  NOR2_X1 U17 ( .A1(n4), .A2(reset), .ZN(n11) );
  NAND2_X1 U18 ( .A1(n13), .A2(n6), .ZN(n9) );
  INV_X1 U19 ( .A(reset), .ZN(n6) );
  AND2_X1 U20 ( .A1(n11), .A2(opcode[2]), .ZN(branch) );
  INV_X1 U21 ( .A(opcode[1]), .ZN(n4) );
  INV_X1 U22 ( .A(opcode[2]), .ZN(n5) );
  INV_X1 U23 ( .A(opcode[0]), .ZN(n2) );
  NOR3_X1 U24 ( .A1(opcode[0]), .A2(opcode[1]), .A3(n5), .ZN(n13) );
endmodule


module register_file ( clk, rst, reg_write_en, reg_write_dest, reg_write_data, 
        reg_read_addr_1, reg_read_data_1, reg_read_addr_2, reg_read_data_2 );
  input [2:0] reg_write_dest;
  input [15:0] reg_write_data;
  input [2:0] reg_read_addr_1;
  output [15:0] reg_read_data_1;
  input [2:0] reg_read_addr_2;
  output [15:0] reg_read_data_2;
  input clk, rst, reg_write_en;
  wire   N29, N30, N31, N32, N33, N34, N35, N36, N37, N38, N39, N40, N41, N42,
         N43, N44, N45, N46, N47, N48, N49, N50, N51, N52, N53, N54, N55, N56,
         N57, N58, N59, N60, n21, n22, n23, n24, n25, n26, n27, n28, n2900,
         n3000, n3100, n3200, n3300, n3400, n3500, n3600, n3700, n3800, n3900,
         n4000, n4100, n4200, n4300, n4400, n4500, n4600, n4700, n4800, n4900,
         n5000, n510, n520, n530, n540, n550, n560, n570, n580, n590, n600,
         n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74,
         n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88,
         n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101,
         n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112,
         n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123,
         n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134,
         n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145,
         n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156,
         n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167,
         n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178,
         n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189,
         n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200,
         n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211,
         n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222,
         n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233,
         n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244,
         n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255,
         n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266,
         n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277,
         n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n1410, n1510,
         n1610, n1710, n1810, n1910, n20, n289, n2901, n291, n292, n293, n294,
         n295, n296, n297, n298, n299, n3001, n301, n302, n303, n304, n305,
         n306, n307, n308, n309, n3101, n311, n312, n313, n314, n315, n316,
         n317, n318, n319, n3201, n321, n322, n323, n324, n325, n326, n327,
         n328, n329, n3301, n331, n332, n333, n334, n335, n336, n337, n338,
         n339, n3401, n341, n342, n343, n344, n345, n346, n347, n348, n349,
         n3501, n351, n352, n353, n354, n355, n356, n357, n358, n359, n3601,
         n361, n362, n363, n364, n365, n366, n367, n368, n369, n3701, n371,
         n372, n373, n374, n375, n376, n377, n378, n379, n3801, n381, n382,
         n383, n384, n385, n386, n387, n388, n389, n3901, n391, n392, n393,
         n394, n395, n396, n397, n398, n399, n4001, n401, n402, n403, n404,
         n405, n406, n407, n408, n409, n4101, n411, n412, n413, n414, n415,
         n416, n417, n418, n419, n4201, n421, n422, n423, n424, n425, n426,
         n427, n428, n429, n4301, n431, n432, n433, n434, n435, n436, n437,
         n438, n439, n4401, n441, n442, n443, n444, n445, n446, n447, n448,
         n449, n4501, n451, n452, n453, n454, n455, n456, n457, n458, n459,
         n4601, n461, n462, n463, n464, n465, n466, n467, n468, n469, n4701,
         n471, n472, n473, n474, n475, n476, n477, n478, n479, n4801, n481,
         n482, n483, n484, n485, n486, n487, n488, n489, n4901, n491, n492,
         n493, n494, n495, n496, n497, n498, n499, n5001, n501, n502, n503,
         n504;
  wire   [127:0] reg_array;

  DFFR_X1 reg_array_reg_7__15_ ( .D(n288), .CK(clk), .RN(n504), .Q(
        reg_array[127]) );
  DFFR_X1 reg_array_reg_7__14_ ( .D(n287), .CK(clk), .RN(n504), .Q(
        reg_array[126]) );
  DFFR_X1 reg_array_reg_7__13_ ( .D(n286), .CK(clk), .RN(n504), .Q(
        reg_array[125]) );
  DFFR_X1 reg_array_reg_7__12_ ( .D(n285), .CK(clk), .RN(n504), .Q(
        reg_array[124]) );
  DFFR_X1 reg_array_reg_7__11_ ( .D(n284), .CK(clk), .RN(n504), .Q(
        reg_array[123]) );
  DFFR_X1 reg_array_reg_7__10_ ( .D(n283), .CK(clk), .RN(n504), .Q(
        reg_array[122]) );
  DFFR_X1 reg_array_reg_7__9_ ( .D(n282), .CK(clk), .RN(n504), .Q(
        reg_array[121]) );
  DFFR_X1 reg_array_reg_7__8_ ( .D(n281), .CK(clk), .RN(n504), .Q(
        reg_array[120]) );
  DFFR_X1 reg_array_reg_7__7_ ( .D(n280), .CK(clk), .RN(n504), .Q(
        reg_array[119]) );
  DFFR_X1 reg_array_reg_7__6_ ( .D(n279), .CK(clk), .RN(n504), .Q(
        reg_array[118]) );
  DFFR_X1 reg_array_reg_7__5_ ( .D(n278), .CK(clk), .RN(n504), .Q(
        reg_array[117]) );
  DFFR_X1 reg_array_reg_7__4_ ( .D(n277), .CK(clk), .RN(n504), .Q(
        reg_array[116]) );
  DFFR_X1 reg_array_reg_7__3_ ( .D(n276), .CK(clk), .RN(n504), .Q(
        reg_array[115]) );
  DFFR_X1 reg_array_reg_7__2_ ( .D(n275), .CK(clk), .RN(n504), .Q(
        reg_array[114]) );
  DFFR_X1 reg_array_reg_7__1_ ( .D(n274), .CK(clk), .RN(n504), .Q(
        reg_array[113]) );
  DFFR_X1 reg_array_reg_7__0_ ( .D(n273), .CK(clk), .RN(n504), .Q(
        reg_array[112]) );
  DFFR_X1 reg_array_reg_5__15_ ( .D(n256), .CK(clk), .RN(n504), .Q(
        reg_array[95]) );
  DFFR_X1 reg_array_reg_5__14_ ( .D(n255), .CK(clk), .RN(n504), .Q(
        reg_array[94]) );
  DFFR_X1 reg_array_reg_5__13_ ( .D(n254), .CK(clk), .RN(n504), .Q(
        reg_array[93]) );
  DFFR_X1 reg_array_reg_5__12_ ( .D(n253), .CK(clk), .RN(n504), .Q(
        reg_array[92]) );
  DFFR_X1 reg_array_reg_5__11_ ( .D(n252), .CK(clk), .RN(n504), .Q(
        reg_array[91]) );
  DFFR_X1 reg_array_reg_5__10_ ( .D(n251), .CK(clk), .RN(n504), .Q(
        reg_array[90]) );
  DFFR_X1 reg_array_reg_5__9_ ( .D(n250), .CK(clk), .RN(n504), .Q(
        reg_array[89]) );
  DFFR_X1 reg_array_reg_5__8_ ( .D(n249), .CK(clk), .RN(n504), .Q(
        reg_array[88]) );
  DFFR_X1 reg_array_reg_5__7_ ( .D(n248), .CK(clk), .RN(n504), .Q(
        reg_array[87]) );
  DFFR_X1 reg_array_reg_5__6_ ( .D(n247), .CK(clk), .RN(n504), .Q(
        reg_array[86]) );
  DFFR_X1 reg_array_reg_5__5_ ( .D(n246), .CK(clk), .RN(n504), .Q(
        reg_array[85]) );
  DFFR_X1 reg_array_reg_5__4_ ( .D(n245), .CK(clk), .RN(n504), .Q(
        reg_array[84]) );
  DFFR_X1 reg_array_reg_5__3_ ( .D(n244), .CK(clk), .RN(n504), .Q(
        reg_array[83]) );
  DFFR_X1 reg_array_reg_5__2_ ( .D(n243), .CK(clk), .RN(n504), .Q(
        reg_array[82]) );
  DFFR_X1 reg_array_reg_5__1_ ( .D(n242), .CK(clk), .RN(n504), .Q(
        reg_array[81]) );
  DFFR_X1 reg_array_reg_5__0_ ( .D(n241), .CK(clk), .RN(n504), .Q(
        reg_array[80]) );
  DFFR_X1 reg_array_reg_3__15_ ( .D(n224), .CK(clk), .RN(n504), .Q(
        reg_array[63]) );
  DFFR_X1 reg_array_reg_3__14_ ( .D(n223), .CK(clk), .RN(n504), .Q(
        reg_array[62]) );
  DFFR_X1 reg_array_reg_3__13_ ( .D(n222), .CK(clk), .RN(n504), .Q(
        reg_array[61]) );
  DFFR_X1 reg_array_reg_3__12_ ( .D(n221), .CK(clk), .RN(n504), .Q(
        reg_array[60]) );
  DFFR_X1 reg_array_reg_3__11_ ( .D(n220), .CK(clk), .RN(n504), .Q(
        reg_array[59]) );
  DFFR_X1 reg_array_reg_3__10_ ( .D(n219), .CK(clk), .RN(n504), .Q(
        reg_array[58]) );
  DFFR_X1 reg_array_reg_3__9_ ( .D(n218), .CK(clk), .RN(n504), .Q(
        reg_array[57]) );
  DFFR_X1 reg_array_reg_3__8_ ( .D(n217), .CK(clk), .RN(n504), .Q(
        reg_array[56]) );
  DFFR_X1 reg_array_reg_3__7_ ( .D(n216), .CK(clk), .RN(n504), .Q(
        reg_array[55]) );
  DFFR_X1 reg_array_reg_3__6_ ( .D(n215), .CK(clk), .RN(n504), .Q(
        reg_array[54]) );
  DFFR_X1 reg_array_reg_3__5_ ( .D(n214), .CK(clk), .RN(n504), .Q(
        reg_array[53]) );
  DFFR_X1 reg_array_reg_3__4_ ( .D(n213), .CK(clk), .RN(n504), .Q(
        reg_array[52]) );
  DFFR_X1 reg_array_reg_3__3_ ( .D(n212), .CK(clk), .RN(n504), .Q(
        reg_array[51]) );
  DFFR_X1 reg_array_reg_3__2_ ( .D(n211), .CK(clk), .RN(n504), .Q(
        reg_array[50]) );
  DFFR_X1 reg_array_reg_3__1_ ( .D(n210), .CK(clk), .RN(n504), .Q(
        reg_array[49]) );
  DFFR_X1 reg_array_reg_3__0_ ( .D(n209), .CK(clk), .RN(n504), .Q(
        reg_array[48]) );
  DFFR_X1 reg_array_reg_1__15_ ( .D(n192), .CK(clk), .RN(n504), .Q(
        reg_array[31]) );
  DFFR_X1 reg_array_reg_1__14_ ( .D(n191), .CK(clk), .RN(n504), .Q(
        reg_array[30]) );
  DFFR_X1 reg_array_reg_1__13_ ( .D(n190), .CK(clk), .RN(n504), .Q(
        reg_array[29]) );
  DFFR_X1 reg_array_reg_1__12_ ( .D(n189), .CK(clk), .RN(n504), .Q(
        reg_array[28]) );
  DFFR_X1 reg_array_reg_1__11_ ( .D(n188), .CK(clk), .RN(n504), .Q(
        reg_array[27]) );
  DFFR_X1 reg_array_reg_1__10_ ( .D(n187), .CK(clk), .RN(n504), .Q(
        reg_array[26]) );
  DFFR_X1 reg_array_reg_1__9_ ( .D(n186), .CK(clk), .RN(n504), .Q(
        reg_array[25]) );
  DFFR_X1 reg_array_reg_1__8_ ( .D(n185), .CK(clk), .RN(n504), .Q(
        reg_array[24]) );
  DFFR_X1 reg_array_reg_1__7_ ( .D(n184), .CK(clk), .RN(n504), .Q(
        reg_array[23]) );
  DFFR_X1 reg_array_reg_1__6_ ( .D(n183), .CK(clk), .RN(n504), .Q(
        reg_array[22]) );
  DFFR_X1 reg_array_reg_1__5_ ( .D(n182), .CK(clk), .RN(n504), .Q(
        reg_array[21]) );
  DFFR_X1 reg_array_reg_1__4_ ( .D(n181), .CK(clk), .RN(n504), .Q(
        reg_array[20]) );
  DFFR_X1 reg_array_reg_1__3_ ( .D(n180), .CK(clk), .RN(n504), .Q(
        reg_array[19]) );
  DFFR_X1 reg_array_reg_1__2_ ( .D(n179), .CK(clk), .RN(n504), .Q(
        reg_array[18]) );
  DFFR_X1 reg_array_reg_1__1_ ( .D(n178), .CK(clk), .RN(n504), .Q(
        reg_array[17]) );
  DFFR_X1 reg_array_reg_1__0_ ( .D(n177), .CK(clk), .RN(n504), .Q(
        reg_array[16]) );
  DFFR_X1 reg_array_reg_6__15_ ( .D(n272), .CK(clk), .RN(n504), .Q(
        reg_array[111]) );
  DFFR_X1 reg_array_reg_6__14_ ( .D(n271), .CK(clk), .RN(n504), .Q(
        reg_array[110]) );
  DFFR_X1 reg_array_reg_6__13_ ( .D(n270), .CK(clk), .RN(n504), .Q(
        reg_array[109]) );
  DFFR_X1 reg_array_reg_6__12_ ( .D(n269), .CK(clk), .RN(n504), .Q(
        reg_array[108]) );
  DFFR_X1 reg_array_reg_6__11_ ( .D(n268), .CK(clk), .RN(n504), .Q(
        reg_array[107]) );
  DFFR_X1 reg_array_reg_6__10_ ( .D(n267), .CK(clk), .RN(n504), .Q(
        reg_array[106]) );
  DFFR_X1 reg_array_reg_6__9_ ( .D(n266), .CK(clk), .RN(n504), .Q(
        reg_array[105]) );
  DFFR_X1 reg_array_reg_6__8_ ( .D(n265), .CK(clk), .RN(n504), .Q(
        reg_array[104]) );
  DFFR_X1 reg_array_reg_6__7_ ( .D(n264), .CK(clk), .RN(n504), .Q(
        reg_array[103]) );
  DFFR_X1 reg_array_reg_6__6_ ( .D(n263), .CK(clk), .RN(n504), .Q(
        reg_array[102]) );
  DFFR_X1 reg_array_reg_6__5_ ( .D(n262), .CK(clk), .RN(n504), .Q(
        reg_array[101]) );
  DFFR_X1 reg_array_reg_6__4_ ( .D(n261), .CK(clk), .RN(n504), .Q(
        reg_array[100]) );
  DFFR_X1 reg_array_reg_6__3_ ( .D(n260), .CK(clk), .RN(n504), .Q(
        reg_array[99]) );
  DFFR_X1 reg_array_reg_6__2_ ( .D(n259), .CK(clk), .RN(n504), .Q(
        reg_array[98]) );
  DFFR_X1 reg_array_reg_6__1_ ( .D(n258), .CK(clk), .RN(n504), .Q(
        reg_array[97]) );
  DFFR_X1 reg_array_reg_6__0_ ( .D(n257), .CK(clk), .RN(n504), .Q(
        reg_array[96]) );
  DFFR_X1 reg_array_reg_4__15_ ( .D(n240), .CK(clk), .RN(n504), .Q(
        reg_array[79]) );
  DFFR_X1 reg_array_reg_4__14_ ( .D(n239), .CK(clk), .RN(n504), .Q(
        reg_array[78]) );
  DFFR_X1 reg_array_reg_4__13_ ( .D(n238), .CK(clk), .RN(n504), .Q(
        reg_array[77]) );
  DFFR_X1 reg_array_reg_4__12_ ( .D(n237), .CK(clk), .RN(n504), .Q(
        reg_array[76]) );
  DFFR_X1 reg_array_reg_4__11_ ( .D(n236), .CK(clk), .RN(n504), .Q(
        reg_array[75]) );
  DFFR_X1 reg_array_reg_4__10_ ( .D(n235), .CK(clk), .RN(n504), .Q(
        reg_array[74]) );
  DFFR_X1 reg_array_reg_4__9_ ( .D(n234), .CK(clk), .RN(n504), .Q(
        reg_array[73]) );
  DFFR_X1 reg_array_reg_4__8_ ( .D(n233), .CK(clk), .RN(n504), .Q(
        reg_array[72]) );
  DFFR_X1 reg_array_reg_4__7_ ( .D(n232), .CK(clk), .RN(n504), .Q(
        reg_array[71]) );
  DFFR_X1 reg_array_reg_4__6_ ( .D(n231), .CK(clk), .RN(n504), .Q(
        reg_array[70]) );
  DFFR_X1 reg_array_reg_4__5_ ( .D(n230), .CK(clk), .RN(n504), .Q(
        reg_array[69]) );
  DFFR_X1 reg_array_reg_4__4_ ( .D(n229), .CK(clk), .RN(n504), .Q(
        reg_array[68]) );
  DFFR_X1 reg_array_reg_4__3_ ( .D(n228), .CK(clk), .RN(n504), .Q(
        reg_array[67]) );
  DFFR_X1 reg_array_reg_4__2_ ( .D(n227), .CK(clk), .RN(n504), .Q(
        reg_array[66]) );
  DFFR_X1 reg_array_reg_4__1_ ( .D(n226), .CK(clk), .RN(n504), .Q(
        reg_array[65]) );
  DFFR_X1 reg_array_reg_4__0_ ( .D(n225), .CK(clk), .RN(n504), .Q(
        reg_array[64]) );
  DFFR_X1 reg_array_reg_2__15_ ( .D(n208), .CK(clk), .RN(n504), .Q(
        reg_array[47]) );
  DFFR_X1 reg_array_reg_2__14_ ( .D(n207), .CK(clk), .RN(n504), .Q(
        reg_array[46]) );
  DFFR_X1 reg_array_reg_2__13_ ( .D(n206), .CK(clk), .RN(n504), .Q(
        reg_array[45]) );
  DFFR_X1 reg_array_reg_2__12_ ( .D(n205), .CK(clk), .RN(n504), .Q(
        reg_array[44]) );
  DFFR_X1 reg_array_reg_2__11_ ( .D(n204), .CK(clk), .RN(n504), .Q(
        reg_array[43]) );
  DFFR_X1 reg_array_reg_2__10_ ( .D(n203), .CK(clk), .RN(n504), .Q(
        reg_array[42]) );
  DFFR_X1 reg_array_reg_2__9_ ( .D(n202), .CK(clk), .RN(n504), .Q(
        reg_array[41]) );
  DFFR_X1 reg_array_reg_2__8_ ( .D(n201), .CK(clk), .RN(n504), .Q(
        reg_array[40]) );
  DFFR_X1 reg_array_reg_2__7_ ( .D(n200), .CK(clk), .RN(n504), .Q(
        reg_array[39]) );
  DFFR_X1 reg_array_reg_2__6_ ( .D(n199), .CK(clk), .RN(n504), .Q(
        reg_array[38]) );
  DFFR_X1 reg_array_reg_2__5_ ( .D(n198), .CK(clk), .RN(n504), .Q(
        reg_array[37]) );
  DFFR_X1 reg_array_reg_2__4_ ( .D(n197), .CK(clk), .RN(n504), .Q(
        reg_array[36]) );
  DFFR_X1 reg_array_reg_2__3_ ( .D(n196), .CK(clk), .RN(n504), .Q(
        reg_array[35]) );
  DFFR_X1 reg_array_reg_2__2_ ( .D(n195), .CK(clk), .RN(n504), .Q(
        reg_array[34]) );
  DFFR_X1 reg_array_reg_2__1_ ( .D(n194), .CK(clk), .RN(n504), .Q(
        reg_array[33]) );
  DFFR_X1 reg_array_reg_2__0_ ( .D(n193), .CK(clk), .RN(n504), .Q(
        reg_array[32]) );
  DFFR_X1 reg_array_reg_0__15_ ( .D(n176), .CK(clk), .RN(n504), .Q(
        reg_array[15]) );
  DFFR_X1 reg_array_reg_0__14_ ( .D(n175), .CK(clk), .RN(n504), .Q(
        reg_array[14]) );
  DFFR_X1 reg_array_reg_0__13_ ( .D(n174), .CK(clk), .RN(n504), .Q(
        reg_array[13]) );
  DFFR_X1 reg_array_reg_0__12_ ( .D(n173), .CK(clk), .RN(n504), .Q(
        reg_array[12]) );
  DFFR_X1 reg_array_reg_0__11_ ( .D(n172), .CK(clk), .RN(n504), .Q(
        reg_array[11]) );
  DFFR_X1 reg_array_reg_0__10_ ( .D(n171), .CK(clk), .RN(n504), .Q(
        reg_array[10]) );
  DFFR_X1 reg_array_reg_0__9_ ( .D(n170), .CK(clk), .RN(n504), .Q(reg_array[9]) );
  DFFR_X1 reg_array_reg_0__8_ ( .D(n169), .CK(clk), .RN(n504), .Q(reg_array[8]) );
  DFFR_X1 reg_array_reg_0__3_ ( .D(n164), .CK(clk), .RN(n504), .Q(reg_array[3]) );
  DFFR_X1 reg_array_reg_0__2_ ( .D(n163), .CK(clk), .RN(n504), .Q(reg_array[2]) );
  DFFR_X1 reg_array_reg_0__1_ ( .D(n162), .CK(clk), .RN(n504), .Q(reg_array[1]) );
  DFFR_X1 reg_array_reg_0__0_ ( .D(n161), .CK(clk), .RN(n504), .Q(reg_array[0]) );
  DFFR_X1 reg_array_reg_0__7_ ( .D(n168), .CK(clk), .RN(n504), .Q(reg_array[7]) );
  DFFR_X1 reg_array_reg_0__6_ ( .D(n167), .CK(clk), .RN(n504), .Q(reg_array[6]) );
  DFFR_X1 reg_array_reg_0__5_ ( .D(n166), .CK(clk), .RN(n504), .Q(reg_array[5]) );
  DFFR_X1 reg_array_reg_0__4_ ( .D(n165), .CK(clk), .RN(n504), .Q(reg_array[4]) );
  INV_X8 U2 ( .A(rst), .ZN(n504) );
  BUF_X1 U3 ( .A(n23), .Z(n483) );
  BUF_X1 U4 ( .A(n23), .Z(n482) );
  BUF_X1 U5 ( .A(n4100), .Z(n481) );
  BUF_X1 U6 ( .A(n580), .Z(n478) );
  BUF_X1 U7 ( .A(n75), .Z(n475) );
  BUF_X1 U8 ( .A(n92), .Z(n472) );
  BUF_X1 U9 ( .A(n110), .Z(n469) );
  BUF_X1 U10 ( .A(n127), .Z(n466) );
  BUF_X1 U11 ( .A(n144), .Z(n463) );
  BUF_X1 U12 ( .A(n23), .Z(n484) );
  BUF_X1 U13 ( .A(n4100), .Z(n479) );
  BUF_X1 U14 ( .A(n580), .Z(n476) );
  BUF_X1 U15 ( .A(n75), .Z(n473) );
  BUF_X1 U16 ( .A(n92), .Z(n4701) );
  BUF_X1 U17 ( .A(n110), .Z(n467) );
  BUF_X1 U18 ( .A(n127), .Z(n464) );
  BUF_X1 U19 ( .A(n144), .Z(n461) );
  BUF_X1 U20 ( .A(n4100), .Z(n4801) );
  BUF_X1 U21 ( .A(n580), .Z(n477) );
  BUF_X1 U22 ( .A(n75), .Z(n474) );
  BUF_X1 U23 ( .A(n92), .Z(n471) );
  BUF_X1 U24 ( .A(n110), .Z(n468) );
  BUF_X1 U25 ( .A(n127), .Z(n465) );
  BUF_X1 U26 ( .A(n144), .Z(n462) );
  INV_X1 U27 ( .A(reg_write_dest[1]), .ZN(n502) );
  INV_X1 U28 ( .A(reg_write_dest[0]), .ZN(n501) );
  NAND3_X1 U29 ( .A1(n501), .A2(n502), .A3(n4000), .ZN(n23) );
  INV_X1 U30 ( .A(reg_write_data[15]), .ZN(n485) );
  NAND3_X1 U31 ( .A1(n4000), .A2(n502), .A3(reg_write_dest[0]), .ZN(n4100) );
  NAND3_X1 U32 ( .A1(n4000), .A2(n501), .A3(reg_write_dest[1]), .ZN(n580) );
  NAND3_X1 U33 ( .A1(reg_write_dest[0]), .A2(n4000), .A3(reg_write_dest[1]), 
        .ZN(n75) );
  NAND3_X1 U34 ( .A1(reg_write_dest[1]), .A2(n501), .A3(n109), .ZN(n127) );
  NAND3_X1 U35 ( .A1(reg_write_dest[1]), .A2(reg_write_dest[0]), .A3(n109), 
        .ZN(n144) );
  NAND3_X1 U36 ( .A1(reg_write_dest[0]), .A2(n502), .A3(n109), .ZN(n110) );
  NAND3_X1 U37 ( .A1(n501), .A2(n502), .A3(n109), .ZN(n92) );
  NOR2_X1 U38 ( .A1(n503), .A2(reg_write_dest[2]), .ZN(n4000) );
  INV_X1 U39 ( .A(reg_write_en), .ZN(n503) );
  INV_X1 U40 ( .A(reg_write_data[2]), .ZN(n498) );
  INV_X1 U41 ( .A(reg_write_data[3]), .ZN(n497) );
  INV_X1 U42 ( .A(reg_write_data[4]), .ZN(n496) );
  INV_X1 U43 ( .A(reg_write_data[5]), .ZN(n495) );
  INV_X1 U44 ( .A(reg_write_data[6]), .ZN(n494) );
  INV_X1 U45 ( .A(reg_write_data[7]), .ZN(n493) );
  INV_X1 U46 ( .A(reg_write_data[8]), .ZN(n492) );
  INV_X1 U47 ( .A(reg_write_data[9]), .ZN(n491) );
  INV_X1 U48 ( .A(reg_write_data[10]), .ZN(n4901) );
  INV_X1 U49 ( .A(reg_write_data[11]), .ZN(n489) );
  INV_X1 U50 ( .A(reg_write_data[12]), .ZN(n488) );
  INV_X1 U51 ( .A(reg_write_data[13]), .ZN(n487) );
  INV_X1 U52 ( .A(reg_write_data[14]), .ZN(n486) );
  AND2_X1 U53 ( .A1(reg_write_dest[2]), .A2(reg_write_en), .ZN(n109) );
  OAI21_X1 U54 ( .B1(n483), .B2(n496), .A(n28), .ZN(n165) );
  NAND2_X1 U55 ( .A1(reg_array[4]), .A2(n483), .ZN(n28) );
  OAI21_X1 U56 ( .B1(n483), .B2(n495), .A(n2900), .ZN(n166) );
  NAND2_X1 U57 ( .A1(reg_array[5]), .A2(n483), .ZN(n2900) );
  OAI21_X1 U58 ( .B1(n483), .B2(n494), .A(n3000), .ZN(n167) );
  NAND2_X1 U59 ( .A1(reg_array[6]), .A2(n483), .ZN(n3000) );
  OAI21_X1 U60 ( .B1(n483), .B2(n493), .A(n3100), .ZN(n168) );
  NAND2_X1 U61 ( .A1(reg_array[7]), .A2(n483), .ZN(n3100) );
  OAI21_X1 U62 ( .B1(n483), .B2(n5001), .A(n24), .ZN(n161) );
  NAND2_X1 U63 ( .A1(reg_array[0]), .A2(n482), .ZN(n24) );
  OAI21_X1 U64 ( .B1(n483), .B2(n499), .A(n25), .ZN(n162) );
  NAND2_X1 U65 ( .A1(reg_array[1]), .A2(n482), .ZN(n25) );
  OAI21_X1 U66 ( .B1(n483), .B2(n498), .A(n26), .ZN(n163) );
  NAND2_X1 U67 ( .A1(reg_array[2]), .A2(n482), .ZN(n26) );
  OAI21_X1 U68 ( .B1(n483), .B2(n497), .A(n27), .ZN(n164) );
  NAND2_X1 U69 ( .A1(reg_array[3]), .A2(n482), .ZN(n27) );
  OAI21_X1 U70 ( .B1(n484), .B2(n492), .A(n3200), .ZN(n169) );
  NAND2_X1 U71 ( .A1(reg_array[8]), .A2(n482), .ZN(n3200) );
  OAI21_X1 U72 ( .B1(n484), .B2(n491), .A(n3300), .ZN(n170) );
  NAND2_X1 U73 ( .A1(reg_array[9]), .A2(n482), .ZN(n3300) );
  OAI21_X1 U74 ( .B1(n484), .B2(n4901), .A(n3400), .ZN(n171) );
  NAND2_X1 U75 ( .A1(reg_array[10]), .A2(n482), .ZN(n3400) );
  OAI21_X1 U76 ( .B1(n484), .B2(n489), .A(n3500), .ZN(n172) );
  NAND2_X1 U77 ( .A1(reg_array[11]), .A2(n482), .ZN(n3500) );
  OAI21_X1 U78 ( .B1(n484), .B2(n488), .A(n3600), .ZN(n173) );
  NAND2_X1 U79 ( .A1(reg_array[12]), .A2(n482), .ZN(n3600) );
  OAI21_X1 U80 ( .B1(n484), .B2(n487), .A(n3700), .ZN(n174) );
  NAND2_X1 U81 ( .A1(reg_array[13]), .A2(n482), .ZN(n3700) );
  OAI21_X1 U82 ( .B1(n484), .B2(n486), .A(n3800), .ZN(n175) );
  NAND2_X1 U83 ( .A1(reg_array[14]), .A2(n482), .ZN(n3800) );
  OAI21_X1 U84 ( .B1(n483), .B2(n485), .A(n3900), .ZN(n176) );
  NAND2_X1 U85 ( .A1(reg_array[15]), .A2(n482), .ZN(n3900) );
  OAI21_X1 U86 ( .B1(n5001), .B2(n4801), .A(n4200), .ZN(n177) );
  NAND2_X1 U87 ( .A1(reg_array[16]), .A2(n479), .ZN(n4200) );
  OAI21_X1 U88 ( .B1(n499), .B2(n4801), .A(n4300), .ZN(n178) );
  NAND2_X1 U89 ( .A1(reg_array[17]), .A2(n479), .ZN(n4300) );
  OAI21_X1 U90 ( .B1(n498), .B2(n4801), .A(n4400), .ZN(n179) );
  NAND2_X1 U91 ( .A1(reg_array[18]), .A2(n479), .ZN(n4400) );
  OAI21_X1 U92 ( .B1(n497), .B2(n4801), .A(n4500), .ZN(n180) );
  NAND2_X1 U93 ( .A1(reg_array[19]), .A2(n479), .ZN(n4500) );
  OAI21_X1 U94 ( .B1(n496), .B2(n4801), .A(n4600), .ZN(n181) );
  NAND2_X1 U95 ( .A1(reg_array[20]), .A2(n4801), .ZN(n4600) );
  OAI21_X1 U96 ( .B1(n495), .B2(n4801), .A(n4700), .ZN(n182) );
  NAND2_X1 U97 ( .A1(reg_array[21]), .A2(n4801), .ZN(n4700) );
  OAI21_X1 U98 ( .B1(n494), .B2(n4801), .A(n4800), .ZN(n183) );
  NAND2_X1 U99 ( .A1(reg_array[22]), .A2(n4801), .ZN(n4800) );
  OAI21_X1 U100 ( .B1(n493), .B2(n481), .A(n4900), .ZN(n184) );
  NAND2_X1 U101 ( .A1(reg_array[23]), .A2(n4801), .ZN(n4900) );
  OAI21_X1 U102 ( .B1(n492), .B2(n481), .A(n5000), .ZN(n185) );
  NAND2_X1 U103 ( .A1(reg_array[24]), .A2(n479), .ZN(n5000) );
  OAI21_X1 U104 ( .B1(n491), .B2(n481), .A(n510), .ZN(n186) );
  NAND2_X1 U105 ( .A1(reg_array[25]), .A2(n479), .ZN(n510) );
  OAI21_X1 U106 ( .B1(n4901), .B2(n481), .A(n520), .ZN(n187) );
  NAND2_X1 U107 ( .A1(reg_array[26]), .A2(n479), .ZN(n520) );
  OAI21_X1 U108 ( .B1(n489), .B2(n481), .A(n530), .ZN(n188) );
  NAND2_X1 U109 ( .A1(reg_array[27]), .A2(n479), .ZN(n530) );
  OAI21_X1 U110 ( .B1(n488), .B2(n481), .A(n540), .ZN(n189) );
  NAND2_X1 U111 ( .A1(reg_array[28]), .A2(n479), .ZN(n540) );
  OAI21_X1 U112 ( .B1(n487), .B2(n481), .A(n550), .ZN(n190) );
  NAND2_X1 U113 ( .A1(reg_array[29]), .A2(n479), .ZN(n550) );
  OAI21_X1 U114 ( .B1(n486), .B2(n481), .A(n560), .ZN(n191) );
  NAND2_X1 U115 ( .A1(reg_array[30]), .A2(n479), .ZN(n560) );
  OAI21_X1 U116 ( .B1(n485), .B2(n4801), .A(n570), .ZN(n192) );
  NAND2_X1 U117 ( .A1(reg_array[31]), .A2(n479), .ZN(n570) );
  OAI21_X1 U118 ( .B1(n5001), .B2(n477), .A(n590), .ZN(n193) );
  NAND2_X1 U119 ( .A1(reg_array[32]), .A2(n476), .ZN(n590) );
  OAI21_X1 U120 ( .B1(n499), .B2(n477), .A(n600), .ZN(n194) );
  NAND2_X1 U121 ( .A1(reg_array[33]), .A2(n476), .ZN(n600) );
  OAI21_X1 U122 ( .B1(n498), .B2(n477), .A(n61), .ZN(n195) );
  NAND2_X1 U123 ( .A1(reg_array[34]), .A2(n476), .ZN(n61) );
  OAI21_X1 U124 ( .B1(n497), .B2(n477), .A(n62), .ZN(n196) );
  NAND2_X1 U125 ( .A1(reg_array[35]), .A2(n476), .ZN(n62) );
  OAI21_X1 U126 ( .B1(n496), .B2(n477), .A(n63), .ZN(n197) );
  NAND2_X1 U127 ( .A1(reg_array[36]), .A2(n477), .ZN(n63) );
  OAI21_X1 U128 ( .B1(n495), .B2(n477), .A(n64), .ZN(n198) );
  NAND2_X1 U129 ( .A1(reg_array[37]), .A2(n477), .ZN(n64) );
  OAI21_X1 U130 ( .B1(n494), .B2(n477), .A(n65), .ZN(n199) );
  NAND2_X1 U131 ( .A1(reg_array[38]), .A2(n477), .ZN(n65) );
  OAI21_X1 U132 ( .B1(n493), .B2(n478), .A(n66), .ZN(n200) );
  NAND2_X1 U133 ( .A1(reg_array[39]), .A2(n477), .ZN(n66) );
  OAI21_X1 U134 ( .B1(n492), .B2(n478), .A(n67), .ZN(n201) );
  NAND2_X1 U135 ( .A1(reg_array[40]), .A2(n476), .ZN(n67) );
  OAI21_X1 U136 ( .B1(n491), .B2(n478), .A(n68), .ZN(n202) );
  NAND2_X1 U137 ( .A1(reg_array[41]), .A2(n476), .ZN(n68) );
  OAI21_X1 U138 ( .B1(n4901), .B2(n478), .A(n69), .ZN(n203) );
  NAND2_X1 U139 ( .A1(reg_array[42]), .A2(n476), .ZN(n69) );
  OAI21_X1 U140 ( .B1(n489), .B2(n478), .A(n70), .ZN(n204) );
  NAND2_X1 U141 ( .A1(reg_array[43]), .A2(n476), .ZN(n70) );
  OAI21_X1 U142 ( .B1(n488), .B2(n478), .A(n71), .ZN(n205) );
  NAND2_X1 U143 ( .A1(reg_array[44]), .A2(n476), .ZN(n71) );
  OAI21_X1 U144 ( .B1(n487), .B2(n478), .A(n72), .ZN(n206) );
  NAND2_X1 U145 ( .A1(reg_array[45]), .A2(n476), .ZN(n72) );
  OAI21_X1 U146 ( .B1(n486), .B2(n478), .A(n73), .ZN(n207) );
  NAND2_X1 U147 ( .A1(reg_array[46]), .A2(n476), .ZN(n73) );
  OAI21_X1 U148 ( .B1(n485), .B2(n477), .A(n74), .ZN(n208) );
  NAND2_X1 U149 ( .A1(reg_array[47]), .A2(n476), .ZN(n74) );
  OAI21_X1 U150 ( .B1(n5001), .B2(n474), .A(n76), .ZN(n209) );
  NAND2_X1 U151 ( .A1(reg_array[48]), .A2(n473), .ZN(n76) );
  OAI21_X1 U152 ( .B1(n499), .B2(n474), .A(n77), .ZN(n210) );
  NAND2_X1 U153 ( .A1(reg_array[49]), .A2(n473), .ZN(n77) );
  OAI21_X1 U154 ( .B1(n498), .B2(n474), .A(n78), .ZN(n211) );
  NAND2_X1 U155 ( .A1(reg_array[50]), .A2(n473), .ZN(n78) );
  OAI21_X1 U156 ( .B1(n497), .B2(n474), .A(n79), .ZN(n212) );
  NAND2_X1 U157 ( .A1(reg_array[51]), .A2(n473), .ZN(n79) );
  OAI21_X1 U158 ( .B1(n496), .B2(n474), .A(n80), .ZN(n213) );
  NAND2_X1 U159 ( .A1(reg_array[52]), .A2(n474), .ZN(n80) );
  OAI21_X1 U160 ( .B1(n495), .B2(n474), .A(n81), .ZN(n214) );
  NAND2_X1 U161 ( .A1(reg_array[53]), .A2(n474), .ZN(n81) );
  OAI21_X1 U162 ( .B1(n494), .B2(n474), .A(n82), .ZN(n215) );
  NAND2_X1 U163 ( .A1(reg_array[54]), .A2(n474), .ZN(n82) );
  OAI21_X1 U164 ( .B1(n493), .B2(n475), .A(n83), .ZN(n216) );
  NAND2_X1 U165 ( .A1(reg_array[55]), .A2(n474), .ZN(n83) );
  OAI21_X1 U166 ( .B1(n492), .B2(n475), .A(n84), .ZN(n217) );
  NAND2_X1 U167 ( .A1(reg_array[56]), .A2(n473), .ZN(n84) );
  OAI21_X1 U168 ( .B1(n491), .B2(n475), .A(n85), .ZN(n218) );
  NAND2_X1 U169 ( .A1(reg_array[57]), .A2(n473), .ZN(n85) );
  OAI21_X1 U170 ( .B1(n4901), .B2(n475), .A(n86), .ZN(n219) );
  NAND2_X1 U171 ( .A1(reg_array[58]), .A2(n473), .ZN(n86) );
  OAI21_X1 U172 ( .B1(n489), .B2(n475), .A(n87), .ZN(n220) );
  NAND2_X1 U173 ( .A1(reg_array[59]), .A2(n473), .ZN(n87) );
  OAI21_X1 U174 ( .B1(n488), .B2(n475), .A(n88), .ZN(n221) );
  NAND2_X1 U175 ( .A1(reg_array[60]), .A2(n473), .ZN(n88) );
  OAI21_X1 U176 ( .B1(n487), .B2(n475), .A(n89), .ZN(n222) );
  NAND2_X1 U177 ( .A1(reg_array[61]), .A2(n473), .ZN(n89) );
  OAI21_X1 U178 ( .B1(n486), .B2(n475), .A(n90), .ZN(n223) );
  NAND2_X1 U179 ( .A1(reg_array[62]), .A2(n473), .ZN(n90) );
  OAI21_X1 U180 ( .B1(n485), .B2(n474), .A(n91), .ZN(n224) );
  NAND2_X1 U181 ( .A1(reg_array[63]), .A2(n473), .ZN(n91) );
  OAI21_X1 U182 ( .B1(n5001), .B2(n471), .A(n93), .ZN(n225) );
  NAND2_X1 U183 ( .A1(reg_array[64]), .A2(n4701), .ZN(n93) );
  OAI21_X1 U184 ( .B1(n499), .B2(n471), .A(n94), .ZN(n226) );
  NAND2_X1 U185 ( .A1(reg_array[65]), .A2(n4701), .ZN(n94) );
  OAI21_X1 U186 ( .B1(n498), .B2(n471), .A(n95), .ZN(n227) );
  NAND2_X1 U187 ( .A1(reg_array[66]), .A2(n4701), .ZN(n95) );
  OAI21_X1 U188 ( .B1(n497), .B2(n471), .A(n96), .ZN(n228) );
  NAND2_X1 U189 ( .A1(reg_array[67]), .A2(n4701), .ZN(n96) );
  OAI21_X1 U190 ( .B1(n496), .B2(n471), .A(n97), .ZN(n229) );
  NAND2_X1 U191 ( .A1(reg_array[68]), .A2(n471), .ZN(n97) );
  OAI21_X1 U192 ( .B1(n495), .B2(n471), .A(n98), .ZN(n230) );
  NAND2_X1 U193 ( .A1(reg_array[69]), .A2(n471), .ZN(n98) );
  OAI21_X1 U194 ( .B1(n494), .B2(n471), .A(n99), .ZN(n231) );
  NAND2_X1 U195 ( .A1(reg_array[70]), .A2(n471), .ZN(n99) );
  OAI21_X1 U196 ( .B1(n493), .B2(n472), .A(n100), .ZN(n232) );
  NAND2_X1 U197 ( .A1(reg_array[71]), .A2(n471), .ZN(n100) );
  OAI21_X1 U198 ( .B1(n492), .B2(n472), .A(n101), .ZN(n233) );
  NAND2_X1 U199 ( .A1(reg_array[72]), .A2(n4701), .ZN(n101) );
  OAI21_X1 U200 ( .B1(n491), .B2(n472), .A(n102), .ZN(n234) );
  NAND2_X1 U201 ( .A1(reg_array[73]), .A2(n4701), .ZN(n102) );
  OAI21_X1 U202 ( .B1(n4901), .B2(n472), .A(n103), .ZN(n235) );
  NAND2_X1 U203 ( .A1(reg_array[74]), .A2(n4701), .ZN(n103) );
  OAI21_X1 U204 ( .B1(n489), .B2(n472), .A(n104), .ZN(n236) );
  NAND2_X1 U205 ( .A1(reg_array[75]), .A2(n4701), .ZN(n104) );
  OAI21_X1 U206 ( .B1(n488), .B2(n472), .A(n105), .ZN(n237) );
  NAND2_X1 U207 ( .A1(reg_array[76]), .A2(n4701), .ZN(n105) );
  OAI21_X1 U208 ( .B1(n487), .B2(n472), .A(n106), .ZN(n238) );
  NAND2_X1 U209 ( .A1(reg_array[77]), .A2(n4701), .ZN(n106) );
  OAI21_X1 U210 ( .B1(n486), .B2(n472), .A(n107), .ZN(n239) );
  NAND2_X1 U211 ( .A1(reg_array[78]), .A2(n4701), .ZN(n107) );
  OAI21_X1 U212 ( .B1(n485), .B2(n471), .A(n108), .ZN(n240) );
  NAND2_X1 U213 ( .A1(reg_array[79]), .A2(n4701), .ZN(n108) );
  OAI21_X1 U214 ( .B1(n5001), .B2(n468), .A(n111), .ZN(n241) );
  NAND2_X1 U215 ( .A1(reg_array[80]), .A2(n467), .ZN(n111) );
  OAI21_X1 U216 ( .B1(n499), .B2(n468), .A(n112), .ZN(n242) );
  NAND2_X1 U217 ( .A1(reg_array[81]), .A2(n467), .ZN(n112) );
  OAI21_X1 U218 ( .B1(n498), .B2(n468), .A(n113), .ZN(n243) );
  NAND2_X1 U219 ( .A1(reg_array[82]), .A2(n467), .ZN(n113) );
  OAI21_X1 U220 ( .B1(n497), .B2(n468), .A(n114), .ZN(n244) );
  NAND2_X1 U221 ( .A1(reg_array[83]), .A2(n467), .ZN(n114) );
  OAI21_X1 U222 ( .B1(n496), .B2(n468), .A(n115), .ZN(n245) );
  NAND2_X1 U223 ( .A1(reg_array[84]), .A2(n468), .ZN(n115) );
  OAI21_X1 U224 ( .B1(n495), .B2(n468), .A(n116), .ZN(n246) );
  NAND2_X1 U225 ( .A1(reg_array[85]), .A2(n468), .ZN(n116) );
  OAI21_X1 U226 ( .B1(n494), .B2(n468), .A(n117), .ZN(n247) );
  NAND2_X1 U227 ( .A1(reg_array[86]), .A2(n468), .ZN(n117) );
  OAI21_X1 U228 ( .B1(n493), .B2(n469), .A(n118), .ZN(n248) );
  NAND2_X1 U229 ( .A1(reg_array[87]), .A2(n468), .ZN(n118) );
  OAI21_X1 U230 ( .B1(n492), .B2(n469), .A(n119), .ZN(n249) );
  NAND2_X1 U231 ( .A1(reg_array[88]), .A2(n467), .ZN(n119) );
  OAI21_X1 U232 ( .B1(n491), .B2(n469), .A(n120), .ZN(n250) );
  NAND2_X1 U233 ( .A1(reg_array[89]), .A2(n467), .ZN(n120) );
  OAI21_X1 U234 ( .B1(n4901), .B2(n469), .A(n121), .ZN(n251) );
  NAND2_X1 U235 ( .A1(reg_array[90]), .A2(n467), .ZN(n121) );
  OAI21_X1 U236 ( .B1(n489), .B2(n469), .A(n122), .ZN(n252) );
  NAND2_X1 U237 ( .A1(reg_array[91]), .A2(n467), .ZN(n122) );
  OAI21_X1 U238 ( .B1(n488), .B2(n469), .A(n123), .ZN(n253) );
  NAND2_X1 U239 ( .A1(reg_array[92]), .A2(n467), .ZN(n123) );
  OAI21_X1 U240 ( .B1(n487), .B2(n469), .A(n124), .ZN(n254) );
  NAND2_X1 U241 ( .A1(reg_array[93]), .A2(n467), .ZN(n124) );
  OAI21_X1 U242 ( .B1(n486), .B2(n469), .A(n125), .ZN(n255) );
  NAND2_X1 U243 ( .A1(reg_array[94]), .A2(n467), .ZN(n125) );
  OAI21_X1 U244 ( .B1(n485), .B2(n468), .A(n126), .ZN(n256) );
  NAND2_X1 U245 ( .A1(reg_array[95]), .A2(n467), .ZN(n126) );
  OAI21_X1 U246 ( .B1(n5001), .B2(n465), .A(n128), .ZN(n257) );
  NAND2_X1 U247 ( .A1(reg_array[96]), .A2(n464), .ZN(n128) );
  OAI21_X1 U248 ( .B1(n499), .B2(n465), .A(n129), .ZN(n258) );
  NAND2_X1 U249 ( .A1(reg_array[97]), .A2(n464), .ZN(n129) );
  OAI21_X1 U250 ( .B1(n498), .B2(n465), .A(n130), .ZN(n259) );
  NAND2_X1 U251 ( .A1(reg_array[98]), .A2(n464), .ZN(n130) );
  OAI21_X1 U252 ( .B1(n497), .B2(n465), .A(n131), .ZN(n260) );
  NAND2_X1 U253 ( .A1(reg_array[99]), .A2(n464), .ZN(n131) );
  OAI21_X1 U254 ( .B1(n496), .B2(n465), .A(n132), .ZN(n261) );
  NAND2_X1 U255 ( .A1(reg_array[100]), .A2(n465), .ZN(n132) );
  OAI21_X1 U256 ( .B1(n495), .B2(n465), .A(n133), .ZN(n262) );
  NAND2_X1 U257 ( .A1(reg_array[101]), .A2(n465), .ZN(n133) );
  OAI21_X1 U258 ( .B1(n494), .B2(n465), .A(n134), .ZN(n263) );
  NAND2_X1 U259 ( .A1(reg_array[102]), .A2(n465), .ZN(n134) );
  OAI21_X1 U260 ( .B1(n493), .B2(n466), .A(n135), .ZN(n264) );
  NAND2_X1 U261 ( .A1(reg_array[103]), .A2(n465), .ZN(n135) );
  OAI21_X1 U262 ( .B1(n492), .B2(n466), .A(n136), .ZN(n265) );
  NAND2_X1 U263 ( .A1(reg_array[104]), .A2(n464), .ZN(n136) );
  OAI21_X1 U264 ( .B1(n491), .B2(n466), .A(n137), .ZN(n266) );
  NAND2_X1 U265 ( .A1(reg_array[105]), .A2(n464), .ZN(n137) );
  OAI21_X1 U266 ( .B1(n4901), .B2(n466), .A(n138), .ZN(n267) );
  NAND2_X1 U267 ( .A1(reg_array[106]), .A2(n464), .ZN(n138) );
  OAI21_X1 U268 ( .B1(n489), .B2(n466), .A(n139), .ZN(n268) );
  NAND2_X1 U269 ( .A1(reg_array[107]), .A2(n464), .ZN(n139) );
  OAI21_X1 U270 ( .B1(n488), .B2(n466), .A(n140), .ZN(n269) );
  NAND2_X1 U271 ( .A1(reg_array[108]), .A2(n464), .ZN(n140) );
  OAI21_X1 U272 ( .B1(n487), .B2(n466), .A(n141), .ZN(n270) );
  NAND2_X1 U273 ( .A1(reg_array[109]), .A2(n464), .ZN(n141) );
  OAI21_X1 U274 ( .B1(n486), .B2(n466), .A(n142), .ZN(n271) );
  NAND2_X1 U275 ( .A1(reg_array[110]), .A2(n464), .ZN(n142) );
  OAI21_X1 U276 ( .B1(n485), .B2(n465), .A(n143), .ZN(n272) );
  NAND2_X1 U277 ( .A1(reg_array[111]), .A2(n464), .ZN(n143) );
  OAI21_X1 U278 ( .B1(n5001), .B2(n462), .A(n145), .ZN(n273) );
  NAND2_X1 U279 ( .A1(reg_array[112]), .A2(n461), .ZN(n145) );
  OAI21_X1 U280 ( .B1(n499), .B2(n462), .A(n146), .ZN(n274) );
  NAND2_X1 U281 ( .A1(reg_array[113]), .A2(n461), .ZN(n146) );
  OAI21_X1 U282 ( .B1(n498), .B2(n462), .A(n147), .ZN(n275) );
  NAND2_X1 U283 ( .A1(reg_array[114]), .A2(n461), .ZN(n147) );
  OAI21_X1 U284 ( .B1(n497), .B2(n462), .A(n148), .ZN(n276) );
  NAND2_X1 U285 ( .A1(reg_array[115]), .A2(n461), .ZN(n148) );
  OAI21_X1 U286 ( .B1(n496), .B2(n462), .A(n149), .ZN(n277) );
  NAND2_X1 U287 ( .A1(reg_array[116]), .A2(n462), .ZN(n149) );
  OAI21_X1 U288 ( .B1(n495), .B2(n462), .A(n150), .ZN(n278) );
  NAND2_X1 U289 ( .A1(reg_array[117]), .A2(n462), .ZN(n150) );
  OAI21_X1 U290 ( .B1(n494), .B2(n462), .A(n151), .ZN(n279) );
  NAND2_X1 U291 ( .A1(reg_array[118]), .A2(n462), .ZN(n151) );
  OAI21_X1 U292 ( .B1(n493), .B2(n463), .A(n152), .ZN(n280) );
  NAND2_X1 U293 ( .A1(reg_array[119]), .A2(n462), .ZN(n152) );
  OAI21_X1 U294 ( .B1(n492), .B2(n463), .A(n153), .ZN(n281) );
  NAND2_X1 U295 ( .A1(reg_array[120]), .A2(n461), .ZN(n153) );
  OAI21_X1 U296 ( .B1(n491), .B2(n463), .A(n154), .ZN(n282) );
  NAND2_X1 U297 ( .A1(reg_array[121]), .A2(n461), .ZN(n154) );
  OAI21_X1 U298 ( .B1(n4901), .B2(n463), .A(n155), .ZN(n283) );
  NAND2_X1 U299 ( .A1(reg_array[122]), .A2(n461), .ZN(n155) );
  OAI21_X1 U300 ( .B1(n489), .B2(n463), .A(n156), .ZN(n284) );
  NAND2_X1 U301 ( .A1(reg_array[123]), .A2(n461), .ZN(n156) );
  OAI21_X1 U302 ( .B1(n488), .B2(n463), .A(n157), .ZN(n285) );
  NAND2_X1 U303 ( .A1(reg_array[124]), .A2(n461), .ZN(n157) );
  OAI21_X1 U304 ( .B1(n487), .B2(n463), .A(n158), .ZN(n286) );
  NAND2_X1 U305 ( .A1(reg_array[125]), .A2(n461), .ZN(n158) );
  OAI21_X1 U306 ( .B1(n486), .B2(n463), .A(n159), .ZN(n287) );
  NAND2_X1 U307 ( .A1(reg_array[126]), .A2(n461), .ZN(n159) );
  OAI21_X1 U308 ( .B1(n485), .B2(n462), .A(n160), .ZN(n288) );
  NAND2_X1 U309 ( .A1(reg_array[127]), .A2(n461), .ZN(n160) );
  INV_X1 U310 ( .A(reg_write_data[0]), .ZN(n5001) );
  INV_X1 U311 ( .A(reg_write_data[1]), .ZN(n499) );
  AND2_X1 U312 ( .A1(N44), .A2(n22), .ZN(reg_read_data_1[0]) );
  AND2_X1 U313 ( .A1(N29), .A2(n22), .ZN(reg_read_data_1[15]) );
  AND2_X1 U314 ( .A1(N37), .A2(n22), .ZN(reg_read_data_1[7]) );
  AND2_X1 U315 ( .A1(N34), .A2(n22), .ZN(reg_read_data_1[10]) );
  AND2_X1 U316 ( .A1(N33), .A2(n22), .ZN(reg_read_data_1[11]) );
  AND2_X1 U317 ( .A1(N31), .A2(n22), .ZN(reg_read_data_1[13]) );
  AND2_X1 U318 ( .A1(N41), .A2(n22), .ZN(reg_read_data_1[3]) );
  AND2_X1 U319 ( .A1(N39), .A2(n22), .ZN(reg_read_data_1[5]) );
  AND2_X1 U320 ( .A1(N43), .A2(n22), .ZN(reg_read_data_1[1]) );
  AND2_X1 U321 ( .A1(N38), .A2(n22), .ZN(reg_read_data_1[6]) );
  AND2_X1 U322 ( .A1(N36), .A2(n22), .ZN(reg_read_data_1[8]) );
  AND2_X1 U323 ( .A1(N35), .A2(n22), .ZN(reg_read_data_1[9]) );
  AND2_X1 U324 ( .A1(N32), .A2(n22), .ZN(reg_read_data_1[12]) );
  AND2_X1 U325 ( .A1(N42), .A2(n22), .ZN(reg_read_data_1[2]) );
  AND2_X1 U326 ( .A1(N40), .A2(n22), .ZN(reg_read_data_1[4]) );
  AND2_X1 U327 ( .A1(N30), .A2(n22), .ZN(reg_read_data_1[14]) );
  AND2_X1 U328 ( .A1(N53), .A2(n21), .ZN(reg_read_data_2[7]) );
  AND2_X1 U329 ( .A1(N52), .A2(n21), .ZN(reg_read_data_2[8]) );
  AND2_X1 U330 ( .A1(N51), .A2(n21), .ZN(reg_read_data_2[9]) );
  AND2_X1 U331 ( .A1(N50), .A2(n21), .ZN(reg_read_data_2[10]) );
  AND2_X1 U332 ( .A1(N49), .A2(n21), .ZN(reg_read_data_2[11]) );
  AND2_X1 U333 ( .A1(N48), .A2(n21), .ZN(reg_read_data_2[12]) );
  AND2_X1 U334 ( .A1(N47), .A2(n21), .ZN(reg_read_data_2[13]) );
  AND2_X1 U335 ( .A1(N46), .A2(n21), .ZN(reg_read_data_2[14]) );
  AND2_X1 U336 ( .A1(N45), .A2(n21), .ZN(reg_read_data_2[15]) );
  AND2_X1 U337 ( .A1(N60), .A2(n21), .ZN(reg_read_data_2[0]) );
  AND2_X1 U338 ( .A1(N59), .A2(n21), .ZN(reg_read_data_2[1]) );
  AND2_X1 U339 ( .A1(N58), .A2(n21), .ZN(reg_read_data_2[2]) );
  AND2_X1 U340 ( .A1(N57), .A2(n21), .ZN(reg_read_data_2[3]) );
  AND2_X1 U341 ( .A1(N56), .A2(n21), .ZN(reg_read_data_2[4]) );
  AND2_X1 U342 ( .A1(N55), .A2(n21), .ZN(reg_read_data_2[5]) );
  AND2_X1 U343 ( .A1(N54), .A2(n21), .ZN(reg_read_data_2[6]) );
  OR3_X1 U344 ( .A1(reg_read_addr_2[1]), .A2(reg_read_addr_2[2]), .A3(
        reg_read_addr_2[0]), .ZN(n21) );
  OR3_X1 U345 ( .A1(reg_read_addr_1[1]), .A2(reg_read_addr_1[2]), .A3(
        reg_read_addr_1[0]), .ZN(n22) );
  MUX2_X1 U346 ( .A(reg_array[96]), .B(reg_array[112]), .S(reg_read_addr_1[0]), 
        .Z(n1) );
  MUX2_X1 U347 ( .A(reg_array[64]), .B(reg_array[80]), .S(reg_read_addr_1[0]), 
        .Z(n2) );
  MUX2_X1 U348 ( .A(n2), .B(n1), .S(reg_read_addr_1[1]), .Z(n3) );
  MUX2_X1 U349 ( .A(reg_array[32]), .B(reg_array[48]), .S(reg_read_addr_1[0]), 
        .Z(n4) );
  MUX2_X1 U350 ( .A(reg_array[0]), .B(reg_array[16]), .S(reg_read_addr_1[0]), 
        .Z(n5) );
  MUX2_X1 U351 ( .A(n5), .B(n4), .S(reg_read_addr_1[1]), .Z(n6) );
  MUX2_X1 U352 ( .A(n6), .B(n3), .S(reg_read_addr_1[2]), .Z(N44) );
  MUX2_X1 U353 ( .A(reg_array[97]), .B(reg_array[113]), .S(reg_read_addr_1[0]), 
        .Z(n7) );
  MUX2_X1 U354 ( .A(reg_array[65]), .B(reg_array[81]), .S(reg_read_addr_1[0]), 
        .Z(n8) );
  MUX2_X1 U355 ( .A(n8), .B(n7), .S(reg_read_addr_1[1]), .Z(n9) );
  MUX2_X1 U356 ( .A(reg_array[33]), .B(reg_array[49]), .S(reg_read_addr_1[0]), 
        .Z(n10) );
  MUX2_X1 U357 ( .A(reg_array[1]), .B(reg_array[17]), .S(reg_read_addr_1[0]), 
        .Z(n11) );
  MUX2_X1 U358 ( .A(n11), .B(n10), .S(reg_read_addr_1[1]), .Z(n12) );
  MUX2_X1 U359 ( .A(n12), .B(n9), .S(reg_read_addr_1[2]), .Z(N43) );
  MUX2_X1 U360 ( .A(reg_array[98]), .B(reg_array[114]), .S(reg_read_addr_1[0]), 
        .Z(n13) );
  MUX2_X1 U361 ( .A(reg_array[66]), .B(reg_array[82]), .S(reg_read_addr_1[0]), 
        .Z(n1410) );
  MUX2_X1 U362 ( .A(n1410), .B(n13), .S(reg_read_addr_1[1]), .Z(n1510) );
  MUX2_X1 U363 ( .A(reg_array[34]), .B(reg_array[50]), .S(reg_read_addr_1[0]), 
        .Z(n1610) );
  MUX2_X1 U364 ( .A(reg_array[2]), .B(reg_array[18]), .S(reg_read_addr_1[0]), 
        .Z(n1710) );
  MUX2_X1 U365 ( .A(n1710), .B(n1610), .S(reg_read_addr_1[1]), .Z(n1810) );
  MUX2_X1 U366 ( .A(n1810), .B(n1510), .S(reg_read_addr_1[2]), .Z(N42) );
  MUX2_X1 U367 ( .A(reg_array[99]), .B(reg_array[115]), .S(reg_read_addr_1[0]), 
        .Z(n1910) );
  MUX2_X1 U368 ( .A(reg_array[67]), .B(reg_array[83]), .S(reg_read_addr_1[0]), 
        .Z(n20) );
  MUX2_X1 U369 ( .A(n20), .B(n1910), .S(reg_read_addr_1[1]), .Z(n289) );
  MUX2_X1 U370 ( .A(reg_array[35]), .B(reg_array[51]), .S(reg_read_addr_1[0]), 
        .Z(n2901) );
  MUX2_X1 U371 ( .A(reg_array[3]), .B(reg_array[19]), .S(reg_read_addr_1[0]), 
        .Z(n291) );
  MUX2_X1 U372 ( .A(n291), .B(n2901), .S(reg_read_addr_1[1]), .Z(n292) );
  MUX2_X1 U373 ( .A(n292), .B(n289), .S(reg_read_addr_1[2]), .Z(N41) );
  MUX2_X1 U374 ( .A(reg_array[100]), .B(reg_array[116]), .S(reg_read_addr_1[0]), .Z(n293) );
  MUX2_X1 U375 ( .A(reg_array[68]), .B(reg_array[84]), .S(reg_read_addr_1[0]), 
        .Z(n294) );
  MUX2_X1 U376 ( .A(n294), .B(n293), .S(reg_read_addr_1[1]), .Z(n295) );
  MUX2_X1 U377 ( .A(reg_array[36]), .B(reg_array[52]), .S(reg_read_addr_1[0]), 
        .Z(n296) );
  MUX2_X1 U378 ( .A(reg_array[4]), .B(reg_array[20]), .S(reg_read_addr_1[0]), 
        .Z(n297) );
  MUX2_X1 U379 ( .A(n297), .B(n296), .S(reg_read_addr_1[1]), .Z(n298) );
  MUX2_X1 U380 ( .A(n298), .B(n295), .S(reg_read_addr_1[2]), .Z(N40) );
  MUX2_X1 U381 ( .A(reg_array[101]), .B(reg_array[117]), .S(reg_read_addr_1[0]), .Z(n299) );
  MUX2_X1 U382 ( .A(reg_array[69]), .B(reg_array[85]), .S(reg_read_addr_1[0]), 
        .Z(n3001) );
  MUX2_X1 U383 ( .A(n3001), .B(n299), .S(reg_read_addr_1[1]), .Z(n301) );
  MUX2_X1 U384 ( .A(reg_array[37]), .B(reg_array[53]), .S(reg_read_addr_1[0]), 
        .Z(n302) );
  MUX2_X1 U385 ( .A(reg_array[5]), .B(reg_array[21]), .S(reg_read_addr_1[0]), 
        .Z(n303) );
  MUX2_X1 U386 ( .A(n303), .B(n302), .S(reg_read_addr_1[1]), .Z(n304) );
  MUX2_X1 U387 ( .A(n304), .B(n301), .S(reg_read_addr_1[2]), .Z(N39) );
  MUX2_X1 U388 ( .A(reg_array[102]), .B(reg_array[118]), .S(reg_read_addr_1[0]), .Z(n305) );
  MUX2_X1 U389 ( .A(reg_array[70]), .B(reg_array[86]), .S(reg_read_addr_1[0]), 
        .Z(n306) );
  MUX2_X1 U390 ( .A(n306), .B(n305), .S(reg_read_addr_1[1]), .Z(n307) );
  MUX2_X1 U391 ( .A(reg_array[38]), .B(reg_array[54]), .S(reg_read_addr_1[0]), 
        .Z(n308) );
  MUX2_X1 U392 ( .A(reg_array[6]), .B(reg_array[22]), .S(reg_read_addr_1[0]), 
        .Z(n309) );
  MUX2_X1 U393 ( .A(n309), .B(n308), .S(reg_read_addr_1[1]), .Z(n3101) );
  MUX2_X1 U394 ( .A(n3101), .B(n307), .S(reg_read_addr_1[2]), .Z(N38) );
  MUX2_X1 U395 ( .A(reg_array[103]), .B(reg_array[119]), .S(reg_read_addr_1[0]), .Z(n311) );
  MUX2_X1 U396 ( .A(reg_array[71]), .B(reg_array[87]), .S(reg_read_addr_1[0]), 
        .Z(n312) );
  MUX2_X1 U397 ( .A(n312), .B(n311), .S(reg_read_addr_1[1]), .Z(n313) );
  MUX2_X1 U398 ( .A(reg_array[39]), .B(reg_array[55]), .S(reg_read_addr_1[0]), 
        .Z(n314) );
  MUX2_X1 U399 ( .A(reg_array[7]), .B(reg_array[23]), .S(reg_read_addr_1[0]), 
        .Z(n315) );
  MUX2_X1 U400 ( .A(n315), .B(n314), .S(reg_read_addr_1[1]), .Z(n316) );
  MUX2_X1 U401 ( .A(n316), .B(n313), .S(reg_read_addr_1[2]), .Z(N37) );
  MUX2_X1 U402 ( .A(reg_array[104]), .B(reg_array[120]), .S(reg_read_addr_1[0]), .Z(n317) );
  MUX2_X1 U403 ( .A(reg_array[72]), .B(reg_array[88]), .S(reg_read_addr_1[0]), 
        .Z(n318) );
  MUX2_X1 U404 ( .A(n318), .B(n317), .S(reg_read_addr_1[1]), .Z(n319) );
  MUX2_X1 U405 ( .A(reg_array[40]), .B(reg_array[56]), .S(reg_read_addr_1[0]), 
        .Z(n3201) );
  MUX2_X1 U406 ( .A(reg_array[8]), .B(reg_array[24]), .S(reg_read_addr_1[0]), 
        .Z(n321) );
  MUX2_X1 U407 ( .A(n321), .B(n3201), .S(reg_read_addr_1[1]), .Z(n322) );
  MUX2_X1 U408 ( .A(n322), .B(n319), .S(reg_read_addr_1[2]), .Z(N36) );
  MUX2_X1 U409 ( .A(reg_array[105]), .B(reg_array[121]), .S(reg_read_addr_1[0]), .Z(n323) );
  MUX2_X1 U410 ( .A(reg_array[73]), .B(reg_array[89]), .S(reg_read_addr_1[0]), 
        .Z(n324) );
  MUX2_X1 U411 ( .A(n324), .B(n323), .S(reg_read_addr_1[1]), .Z(n325) );
  MUX2_X1 U412 ( .A(reg_array[41]), .B(reg_array[57]), .S(reg_read_addr_1[0]), 
        .Z(n326) );
  MUX2_X1 U413 ( .A(reg_array[9]), .B(reg_array[25]), .S(reg_read_addr_1[0]), 
        .Z(n327) );
  MUX2_X1 U414 ( .A(n327), .B(n326), .S(reg_read_addr_1[1]), .Z(n328) );
  MUX2_X1 U415 ( .A(n328), .B(n325), .S(reg_read_addr_1[2]), .Z(N35) );
  MUX2_X1 U416 ( .A(reg_array[106]), .B(reg_array[122]), .S(reg_read_addr_1[0]), .Z(n329) );
  MUX2_X1 U417 ( .A(reg_array[74]), .B(reg_array[90]), .S(reg_read_addr_1[0]), 
        .Z(n3301) );
  MUX2_X1 U418 ( .A(n3301), .B(n329), .S(reg_read_addr_1[1]), .Z(n331) );
  MUX2_X1 U419 ( .A(reg_array[42]), .B(reg_array[58]), .S(reg_read_addr_1[0]), 
        .Z(n332) );
  MUX2_X1 U420 ( .A(reg_array[10]), .B(reg_array[26]), .S(reg_read_addr_1[0]), 
        .Z(n333) );
  MUX2_X1 U421 ( .A(n333), .B(n332), .S(reg_read_addr_1[1]), .Z(n334) );
  MUX2_X1 U422 ( .A(n334), .B(n331), .S(reg_read_addr_1[2]), .Z(N34) );
  MUX2_X1 U423 ( .A(reg_array[107]), .B(reg_array[123]), .S(reg_read_addr_1[0]), .Z(n335) );
  MUX2_X1 U424 ( .A(reg_array[75]), .B(reg_array[91]), .S(reg_read_addr_1[0]), 
        .Z(n336) );
  MUX2_X1 U425 ( .A(n336), .B(n335), .S(reg_read_addr_1[1]), .Z(n337) );
  MUX2_X1 U426 ( .A(reg_array[43]), .B(reg_array[59]), .S(reg_read_addr_1[0]), 
        .Z(n338) );
  MUX2_X1 U427 ( .A(reg_array[11]), .B(reg_array[27]), .S(reg_read_addr_1[0]), 
        .Z(n339) );
  MUX2_X1 U428 ( .A(n339), .B(n338), .S(reg_read_addr_1[1]), .Z(n3401) );
  MUX2_X1 U429 ( .A(n3401), .B(n337), .S(reg_read_addr_1[2]), .Z(N33) );
  MUX2_X1 U430 ( .A(reg_array[108]), .B(reg_array[124]), .S(reg_read_addr_1[0]), .Z(n341) );
  MUX2_X1 U431 ( .A(reg_array[76]), .B(reg_array[92]), .S(reg_read_addr_1[0]), 
        .Z(n342) );
  MUX2_X1 U432 ( .A(n342), .B(n341), .S(reg_read_addr_1[1]), .Z(n343) );
  MUX2_X1 U433 ( .A(reg_array[44]), .B(reg_array[60]), .S(reg_read_addr_1[0]), 
        .Z(n344) );
  MUX2_X1 U434 ( .A(reg_array[12]), .B(reg_array[28]), .S(reg_read_addr_1[0]), 
        .Z(n345) );
  MUX2_X1 U435 ( .A(n345), .B(n344), .S(reg_read_addr_1[1]), .Z(n346) );
  MUX2_X1 U436 ( .A(n346), .B(n343), .S(reg_read_addr_1[2]), .Z(N32) );
  MUX2_X1 U437 ( .A(reg_array[109]), .B(reg_array[125]), .S(reg_read_addr_1[0]), .Z(n347) );
  MUX2_X1 U438 ( .A(reg_array[77]), .B(reg_array[93]), .S(reg_read_addr_1[0]), 
        .Z(n348) );
  MUX2_X1 U439 ( .A(n348), .B(n347), .S(reg_read_addr_1[1]), .Z(n349) );
  MUX2_X1 U440 ( .A(reg_array[45]), .B(reg_array[61]), .S(reg_read_addr_1[0]), 
        .Z(n3501) );
  MUX2_X1 U441 ( .A(reg_array[13]), .B(reg_array[29]), .S(reg_read_addr_1[0]), 
        .Z(n351) );
  MUX2_X1 U442 ( .A(n351), .B(n3501), .S(reg_read_addr_1[1]), .Z(n352) );
  MUX2_X1 U443 ( .A(n352), .B(n349), .S(reg_read_addr_1[2]), .Z(N31) );
  MUX2_X1 U444 ( .A(reg_array[110]), .B(reg_array[126]), .S(reg_read_addr_1[0]), .Z(n353) );
  MUX2_X1 U445 ( .A(reg_array[78]), .B(reg_array[94]), .S(reg_read_addr_1[0]), 
        .Z(n354) );
  MUX2_X1 U446 ( .A(n354), .B(n353), .S(reg_read_addr_1[1]), .Z(n355) );
  MUX2_X1 U447 ( .A(reg_array[46]), .B(reg_array[62]), .S(reg_read_addr_1[0]), 
        .Z(n356) );
  MUX2_X1 U448 ( .A(reg_array[14]), .B(reg_array[30]), .S(reg_read_addr_1[0]), 
        .Z(n357) );
  MUX2_X1 U449 ( .A(n357), .B(n356), .S(reg_read_addr_1[1]), .Z(n358) );
  MUX2_X1 U450 ( .A(n358), .B(n355), .S(reg_read_addr_1[2]), .Z(N30) );
  MUX2_X1 U451 ( .A(reg_array[111]), .B(reg_array[127]), .S(reg_read_addr_1[0]), .Z(n359) );
  MUX2_X1 U452 ( .A(reg_array[79]), .B(reg_array[95]), .S(reg_read_addr_1[0]), 
        .Z(n3601) );
  MUX2_X1 U453 ( .A(n3601), .B(n359), .S(reg_read_addr_1[1]), .Z(n361) );
  MUX2_X1 U454 ( .A(reg_array[47]), .B(reg_array[63]), .S(reg_read_addr_1[0]), 
        .Z(n362) );
  MUX2_X1 U455 ( .A(reg_array[15]), .B(reg_array[31]), .S(reg_read_addr_1[0]), 
        .Z(n363) );
  MUX2_X1 U456 ( .A(n363), .B(n362), .S(reg_read_addr_1[1]), .Z(n364) );
  MUX2_X1 U457 ( .A(n364), .B(n361), .S(reg_read_addr_1[2]), .Z(N29) );
  MUX2_X1 U458 ( .A(reg_array[96]), .B(reg_array[112]), .S(reg_read_addr_2[0]), 
        .Z(n365) );
  MUX2_X1 U459 ( .A(reg_array[64]), .B(reg_array[80]), .S(reg_read_addr_2[0]), 
        .Z(n366) );
  MUX2_X1 U460 ( .A(n366), .B(n365), .S(reg_read_addr_2[1]), .Z(n367) );
  MUX2_X1 U461 ( .A(reg_array[32]), .B(reg_array[48]), .S(reg_read_addr_2[0]), 
        .Z(n368) );
  MUX2_X1 U462 ( .A(reg_array[0]), .B(reg_array[16]), .S(reg_read_addr_2[0]), 
        .Z(n369) );
  MUX2_X1 U463 ( .A(n369), .B(n368), .S(reg_read_addr_2[1]), .Z(n3701) );
  MUX2_X1 U464 ( .A(n3701), .B(n367), .S(reg_read_addr_2[2]), .Z(N60) );
  MUX2_X1 U465 ( .A(reg_array[97]), .B(reg_array[113]), .S(reg_read_addr_2[0]), 
        .Z(n371) );
  MUX2_X1 U466 ( .A(reg_array[65]), .B(reg_array[81]), .S(reg_read_addr_2[0]), 
        .Z(n372) );
  MUX2_X1 U467 ( .A(n372), .B(n371), .S(reg_read_addr_2[1]), .Z(n373) );
  MUX2_X1 U468 ( .A(reg_array[33]), .B(reg_array[49]), .S(reg_read_addr_2[0]), 
        .Z(n374) );
  MUX2_X1 U469 ( .A(reg_array[1]), .B(reg_array[17]), .S(reg_read_addr_2[0]), 
        .Z(n375) );
  MUX2_X1 U470 ( .A(n375), .B(n374), .S(reg_read_addr_2[1]), .Z(n376) );
  MUX2_X1 U471 ( .A(n376), .B(n373), .S(reg_read_addr_2[2]), .Z(N59) );
  MUX2_X1 U472 ( .A(reg_array[98]), .B(reg_array[114]), .S(reg_read_addr_2[0]), 
        .Z(n377) );
  MUX2_X1 U473 ( .A(reg_array[66]), .B(reg_array[82]), .S(reg_read_addr_2[0]), 
        .Z(n378) );
  MUX2_X1 U474 ( .A(n378), .B(n377), .S(reg_read_addr_2[1]), .Z(n379) );
  MUX2_X1 U475 ( .A(reg_array[34]), .B(reg_array[50]), .S(reg_read_addr_2[0]), 
        .Z(n3801) );
  MUX2_X1 U476 ( .A(reg_array[2]), .B(reg_array[18]), .S(reg_read_addr_2[0]), 
        .Z(n381) );
  MUX2_X1 U477 ( .A(n381), .B(n3801), .S(reg_read_addr_2[1]), .Z(n382) );
  MUX2_X1 U478 ( .A(n382), .B(n379), .S(reg_read_addr_2[2]), .Z(N58) );
  MUX2_X1 U479 ( .A(reg_array[99]), .B(reg_array[115]), .S(reg_read_addr_2[0]), 
        .Z(n383) );
  MUX2_X1 U480 ( .A(reg_array[67]), .B(reg_array[83]), .S(reg_read_addr_2[0]), 
        .Z(n384) );
  MUX2_X1 U481 ( .A(n384), .B(n383), .S(reg_read_addr_2[1]), .Z(n385) );
  MUX2_X1 U482 ( .A(reg_array[35]), .B(reg_array[51]), .S(reg_read_addr_2[0]), 
        .Z(n386) );
  MUX2_X1 U483 ( .A(reg_array[3]), .B(reg_array[19]), .S(reg_read_addr_2[0]), 
        .Z(n387) );
  MUX2_X1 U484 ( .A(n387), .B(n386), .S(reg_read_addr_2[1]), .Z(n388) );
  MUX2_X1 U485 ( .A(n388), .B(n385), .S(reg_read_addr_2[2]), .Z(N57) );
  MUX2_X1 U486 ( .A(reg_array[100]), .B(reg_array[116]), .S(reg_read_addr_2[0]), .Z(n389) );
  MUX2_X1 U487 ( .A(reg_array[68]), .B(reg_array[84]), .S(reg_read_addr_2[0]), 
        .Z(n3901) );
  MUX2_X1 U488 ( .A(n3901), .B(n389), .S(reg_read_addr_2[1]), .Z(n391) );
  MUX2_X1 U489 ( .A(reg_array[36]), .B(reg_array[52]), .S(reg_read_addr_2[0]), 
        .Z(n392) );
  MUX2_X1 U490 ( .A(reg_array[4]), .B(reg_array[20]), .S(reg_read_addr_2[0]), 
        .Z(n393) );
  MUX2_X1 U491 ( .A(n393), .B(n392), .S(reg_read_addr_2[1]), .Z(n394) );
  MUX2_X1 U492 ( .A(n394), .B(n391), .S(reg_read_addr_2[2]), .Z(N56) );
  MUX2_X1 U493 ( .A(reg_array[101]), .B(reg_array[117]), .S(reg_read_addr_2[0]), .Z(n395) );
  MUX2_X1 U494 ( .A(reg_array[69]), .B(reg_array[85]), .S(reg_read_addr_2[0]), 
        .Z(n396) );
  MUX2_X1 U495 ( .A(n396), .B(n395), .S(reg_read_addr_2[1]), .Z(n397) );
  MUX2_X1 U496 ( .A(reg_array[37]), .B(reg_array[53]), .S(reg_read_addr_2[0]), 
        .Z(n398) );
  MUX2_X1 U497 ( .A(reg_array[5]), .B(reg_array[21]), .S(reg_read_addr_2[0]), 
        .Z(n399) );
  MUX2_X1 U498 ( .A(n399), .B(n398), .S(reg_read_addr_2[1]), .Z(n4001) );
  MUX2_X1 U499 ( .A(n4001), .B(n397), .S(reg_read_addr_2[2]), .Z(N55) );
  MUX2_X1 U500 ( .A(reg_array[102]), .B(reg_array[118]), .S(reg_read_addr_2[0]), .Z(n401) );
  MUX2_X1 U501 ( .A(reg_array[70]), .B(reg_array[86]), .S(reg_read_addr_2[0]), 
        .Z(n402) );
  MUX2_X1 U502 ( .A(n402), .B(n401), .S(reg_read_addr_2[1]), .Z(n403) );
  MUX2_X1 U503 ( .A(reg_array[38]), .B(reg_array[54]), .S(reg_read_addr_2[0]), 
        .Z(n404) );
  MUX2_X1 U504 ( .A(reg_array[6]), .B(reg_array[22]), .S(reg_read_addr_2[0]), 
        .Z(n405) );
  MUX2_X1 U505 ( .A(n405), .B(n404), .S(reg_read_addr_2[1]), .Z(n406) );
  MUX2_X1 U506 ( .A(n406), .B(n403), .S(reg_read_addr_2[2]), .Z(N54) );
  MUX2_X1 U507 ( .A(reg_array[103]), .B(reg_array[119]), .S(reg_read_addr_2[0]), .Z(n407) );
  MUX2_X1 U508 ( .A(reg_array[71]), .B(reg_array[87]), .S(reg_read_addr_2[0]), 
        .Z(n408) );
  MUX2_X1 U509 ( .A(n408), .B(n407), .S(reg_read_addr_2[1]), .Z(n409) );
  MUX2_X1 U510 ( .A(reg_array[39]), .B(reg_array[55]), .S(reg_read_addr_2[0]), 
        .Z(n4101) );
  MUX2_X1 U511 ( .A(reg_array[7]), .B(reg_array[23]), .S(reg_read_addr_2[0]), 
        .Z(n411) );
  MUX2_X1 U512 ( .A(n411), .B(n4101), .S(reg_read_addr_2[1]), .Z(n412) );
  MUX2_X1 U513 ( .A(n412), .B(n409), .S(reg_read_addr_2[2]), .Z(N53) );
  MUX2_X1 U514 ( .A(reg_array[104]), .B(reg_array[120]), .S(reg_read_addr_2[0]), .Z(n413) );
  MUX2_X1 U515 ( .A(reg_array[72]), .B(reg_array[88]), .S(reg_read_addr_2[0]), 
        .Z(n414) );
  MUX2_X1 U516 ( .A(n414), .B(n413), .S(reg_read_addr_2[1]), .Z(n415) );
  MUX2_X1 U517 ( .A(reg_array[40]), .B(reg_array[56]), .S(reg_read_addr_2[0]), 
        .Z(n416) );
  MUX2_X1 U518 ( .A(reg_array[8]), .B(reg_array[24]), .S(reg_read_addr_2[0]), 
        .Z(n417) );
  MUX2_X1 U519 ( .A(n417), .B(n416), .S(reg_read_addr_2[1]), .Z(n418) );
  MUX2_X1 U520 ( .A(n418), .B(n415), .S(reg_read_addr_2[2]), .Z(N52) );
  MUX2_X1 U521 ( .A(reg_array[105]), .B(reg_array[121]), .S(reg_read_addr_2[0]), .Z(n419) );
  MUX2_X1 U522 ( .A(reg_array[73]), .B(reg_array[89]), .S(reg_read_addr_2[0]), 
        .Z(n4201) );
  MUX2_X1 U523 ( .A(n4201), .B(n419), .S(reg_read_addr_2[1]), .Z(n421) );
  MUX2_X1 U524 ( .A(reg_array[41]), .B(reg_array[57]), .S(reg_read_addr_2[0]), 
        .Z(n422) );
  MUX2_X1 U525 ( .A(reg_array[9]), .B(reg_array[25]), .S(reg_read_addr_2[0]), 
        .Z(n423) );
  MUX2_X1 U526 ( .A(n423), .B(n422), .S(reg_read_addr_2[1]), .Z(n424) );
  MUX2_X1 U527 ( .A(n424), .B(n421), .S(reg_read_addr_2[2]), .Z(N51) );
  MUX2_X1 U528 ( .A(reg_array[106]), .B(reg_array[122]), .S(reg_read_addr_2[0]), .Z(n425) );
  MUX2_X1 U529 ( .A(reg_array[74]), .B(reg_array[90]), .S(reg_read_addr_2[0]), 
        .Z(n426) );
  MUX2_X1 U530 ( .A(n426), .B(n425), .S(reg_read_addr_2[1]), .Z(n427) );
  MUX2_X1 U531 ( .A(reg_array[42]), .B(reg_array[58]), .S(reg_read_addr_2[0]), 
        .Z(n428) );
  MUX2_X1 U532 ( .A(reg_array[10]), .B(reg_array[26]), .S(reg_read_addr_2[0]), 
        .Z(n429) );
  MUX2_X1 U533 ( .A(n429), .B(n428), .S(reg_read_addr_2[1]), .Z(n4301) );
  MUX2_X1 U534 ( .A(n4301), .B(n427), .S(reg_read_addr_2[2]), .Z(N50) );
  MUX2_X1 U535 ( .A(reg_array[107]), .B(reg_array[123]), .S(reg_read_addr_2[0]), .Z(n431) );
  MUX2_X1 U536 ( .A(reg_array[75]), .B(reg_array[91]), .S(reg_read_addr_2[0]), 
        .Z(n432) );
  MUX2_X1 U537 ( .A(n432), .B(n431), .S(reg_read_addr_2[1]), .Z(n433) );
  MUX2_X1 U538 ( .A(reg_array[43]), .B(reg_array[59]), .S(reg_read_addr_2[0]), 
        .Z(n434) );
  MUX2_X1 U539 ( .A(reg_array[11]), .B(reg_array[27]), .S(reg_read_addr_2[0]), 
        .Z(n435) );
  MUX2_X1 U540 ( .A(n435), .B(n434), .S(reg_read_addr_2[1]), .Z(n436) );
  MUX2_X1 U541 ( .A(n436), .B(n433), .S(reg_read_addr_2[2]), .Z(N49) );
  MUX2_X1 U542 ( .A(reg_array[108]), .B(reg_array[124]), .S(reg_read_addr_2[0]), .Z(n437) );
  MUX2_X1 U543 ( .A(reg_array[76]), .B(reg_array[92]), .S(reg_read_addr_2[0]), 
        .Z(n438) );
  MUX2_X1 U544 ( .A(n438), .B(n437), .S(reg_read_addr_2[1]), .Z(n439) );
  MUX2_X1 U545 ( .A(reg_array[44]), .B(reg_array[60]), .S(reg_read_addr_2[0]), 
        .Z(n4401) );
  MUX2_X1 U546 ( .A(reg_array[12]), .B(reg_array[28]), .S(reg_read_addr_2[0]), 
        .Z(n441) );
  MUX2_X1 U547 ( .A(n441), .B(n4401), .S(reg_read_addr_2[1]), .Z(n442) );
  MUX2_X1 U548 ( .A(n442), .B(n439), .S(reg_read_addr_2[2]), .Z(N48) );
  MUX2_X1 U549 ( .A(reg_array[109]), .B(reg_array[125]), .S(reg_read_addr_2[0]), .Z(n443) );
  MUX2_X1 U550 ( .A(reg_array[77]), .B(reg_array[93]), .S(reg_read_addr_2[0]), 
        .Z(n444) );
  MUX2_X1 U551 ( .A(n444), .B(n443), .S(reg_read_addr_2[1]), .Z(n445) );
  MUX2_X1 U552 ( .A(reg_array[45]), .B(reg_array[61]), .S(reg_read_addr_2[0]), 
        .Z(n446) );
  MUX2_X1 U553 ( .A(reg_array[13]), .B(reg_array[29]), .S(reg_read_addr_2[0]), 
        .Z(n447) );
  MUX2_X1 U554 ( .A(n447), .B(n446), .S(reg_read_addr_2[1]), .Z(n448) );
  MUX2_X1 U555 ( .A(n448), .B(n445), .S(reg_read_addr_2[2]), .Z(N47) );
  MUX2_X1 U556 ( .A(reg_array[110]), .B(reg_array[126]), .S(reg_read_addr_2[0]), .Z(n449) );
  MUX2_X1 U557 ( .A(reg_array[78]), .B(reg_array[94]), .S(reg_read_addr_2[0]), 
        .Z(n4501) );
  MUX2_X1 U558 ( .A(n4501), .B(n449), .S(reg_read_addr_2[1]), .Z(n451) );
  MUX2_X1 U559 ( .A(reg_array[46]), .B(reg_array[62]), .S(reg_read_addr_2[0]), 
        .Z(n452) );
  MUX2_X1 U560 ( .A(reg_array[14]), .B(reg_array[30]), .S(reg_read_addr_2[0]), 
        .Z(n453) );
  MUX2_X1 U561 ( .A(n453), .B(n452), .S(reg_read_addr_2[1]), .Z(n454) );
  MUX2_X1 U562 ( .A(n454), .B(n451), .S(reg_read_addr_2[2]), .Z(N46) );
  MUX2_X1 U563 ( .A(reg_array[111]), .B(reg_array[127]), .S(reg_read_addr_2[0]), .Z(n455) );
  MUX2_X1 U564 ( .A(reg_array[79]), .B(reg_array[95]), .S(reg_read_addr_2[0]), 
        .Z(n456) );
  MUX2_X1 U565 ( .A(n456), .B(n455), .S(reg_read_addr_2[1]), .Z(n457) );
  MUX2_X1 U566 ( .A(reg_array[47]), .B(reg_array[63]), .S(reg_read_addr_2[0]), 
        .Z(n458) );
  MUX2_X1 U567 ( .A(reg_array[15]), .B(reg_array[31]), .S(reg_read_addr_2[0]), 
        .Z(n459) );
  MUX2_X1 U568 ( .A(n459), .B(n458), .S(reg_read_addr_2[1]), .Z(n4601) );
  MUX2_X1 U569 ( .A(n4601), .B(n457), .S(reg_read_addr_2[2]), .Z(N45) );
endmodule


module JR_Control ( alu_op, funct, JRControl );
  input [1:0] alu_op;
  input [3:0] funct;
  output JRControl;
  wire   n1, n2, n4;

  INV_X1 U1 ( .A(n4), .ZN(JRControl) );
  OR4_X1 U2 ( .A1(n1), .A2(funct[0]), .A3(funct[2]), .A4(funct[1]), .ZN(n4) );
  NAND2_X1 U3 ( .A1(n2), .A2(funct[3]), .ZN(n1) );
  NOR2_X1 U4 ( .A1(alu_op[1]), .A2(alu_op[0]), .ZN(n2) );
endmodule


module ALUControl ( ALU_Control, ALUOp, Function );
  output [2:0] ALU_Control;
  input [1:0] ALUOp;
  input [3:0] Function;
  wire   n6, n7, n1, n2, n3, n4, n5;

  NOR3_X1 U1 ( .A1(n2), .A2(ALUOp[0]), .A3(n7), .ZN(ALU_Control[1]) );
  OAI22_X1 U2 ( .A1(ALUOp[1]), .A2(n5), .B1(n7), .B2(n1), .ZN(ALU_Control[0])
         );
  INV_X1 U3 ( .A(ALUOp[0]), .ZN(n5) );
  AOI21_X1 U4 ( .B1(n4), .B2(n6), .A(ALUOp[0]), .ZN(ALU_Control[2]) );
  NAND4_X1 U5 ( .A1(Function[2]), .A2(n1), .A3(n2), .A4(n3), .ZN(n6) );
  INV_X1 U6 ( .A(ALUOp[1]), .ZN(n4) );
  OR3_X1 U7 ( .A1(Function[2]), .A2(Function[3]), .A3(ALUOp[1]), .ZN(n7) );
  INV_X1 U8 ( .A(Function[1]), .ZN(n2) );
  INV_X1 U9 ( .A(Function[0]), .ZN(n1) );
  INV_X1 U10 ( .A(Function[3]), .ZN(n3) );
endmodule


module alu_DW01_sub_0 ( A, B, CI, DIFF, CO );
  input [15:0] A;
  input [15:0] B;
  output [15:0] DIFF;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17;
  wire   [15:1] carry;

  FA_X1 U2_15 ( .A(A[15]), .B(n2), .CI(carry[15]), .S(DIFF[15]) );
  FA_X1 U2_14 ( .A(A[14]), .B(n3), .CI(carry[14]), .CO(carry[15]), .S(DIFF[14]) );
  FA_X1 U2_13 ( .A(A[13]), .B(n4), .CI(carry[13]), .CO(carry[14]), .S(DIFF[13]) );
  FA_X1 U2_12 ( .A(A[12]), .B(n5), .CI(carry[12]), .CO(carry[13]), .S(DIFF[12]) );
  FA_X1 U2_11 ( .A(A[11]), .B(n6), .CI(carry[11]), .CO(carry[12]), .S(DIFF[11]) );
  FA_X1 U2_10 ( .A(A[10]), .B(n7), .CI(carry[10]), .CO(carry[11]), .S(DIFF[10]) );
  FA_X1 U2_9 ( .A(A[9]), .B(n8), .CI(carry[9]), .CO(carry[10]), .S(DIFF[9]) );
  FA_X1 U2_8 ( .A(A[8]), .B(n9), .CI(carry[8]), .CO(carry[9]), .S(DIFF[8]) );
  FA_X1 U2_7 ( .A(A[7]), .B(n10), .CI(carry[7]), .CO(carry[8]), .S(DIFF[7]) );
  FA_X1 U2_6 ( .A(A[6]), .B(n11), .CI(carry[6]), .CO(carry[7]), .S(DIFF[6]) );
  FA_X1 U2_5 ( .A(A[5]), .B(n12), .CI(carry[5]), .CO(carry[6]), .S(DIFF[5]) );
  FA_X1 U2_4 ( .A(A[4]), .B(n13), .CI(carry[4]), .CO(carry[5]), .S(DIFF[4]) );
  FA_X1 U2_3 ( .A(A[3]), .B(n14), .CI(carry[3]), .CO(carry[4]), .S(DIFF[3]) );
  FA_X1 U2_2 ( .A(A[2]), .B(n15), .CI(carry[2]), .CO(carry[3]), .S(DIFF[2]) );
  FA_X1 U2_1 ( .A(A[1]), .B(n16), .CI(carry[1]), .CO(carry[2]), .S(DIFF[1]) );
  INV_X1 U1 ( .A(B[0]), .ZN(n17) );
  INV_X1 U2 ( .A(B[15]), .ZN(n2) );
  XNOR2_X1 U3 ( .A(n17), .B(A[0]), .ZN(DIFF[0]) );
  INV_X1 U4 ( .A(B[6]), .ZN(n11) );
  INV_X1 U5 ( .A(B[7]), .ZN(n10) );
  INV_X1 U6 ( .A(B[8]), .ZN(n9) );
  INV_X1 U7 ( .A(B[9]), .ZN(n8) );
  INV_X1 U8 ( .A(B[10]), .ZN(n7) );
  NAND2_X1 U9 ( .A1(B[0]), .A2(n1), .ZN(carry[1]) );
  INV_X1 U10 ( .A(B[1]), .ZN(n16) );
  INV_X1 U11 ( .A(B[11]), .ZN(n6) );
  INV_X1 U12 ( .A(B[2]), .ZN(n15) );
  INV_X1 U13 ( .A(B[4]), .ZN(n13) );
  INV_X1 U14 ( .A(B[12]), .ZN(n5) );
  INV_X1 U15 ( .A(B[3]), .ZN(n14) );
  INV_X1 U16 ( .A(B[5]), .ZN(n12) );
  INV_X1 U17 ( .A(B[13]), .ZN(n4) );
  INV_X1 U18 ( .A(B[14]), .ZN(n3) );
  INV_X1 U19 ( .A(A[0]), .ZN(n1) );
endmodule


module alu_DW01_add_0 ( A, B, CI, SUM, CO );
  input [15:0] A;
  input [15:0] B;
  output [15:0] SUM;
  input CI;
  output CO;
  wire   n2;
  wire   [15:2] carry;

  FA_X1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .S(SUM[15]) );
  FA_X1 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  FA_X1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  FA_X1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  FA_X1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  FA_X1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  FA_X1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  FA_X1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  FA_X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  FA_X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  FA_X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  FA_X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  FA_X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  FA_X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  FA_X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(n2), .CO(carry[2]), .S(SUM[1]) );
  XOR2_X1 U1 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
  AND2_X1 U2 ( .A1(B[0]), .A2(A[0]), .ZN(n2) );
endmodule


module alu ( a, b, alu_control, result, zero );
  input [15:0] a;
  input [15:0] b;
  input [2:0] alu_control;
  output [15:0] result;
  output zero;
  wire   n118, n119, N25, N26, N27, N28, N29, N30, N31, N32, N33, N34, N35,
         N36, N37, N38, N39, N40, N41, N42, N43, N44, N45, N46, N47, N48, N49,
         N50, N51, N52, N53, N54, N55, N56, N89, n460, n470, n480, n490, n500,
         n510, n520, n530, n540, n550, n560, n57, n58, n59, n60, n61, n62, n63,
         n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77,
         n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n1, n2, n3, n6, n7,
         n8, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23,
         n24, n250, n260, n270, n280, n290, n300, n310, n320, n330, n340, n350,
         n360, n370, n380, n390, n400, n410, n420, n430, n440, n450, n88, n890,
         n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102,
         n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113,
         n114, n115, n116, n117;

  XNOR2_X2 U61 ( .A(n116), .B(n87), .ZN(n540) );
  alu_DW01_sub_0 sub_14 ( .A(a), .B(b), .CI(1'b0), .DIFF({N56, N55, N54, N53, 
        N52, N51, N50, N49, N48, N47, N46, N45, N44, N43, N42, N41}) );
  alu_DW01_add_0 r53 ( .A(a), .B(b), .CI(1'b0), .SUM({N40, N39, N38, N37, N36, 
        N35, N34, N33, N32, N31, N30, N29, N28, N27, N26, N25}) );
  OAI221_X4 U2 ( .B1(n110), .B2(n2), .C1(n510), .C2(n95), .A(n79), .ZN(
        result[9]) );
  INV_X1 U4 ( .A(N50), .ZN(n95) );
  AOI22_X1 U5 ( .A1(b[9]), .A2(n80), .B1(N34), .B2(n540), .ZN(n79) );
  OAI21_X1 U6 ( .B1(n550), .B2(n110), .A(n2), .ZN(n80) );
  BUF_X1 U8 ( .A(n119), .Z(result[3]) );
  OAI221_X1 U9 ( .B1(n1), .B2(n113), .C1(n510), .C2(n101), .A(n75), .ZN(n119)
         );
  INV_X1 U10 ( .A(N44), .ZN(n101) );
  AOI22_X1 U11 ( .A1(b[3]), .A2(n76), .B1(N28), .B2(n540), .ZN(n75) );
  OAI221_X1 U12 ( .B1(n2), .B2(n111), .C1(n510), .C2(n97), .A(n83), .ZN(
        result[7]) );
  INV_X1 U13 ( .A(N48), .ZN(n97) );
  AOI22_X1 U14 ( .A1(b[7]), .A2(n84), .B1(N32), .B2(n540), .ZN(n83) );
  OAI21_X1 U15 ( .B1(n550), .B2(n111), .A(n3), .ZN(n84) );
  BUF_X1 U16 ( .A(n118), .Z(result[5]) );
  OAI221_X1 U17 ( .B1(n1), .B2(n112), .C1(n510), .C2(n99), .A(n71), .ZN(n118)
         );
  INV_X1 U18 ( .A(N46), .ZN(n99) );
  AOI22_X1 U19 ( .A1(b[5]), .A2(n72), .B1(N30), .B2(n540), .ZN(n71) );
  BUF_X1 U20 ( .A(n500), .Z(n3) );
  BUF_X1 U21 ( .A(n500), .Z(n2) );
  BUF_X1 U22 ( .A(n500), .Z(n1) );
  OAI21_X1 U23 ( .B1(n550), .B2(n115), .A(n3), .ZN(n61) );
  OAI21_X1 U24 ( .B1(n550), .B2(n113), .A(n2), .ZN(n76) );
  OAI21_X1 U25 ( .B1(n550), .B2(n112), .A(n2), .ZN(n72) );
  OAI21_X1 U26 ( .B1(n550), .B2(n106), .A(n2), .ZN(n66) );
  OAI221_X1 U27 ( .B1(n1), .B2(n280), .C1(n510), .C2(n102), .A(n77), .ZN(
        result[2]) );
  INV_X1 U28 ( .A(N43), .ZN(n102) );
  AOI22_X1 U29 ( .A1(b[2]), .A2(n78), .B1(N27), .B2(n540), .ZN(n77) );
  OAI21_X1 U30 ( .B1(n550), .B2(n280), .A(n2), .ZN(n78) );
  OAI221_X1 U31 ( .B1(n1), .B2(n310), .C1(n510), .C2(n100), .A(n73), .ZN(
        result[4]) );
  INV_X1 U32 ( .A(N45), .ZN(n100) );
  AOI22_X1 U33 ( .A1(b[4]), .A2(n74), .B1(N29), .B2(n540), .ZN(n73) );
  OAI21_X1 U34 ( .B1(n550), .B2(n310), .A(n2), .ZN(n74) );
  OAI221_X1 U35 ( .B1(n2), .B2(n370), .C1(n510), .C2(n96), .A(n81), .ZN(
        result[8]) );
  INV_X1 U36 ( .A(N49), .ZN(n96) );
  AOI22_X1 U37 ( .A1(b[8]), .A2(n82), .B1(N33), .B2(n540), .ZN(n81) );
  OAI21_X1 U38 ( .B1(n550), .B2(n370), .A(n3), .ZN(n82) );
  OAI221_X1 U39 ( .B1(n2), .B2(n340), .C1(n510), .C2(n98), .A(n85), .ZN(
        result[6]) );
  INV_X1 U40 ( .A(N47), .ZN(n98) );
  AOI22_X1 U41 ( .A1(b[6]), .A2(n86), .B1(N31), .B2(n540), .ZN(n85) );
  OAI21_X1 U42 ( .B1(n550), .B2(n340), .A(n3), .ZN(n86) );
  OAI221_X1 U43 ( .B1(n1), .B2(n114), .C1(n510), .C2(n103), .A(n63), .ZN(
        result[1]) );
  INV_X1 U44 ( .A(N42), .ZN(n103) );
  AOI22_X1 U45 ( .A1(b[1]), .A2(n64), .B1(N26), .B2(n540), .ZN(n63) );
  OAI21_X1 U46 ( .B1(n550), .B2(n114), .A(n2), .ZN(n64) );
  OAI221_X1 U47 ( .B1(n1), .B2(n430), .C1(n510), .C2(n92), .A(n520), .ZN(
        result[12]) );
  INV_X1 U48 ( .A(N53), .ZN(n92) );
  AOI22_X1 U49 ( .A1(b[12]), .A2(n530), .B1(N37), .B2(n540), .ZN(n520) );
  OAI21_X1 U50 ( .B1(n550), .B2(n430), .A(n3), .ZN(n530) );
  OAI221_X1 U51 ( .B1(n1), .B2(n109), .C1(n510), .C2(n93), .A(n560), .ZN(
        result[11]) );
  INV_X1 U52 ( .A(N52), .ZN(n93) );
  AOI22_X1 U53 ( .A1(b[11]), .A2(n57), .B1(N36), .B2(n540), .ZN(n560) );
  OAI21_X1 U54 ( .B1(n550), .B2(n109), .A(n3), .ZN(n57) );
  OAI221_X1 U55 ( .B1(n1), .B2(n400), .C1(n510), .C2(n94), .A(n58), .ZN(
        result[10]) );
  INV_X1 U56 ( .A(N51), .ZN(n94) );
  AOI22_X1 U57 ( .A1(b[10]), .A2(n59), .B1(N35), .B2(n540), .ZN(n58) );
  OAI21_X1 U58 ( .B1(n550), .B2(n400), .A(n3), .ZN(n59) );
  OAI221_X1 U59 ( .B1(n1), .B2(n107), .C1(n510), .C2(n90), .A(n67), .ZN(
        result[14]) );
  INV_X1 U60 ( .A(N55), .ZN(n90) );
  AOI22_X1 U62 ( .A1(b[14]), .A2(n68), .B1(N39), .B2(n540), .ZN(n67) );
  OAI21_X1 U63 ( .B1(n550), .B2(n107), .A(n2), .ZN(n68) );
  OAI221_X1 U64 ( .B1(n1), .B2(n108), .C1(n510), .C2(n91), .A(n69), .ZN(
        result[13]) );
  INV_X1 U65 ( .A(N54), .ZN(n91) );
  AOI22_X1 U66 ( .A1(b[13]), .A2(n70), .B1(N38), .B2(n540), .ZN(n69) );
  OAI21_X1 U67 ( .B1(n550), .B2(n108), .A(n2), .ZN(n70) );
  OR4_X1 U68 ( .A1(result[0]), .A2(result[10]), .A3(result[11]), .A4(
        result[12]), .ZN(n490) );
  OR4_X1 U69 ( .A1(result[13]), .A2(result[14]), .A3(result[15]), .A4(
        result[1]), .ZN(n480) );
  INV_X1 U70 ( .A(b[3]), .ZN(n290) );
  INV_X1 U71 ( .A(b[5]), .ZN(n320) );
  INV_X1 U72 ( .A(b[2]), .ZN(n270) );
  INV_X1 U73 ( .A(b[4]), .ZN(n300) );
  INV_X1 U74 ( .A(b[6]), .ZN(n330) );
  INV_X1 U75 ( .A(b[14]), .ZN(n450) );
  INV_X1 U76 ( .A(n6), .ZN(n260) );
  INV_X1 U77 ( .A(b[10]), .ZN(n390) );
  INV_X1 U78 ( .A(b[7]), .ZN(n350) );
  INV_X1 U79 ( .A(b[11]), .ZN(n410) );
  INV_X1 U80 ( .A(b[13]), .ZN(n440) );
  INV_X1 U81 ( .A(b[8]), .ZN(n360) );
  INV_X1 U82 ( .A(b[12]), .ZN(n420) );
  INV_X1 U83 ( .A(b[9]), .ZN(n380) );
  NOR2_X1 U84 ( .A1(alu_control[0]), .A2(alu_control[1]), .ZN(n87) );
  NAND2_X1 U85 ( .A1(alu_control[1]), .A2(n116), .ZN(n550) );
  NAND3_X1 U86 ( .A1(n117), .A2(n116), .A3(alu_control[0]), .ZN(n510) );
  INV_X1 U87 ( .A(alu_control[1]), .ZN(n117) );
  NOR4_X1 U88 ( .A1(n105), .A2(n116), .A3(alu_control[0]), .A4(alu_control[1]), 
        .ZN(n62) );
  INV_X1 U89 ( .A(N89), .ZN(n105) );
  INV_X1 U90 ( .A(b[15]), .ZN(n88) );
  NAND3_X1 U91 ( .A1(alu_control[1]), .A2(n116), .A3(alu_control[0]), .ZN(n500) );
  INV_X1 U92 ( .A(a[2]), .ZN(n280) );
  INV_X1 U93 ( .A(a[4]), .ZN(n310) );
  INV_X1 U94 ( .A(a[6]), .ZN(n340) );
  INV_X1 U95 ( .A(a[8]), .ZN(n370) );
  INV_X1 U96 ( .A(a[10]), .ZN(n400) );
  INV_X1 U97 ( .A(a[12]), .ZN(n430) );
  INV_X1 U98 ( .A(b[0]), .ZN(n250) );
  NOR4_X1 U99 ( .A1(n460), .A2(n470), .A3(n480), .A4(n490), .ZN(zero) );
  OR4_X1 U100 ( .A1(result[6]), .A2(result[7]), .A3(result[8]), .A4(result[9]), 
        .ZN(n460) );
  OR4_X1 U101 ( .A1(result[2]), .A2(result[3]), .A3(result[4]), .A4(result[5]), 
        .ZN(n470) );
  OAI221_X1 U102 ( .B1(n1), .B2(n106), .C1(n510), .C2(n890), .A(n65), .ZN(
        result[15]) );
  INV_X1 U103 ( .A(N56), .ZN(n890) );
  AOI22_X1 U104 ( .A1(b[15]), .A2(n66), .B1(N40), .B2(n540), .ZN(n65) );
  OAI221_X1 U105 ( .B1(n1), .B2(n115), .C1(n510), .C2(n104), .A(n60), .ZN(
        result[0]) );
  INV_X1 U106 ( .A(N41), .ZN(n104) );
  AOI221_X1 U107 ( .B1(N25), .B2(n540), .C1(b[0]), .C2(n61), .A(n62), .ZN(n60)
         );
  INV_X1 U108 ( .A(a[0]), .ZN(n115) );
  INV_X1 U109 ( .A(a[9]), .ZN(n110) );
  INV_X1 U110 ( .A(a[15]), .ZN(n106) );
  INV_X1 U111 ( .A(a[3]), .ZN(n113) );
  INV_X1 U112 ( .A(a[5]), .ZN(n112) );
  INV_X1 U113 ( .A(a[1]), .ZN(n114) );
  INV_X1 U114 ( .A(a[7]), .ZN(n111) );
  INV_X1 U115 ( .A(a[11]), .ZN(n109) );
  INV_X1 U116 ( .A(a[13]), .ZN(n108) );
  INV_X1 U117 ( .A(a[14]), .ZN(n107) );
  INV_X1 U118 ( .A(alu_control[2]), .ZN(n116) );
  NOR2_X1 U119 ( .A1(a[14]), .A2(n450), .ZN(n23) );
  NOR2_X1 U120 ( .A1(n250), .A2(a[0]), .ZN(n6) );
  AOI21_X1 U121 ( .B1(n6), .B2(n114), .A(b[1]), .ZN(n7) );
  AOI221_X1 U122 ( .B1(a[2]), .B2(n270), .C1(a[1]), .C2(n260), .A(n7), .ZN(n8)
         );
  AOI221_X1 U123 ( .B1(b[3]), .B2(n113), .C1(b[2]), .C2(n280), .A(n8), .ZN(n11) );
  AOI221_X1 U124 ( .B1(a[4]), .B2(n300), .C1(a[3]), .C2(n290), .A(n11), .ZN(
        n12) );
  AOI221_X1 U125 ( .B1(b[5]), .B2(n112), .C1(b[4]), .C2(n310), .A(n12), .ZN(
        n13) );
  AOI221_X1 U126 ( .B1(a[6]), .B2(n330), .C1(a[5]), .C2(n320), .A(n13), .ZN(
        n14) );
  AOI221_X1 U127 ( .B1(b[7]), .B2(n111), .C1(b[6]), .C2(n340), .A(n14), .ZN(
        n15) );
  AOI221_X1 U128 ( .B1(a[8]), .B2(n360), .C1(a[7]), .C2(n350), .A(n15), .ZN(
        n16) );
  AOI221_X1 U129 ( .B1(b[9]), .B2(n110), .C1(b[8]), .C2(n370), .A(n16), .ZN(
        n17) );
  AOI221_X1 U130 ( .B1(a[9]), .B2(n380), .C1(a[10]), .C2(n390), .A(n17), .ZN(
        n18) );
  AOI221_X1 U131 ( .B1(b[11]), .B2(n109), .C1(b[10]), .C2(n400), .A(n18), .ZN(
        n19) );
  AOI221_X1 U132 ( .B1(a[12]), .B2(n420), .C1(a[11]), .C2(n410), .A(n19), .ZN(
        n20) );
  AOI221_X1 U133 ( .B1(b[13]), .B2(n108), .C1(b[12]), .C2(n430), .A(n20), .ZN(
        n21) );
  AOI221_X1 U134 ( .B1(a[14]), .B2(n450), .C1(a[13]), .C2(n440), .A(n21), .ZN(
        n22) );
  OAI22_X1 U135 ( .A1(n23), .A2(n22), .B1(b[15]), .B2(n106), .ZN(n24) );
  OAI21_X1 U136 ( .B1(a[15]), .B2(n88), .A(n24), .ZN(N89) );
endmodule


module data_memory ( clk, mem_access_addr, mem_write_data, mem_write_en, 
        mem_read, mem_read_data );
  input [15:0] mem_access_addr;
  input [15:0] mem_write_data;
  output [15:0] mem_read_data;
  input clk, mem_write_en, mem_read;
  wire   N286, N287, N288, N289, N290, N291, N292, N293, N294, N295, N296,
         N297, N298, N299, N300, N301, n4357, n4358, n4359, n4360, n4361,
         n4362, n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371,
         n4372, n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381,
         n4382, n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391,
         n4392, n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401,
         n4402, n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411,
         n4412, n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421,
         n4422, n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431,
         n4432, n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441,
         n4442, n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451,
         n4452, n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461,
         n4462, n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471,
         n4472, n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481,
         n4482, n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491,
         n4492, n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501,
         n4502, n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511,
         n4512, n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521,
         n4522, n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531,
         n4532, n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541,
         n4542, n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551,
         n4552, n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561,
         n4562, n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571,
         n4572, n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581,
         n4582, n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591,
         n4592, n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601,
         n4602, n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611,
         n4612, n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621,
         n4622, n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631,
         n4632, n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641,
         n4642, n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651,
         n4652, n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661,
         n4662, n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671,
         n4672, n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681,
         n4682, n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691,
         n4692, n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701,
         n4702, n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711,
         n4712, n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721,
         n4722, n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731,
         n4732, n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741,
         n4742, n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751,
         n4752, n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761,
         n4762, n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771,
         n4772, n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781,
         n4782, n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791,
         n4792, n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801,
         n4802, n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811,
         n4812, n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821,
         n4822, n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831,
         n4832, n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841,
         n4842, n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851,
         n4852, n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861,
         n4862, n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871,
         n4872, n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881,
         n4882, n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891,
         n4892, n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901,
         n4902, n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911,
         n4912, n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921,
         n4922, n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931,
         n4932, n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941,
         n4942, n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951,
         n4952, n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961,
         n4962, n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971,
         n4972, n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981,
         n4982, n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991,
         n4992, n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001,
         n5002, n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011,
         n5012, n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021,
         n5022, n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031,
         n5032, n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041,
         n5042, n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051,
         n5052, n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061,
         n5062, n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071,
         n5072, n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081,
         n5082, n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091,
         n5092, n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101,
         n5102, n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111,
         n5112, n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121,
         n5122, n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131,
         n5132, n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141,
         n5142, n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151,
         n5152, n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161,
         n5162, n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171,
         n5172, n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181,
         n5182, n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191,
         n5192, n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201,
         n5202, n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211,
         n5212, n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221,
         n5222, n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231,
         n5232, n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241,
         n5242, n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251,
         n5252, n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261,
         n5262, n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271,
         n5272, n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281,
         n5282, n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291,
         n5292, n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301,
         n5302, n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311,
         n5312, n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321,
         n5322, n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331,
         n5332, n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341,
         n5342, n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351,
         n5352, n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361,
         n5362, n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371,
         n5372, n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381,
         n5382, n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391,
         n5392, n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401,
         n5402, n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411,
         n5412, n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421,
         n5422, n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431,
         n5432, n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441,
         n5442, n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451,
         n5452, n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461,
         n5462, n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471,
         n5472, n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481,
         n5482, n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491,
         n5492, n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501,
         n5502, n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511,
         n5512, n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521,
         n5522, n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531,
         n5532, n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541,
         n5542, n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551,
         n5552, n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561,
         n5562, n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571,
         n5572, n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581,
         n5582, n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591,
         n5592, n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601,
         n5602, n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611,
         n5612, n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621,
         n5622, n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631,
         n5632, n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641,
         n5642, n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651,
         n5652, n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661,
         n5662, n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671,
         n5672, n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681,
         n5682, n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691,
         n5692, n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701,
         n5702, n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711,
         n5712, n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721,
         n5722, n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731,
         n5732, n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741,
         n5742, n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751,
         n5752, n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761,
         n5762, n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771,
         n5772, n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781,
         n5782, n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791,
         n5792, n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801,
         n5802, n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811,
         n5812, n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821,
         n5822, n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831,
         n5832, n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841,
         n5842, n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851,
         n5852, n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861,
         n5862, n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871,
         n5872, n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881,
         n5882, n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891,
         n5892, n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901,
         n5902, n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911,
         n5912, n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921,
         n5922, n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931,
         n5932, n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941,
         n5942, n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951,
         n5952, n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961,
         n5962, n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971,
         n5972, n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981,
         n5982, n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991,
         n5992, n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001,
         n6002, n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011,
         n6012, n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021,
         n6022, n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031,
         n6032, n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041,
         n6042, n6043, n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051,
         n6052, n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061,
         n6062, n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071,
         n6072, n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081,
         n6082, n6083, n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091,
         n6092, n6093, n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101,
         n6102, n6103, n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111,
         n6112, n6113, n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121,
         n6122, n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131,
         n6132, n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141,
         n6142, n6143, n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151,
         n6152, n6153, n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161,
         n6162, n6163, n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171,
         n6172, n6173, n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181,
         n6182, n6183, n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191,
         n6192, n6193, n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201,
         n6202, n6203, n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211,
         n6212, n6213, n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221,
         n6222, n6223, n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231,
         n6232, n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241,
         n6242, n6243, n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251,
         n6252, n6253, n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261,
         n6262, n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271,
         n6272, n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281,
         n6282, n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291,
         n6292, n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301,
         n6302, n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311,
         n6312, n6313, n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321,
         n6322, n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331,
         n6332, n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341,
         n6342, n6343, n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351,
         n6352, n6353, n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361,
         n6362, n6363, n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371,
         n6372, n6373, n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381,
         n6382, n6383, n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391,
         n6392, n6393, n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401,
         n6402, n6403, n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411,
         n6412, n6413, n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421,
         n6422, n6423, n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431,
         n6432, n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441,
         n6442, n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451,
         n6452, n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461,
         n6462, n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471,
         n6472, n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481,
         n6482, n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491,
         n6492, n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501,
         n6502, n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511,
         n6512, n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521,
         n6522, n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531,
         n6532, n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541,
         n6542, n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551,
         n6552, n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561,
         n6562, n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571,
         n6572, n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581,
         n6582, n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591,
         n6592, n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601,
         n6602, n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611,
         n6612, n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621,
         n6622, n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631,
         n6632, n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641,
         n6642, n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651,
         n6652, n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661,
         n6662, n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671,
         n6672, n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681,
         n6682, n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691,
         n6692, n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701,
         n6702, n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711,
         n6712, n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721,
         n6722, n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731,
         n6732, n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741,
         n6742, n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751,
         n6752, n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761,
         n6762, n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771,
         n6772, n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781,
         n6782, n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791,
         n6792, n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801,
         n6802, n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811,
         n6812, n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821,
         n6822, n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831,
         n6832, n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841,
         n6842, n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851,
         n6852, n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861,
         n6862, n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871,
         n6872, n6873, n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881,
         n6882, n6883, n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891,
         n6892, n6893, n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901,
         n6902, n6903, n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911,
         n6912, n6913, n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921,
         n6922, n6923, n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931,
         n6932, n6933, n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941,
         n6942, n6943, n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951,
         n6952, n6953, n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961,
         n6962, n6963, n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971,
         n6972, n6973, n6974, n6975, n6976, n6977, n6978, n6979, n6980, n6981,
         n6982, n6983, n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991,
         n6992, n6993, n6994, n6995, n6996, n6997, n6998, n6999, n7000, n7001,
         n7002, n7003, n7004, n7005, n7006, n7007, n7008, n7009, n7010, n7011,
         n7012, n7013, n7014, n7015, n7016, n7017, n7018, n7019, n7020, n7021,
         n7022, n7023, n7024, n7025, n7026, n7027, n7028, n7029, n7030, n7031,
         n7032, n7033, n7034, n7035, n7036, n7037, n7038, n7039, n7040, n7041,
         n7042, n7043, n7044, n7045, n7046, n7047, n7048, n7049, n7050, n7051,
         n7052, n7053, n7054, n7055, n7056, n7057, n7058, n7059, n7060, n7061,
         n7062, n7063, n7064, n7065, n7066, n7067, n7068, n7069, n7070, n7071,
         n7072, n7073, n7074, n7075, n7076, n7077, n7078, n7079, n7080, n7081,
         n7082, n7083, n7084, n7085, n7086, n7087, n7088, n7089, n7090, n7091,
         n7092, n7093, n7094, n7095, n7096, n7097, n7098, n7099, n7100, n7101,
         n7102, n7103, n7104, n7105, n7106, n7107, n7108, n7109, n7110, n7111,
         n7112, n7113, n7114, n7115, n7116, n7117, n7118, n7119, n7120, n7121,
         n7122, n7123, n7124, n7125, n7126, n7127, n7128, n7129, n7130, n7131,
         n7132, n7133, n7134, n7135, n7136, n7137, n7138, n7139, n7140, n7141,
         n7142, n7143, n7144, n7145, n7146, n7147, n7148, n7149, n7150, n7151,
         n7152, n7153, n7154, n7155, n7156, n7157, n7158, n7159, n7160, n7161,
         n7162, n7163, n7164, n7165, n7166, n7167, n7168, n7169, n7170, n7171,
         n7172, n7173, n7174, n7175, n7176, n7177, n7178, n7179, n7180, n7181,
         n7182, n7183, n7184, n7185, n7186, n7187, n7188, n7189, n7190, n7191,
         n7192, n7193, n7194, n7195, n7196, n7197, n7198, n7199, n7200, n7201,
         n7202, n7203, n7204, n7205, n7206, n7207, n7208, n7209, n7210, n7211,
         n7212, n7213, n7214, n7215, n7216, n7217, n7218, n7219, n7220, n7221,
         n7222, n7223, n7224, n7225, n7226, n7227, n7228, n7229, n7230, n7231,
         n7232, n7233, n7234, n7235, n7236, n7237, n7238, n7239, n7240, n7241,
         n7242, n7243, n7244, n7245, n7246, n7247, n7248, n7249, n7250, n7251,
         n7252, n7253, n7254, n7255, n7256, n7257, n7258, n7259, n7260, n7261,
         n7262, n7263, n7264, n7265, n7266, n7267, n7268, n7269, n7270, n7271,
         n7272, n7273, n7274, n7275, n7276, n7277, n7278, n7279, n7280, n7281,
         n7282, n7283, n7284, n7285, n7286, n7287, n7288, n7289, n7290, n7291,
         n7292, n7293, n7294, n7295, n7296, n7297, n7298, n7299, n7300, n7301,
         n7302, n7303, n7304, n7305, n7306, n7307, n7308, n7309, n7310, n7311,
         n7312, n7313, n7314, n7315, n7316, n7317, n7318, n7319, n7320, n7321,
         n7322, n7323, n7324, n7325, n7326, n7327, n7328, n7329, n7330, n7331,
         n7332, n7333, n7334, n7335, n7336, n7337, n7338, n7339, n7340, n7341,
         n7342, n7343, n7344, n7345, n7346, n7347, n7348, n7349, n7350, n7351,
         n7352, n7353, n7354, n7355, n7356, n7357, n7358, n7359, n7360, n7361,
         n7362, n7363, n7364, n7365, n7366, n7367, n7368, n7369, n7370, n7371,
         n7372, n7373, n7374, n7375, n7376, n7377, n7378, n7379, n7380, n7381,
         n7382, n7383, n7384, n7385, n7386, n7387, n7388, n7389, n7390, n7391,
         n7392, n7393, n7394, n7395, n7396, n7397, n7398, n7399, n7400, n7401,
         n7402, n7403, n7404, n7405, n7406, n7407, n7408, n7409, n7410, n7411,
         n7412, n7413, n7414, n7415, n7416, n7417, n7418, n7419, n7420, n7421,
         n7422, n7423, n7424, n7425, n7426, n7427, n7428, n7429, n7430, n7431,
         n7432, n7433, n7434, n7435, n7436, n7437, n7438, n7439, n7440, n7441,
         n7442, n7443, n7444, n7445, n7446, n7447, n7448, n7449, n7450, n7451,
         n7452, n7453, n7454, n7455, n7456, n7457, n7458, n7459, n7460, n7461,
         n7462, n7463, n7464, n7465, n7466, n7467, n7468, n7469, n7470, n7471,
         n7472, n7473, n7474, n7475, n7476, n7477, n7478, n7479, n7480, n7481,
         n7482, n7483, n7484, n7485, n7486, n7487, n7488, n7489, n7490, n7491,
         n7492, n7493, n7494, n7495, n7496, n7497, n7498, n7499, n7500, n7501,
         n7502, n7503, n7504, n7505, n7506, n7507, n7508, n7509, n7510, n7511,
         n7512, n7513, n7514, n7515, n7516, n7517, n7518, n7519, n7520, n7521,
         n7522, n7523, n7524, n7525, n7526, n7527, n7528, n7529, n7530, n7531,
         n7532, n7533, n7534, n7535, n7536, n7537, n7538, n7539, n7540, n7541,
         n7542, n7543, n7544, n7545, n7546, n7547, n7548, n7549, n7550, n7551,
         n7552, n7553, n7554, n7555, n7556, n7557, n7558, n7559, n7560, n7561,
         n7562, n7563, n7564, n7565, n7566, n7567, n7568, n7569, n7570, n7571,
         n7572, n7573, n7574, n7575, n7576, n7577, n7578, n7579, n7580, n7581,
         n7582, n7583, n7584, n7585, n7586, n7587, n7588, n7589, n7590, n7591,
         n7592, n7593, n7594, n7595, n7596, n7597, n7598, n7599, n7600, n7601,
         n7602, n7603, n7604, n7605, n7606, n7607, n7608, n7609, n7610, n7611,
         n7612, n7613, n7614, n7615, n7616, n7617, n7618, n7619, n7620, n7621,
         n7622, n7623, n7624, n7625, n7626, n7627, n7628, n7629, n7630, n7631,
         n7632, n7633, n7634, n7635, n7636, n7637, n7638, n7639, n7640, n7641,
         n7642, n7643, n7644, n7645, n7646, n7647, n7648, n7649, n7650, n7651,
         n7652, n7653, n7654, n7655, n7656, n7657, n7658, n7659, n7660, n7661,
         n7662, n7663, n7664, n7665, n7666, n7667, n7668, n7669, n7670, n7671,
         n7672, n7673, n7674, n7675, n7676, n7677, n7678, n7679, n7680, n7681,
         n7682, n7683, n7684, n7685, n7686, n7687, n7688, n7689, n7690, n7691,
         n7692, n7693, n7694, n7695, n7696, n7697, n7698, n7699, n7700, n7701,
         n7702, n7703, n7704, n7705, n7706, n7707, n7708, n7709, n7710, n7711,
         n7712, n7713, n7714, n7715, n7716, n7717, n7718, n7719, n7720, n7721,
         n7722, n7723, n7724, n7725, n7726, n7727, n7728, n7729, n7730, n7731,
         n7732, n7733, n7734, n7735, n7736, n7737, n7738, n7739, n7740, n7741,
         n7742, n7743, n7744, n7745, n7746, n7747, n7748, n7749, n7750, n7751,
         n7752, n7753, n7754, n7755, n7756, n7757, n7758, n7759, n7760, n7761,
         n7762, n7763, n7764, n7765, n7766, n7767, n7768, n7769, n7770, n7771,
         n7772, n7773, n7774, n7775, n7776, n7777, n7778, n7779, n7780, n7781,
         n7782, n7783, n7784, n7785, n7786, n7787, n7788, n7789, n7790, n7791,
         n7792, n7793, n7794, n7795, n7796, n7797, n7798, n7799, n7800, n7801,
         n7802, n7803, n7804, n7805, n7806, n7807, n7808, n7809, n7810, n7811,
         n7812, n7813, n7814, n7815, n7816, n7817, n7818, n7819, n7820, n7821,
         n7822, n7823, n7824, n7825, n7826, n7827, n7828, n7829, n7830, n7831,
         n7832, n7833, n7834, n7835, n7836, n7837, n7838, n7839, n7840, n7841,
         n7842, n7843, n7844, n7845, n7846, n7847, n7848, n7849, n7850, n7851,
         n7852, n7853, n7854, n7855, n7856, n7857, n7858, n7859, n7860, n7861,
         n7862, n7863, n7864, n7865, n7866, n7867, n7868, n7869, n7870, n7871,
         n7872, n7873, n7874, n7875, n7876, n7877, n7878, n7879, n7880, n7881,
         n7882, n7883, n7884, n7885, n7886, n7887, n7888, n7889, n7890, n7891,
         n7892, n7893, n7894, n7895, n7896, n7897, n7898, n7899, n7900, n7901,
         n7902, n7903, n7904, n7905, n7906, n7907, n7908, n7909, n7910, n7911,
         n7912, n7913, n7914, n7915, n7916, n7917, n7918, n7919, n7920, n7921,
         n7922, n7923, n7924, n7925, n7926, n7927, n7928, n7929, n7930, n7931,
         n7932, n7933, n7934, n7935, n7936, n7937, n7938, n7939, n7940, n7941,
         n7942, n7943, n7944, n7945, n7946, n7947, n7948, n7949, n7950, n7951,
         n7952, n7953, n7954, n7955, n7956, n7957, n7958, n7959, n7960, n7961,
         n7962, n7963, n7964, n7965, n7966, n7967, n7968, n7969, n7970, n7971,
         n7972, n7973, n7974, n7975, n7976, n7977, n7978, n7979, n7980, n7981,
         n7982, n7983, n7984, n7985, n7986, n7987, n7988, n7989, n7990, n7991,
         n7992, n7993, n7994, n7995, n7996, n7997, n7998, n7999, n8000, n8001,
         n8002, n8003, n8004, n8005, n8006, n8007, n8008, n8009, n8010, n8011,
         n8012, n8013, n8014, n8015, n8016, n8017, n8018, n8019, n8020, n8021,
         n8022, n8023, n8024, n8025, n8026, n8027, n8028, n8029, n8030, n8031,
         n8032, n8033, n8034, n8035, n8036, n8037, n8038, n8039, n8040, n8041,
         n8042, n8043, n8044, n8045, n8046, n8047, n8048, n8049, n8050, n8051,
         n8052, n8053, n8054, n8055, n8056, n8057, n8058, n8059, n8060, n8061,
         n8062, n8063, n8064, n8065, n8066, n8067, n8068, n8069, n8070, n8071,
         n8072, n8073, n8074, n8075, n8076, n8077, n8078, n8079, n8080, n8081,
         n8082, n8083, n8084, n8085, n8086, n8087, n8088, n8089, n8090, n8091,
         n8092, n8093, n8094, n8095, n8096, n8097, n8098, n8099, n8100, n8101,
         n8102, n8103, n8104, n8105, n8106, n8107, n8108, n8109, n8110, n8111,
         n8112, n8113, n8114, n8115, n8116, n8117, n8118, n8119, n8120, n8121,
         n8122, n8123, n8124, n8125, n8126, n8127, n8128, n8129, n8130, n8131,
         n8132, n8133, n8134, n8135, n8136, n8137, n8138, n8139, n8140, n8141,
         n8142, n8143, n8144, n8145, n8146, n8147, n8148, n8149, n8150, n8151,
         n8152, n8153, n8154, n8155, n8156, n8157, n8158, n8159, n8160, n8161,
         n8162, n8163, n8164, n8165, n8166, n8167, n8168, n8169, n8170, n8171,
         n8172, n8173, n8174, n8175, n8176, n8177, n8178, n8179, n8180, n8181,
         n8182, n8183, n8184, n8185, n8186, n8187, n8188, n8189, n8190, n8191,
         n8192, n8193, n8194, n8195, n8196, n8197, n8198, n8199, n8200, n8201,
         n8202, n8203, n8204, n8205, n8206, n8207, n8208, n8209, n8210, n8211,
         n8212, n8213, n8214, n8215, n8216, n8217, n8218, n8219, n8220, n8221,
         n8222, n8223, n8224, n8225, n8226, n8227, n8228, n8229, n8230, n8231,
         n8232, n8233, n8234, n8235, n8236, n8237, n8238, n8239, n8240, n8241,
         n8242, n8243, n8244, n8245, n8246, n8247, n8248, n8249, n8250, n8251,
         n8252, n8253, n8254, n8255, n8256, n8257, n8258, n8259, n8260, n8261,
         n8262, n8263, n8264, n8265, n8266, n8267, n8268, n8269, n8270, n8271,
         n8272, n8273, n8274, n8275, n8276, n8277, n8278, n8279, n8280, n8281,
         n8282, n8283, n8284, n8285, n8286, n8287, n8288, n8289, n8290, n8291,
         n8292, n8293, n8294, n8295, n8296, n8297, n8298, n8299, n8300, n8301,
         n8302, n8303, n8304, n8305, n8306, n8307, n8308, n8309, n8310, n8311,
         n8312, n8313, n8314, n8315, n8316, n8317, n8318, n8319, n8320, n8321,
         n8322, n8323, n8324, n8325, n8326, n8327, n8328, n8329, n8330, n8331,
         n8332, n8333, n8334, n8335, n8336, n8337, n8338, n8339, n8340, n8341,
         n8342, n8343, n8344, n8345, n8346, n8347, n8348, n8349, n8350, n8351,
         n8352, n8353, n8354, n8355, n8356, n8357, n8358, n8359, n8360, n8361,
         n8362, n8363, n8364, n8365, n8366, n8367, n8368, n8369, n8370, n8371,
         n8372, n8373, n8374, n8375, n8376, n8377, n8378, n8379, n8380, n8381,
         n8382, n8383, n8384, n8385, n8386, n8387, n8388, n8389, n8390, n8391,
         n8392, n8393, n8394, n8395, n8396, n8397, n8398, n8399, n8400, n8401,
         n8402, n8403, n8404, n8405, n8406, n8407, n8408, n8409, n8410, n8411,
         n8412, n8413, n8414, n8415, n8416, n8417, n8418, n8419, n8420, n8421,
         n8422, n8423, n8424, n8425, n8426, n8427, n8428, n8429, n8430, n8431,
         n8432, n8433, n8434, n8435, n8436, n8437, n8438, n8439, n8440, n8441,
         n8442, n8443, n8444, n8445, n8446, n8447, n8448, n8449, n8450, n8451,
         n8452, n8453, n8454, n8455, n8456, n8457, n8458, n8459, n8460, n8461,
         n8462, n8463, n8464, n8465, n8466, n8467, n8468, n8469, n8470, n8471,
         n8472, n8473, n8474, n8475, n8476, n8477, n8478, n8479, n8480, n8481,
         n8482, n8483, n8484, n8485, n8486, n8487, n8488, n8489, n8490, n8491,
         n8492, n8493, n8494, n8495, n8496, n8497, n8498, n8499, n8500, n8501,
         n8502, n8503, n8504, n8505, n8506, n8507, n8508, n8509, n8510, n8511,
         n8512, n8513, n8514, n8515, n8516, n8517, n8518, n8519, n8520, n8521,
         n8522, n8523, n8524, n8525, n8526, n8527, n8528, n8529, n8530, n8531,
         n8532, n8533, n8534, n8535, n8536, n8537, n8538, n8539, n8540, n8541,
         n8542, n8543, n8544, n8545, n8546, n8547, n8548, n8549, n8550, n8551,
         n8552, n8553, n8554, n8555, n8556, n8557, n8558, n8559, n8560, n8561,
         n8562, n8563, n8564, n8565, n8566, n8567, n8568, n8569, n8570, n8571,
         n8572, n8573, n8574, n8575, n8576, n8577, n8578, n8579, n8580, n8581,
         n8582, n8583, n8584, n8585, n8586, n8587, n8588, n8589, n8590, n8591,
         n8592, n8593, n8594, n8595, n8596, n8597, n8598, n8599, n8600, n8601,
         n8602, n8603, n8604, n8605, n8606, n8607, n8608, n8609, n8610, n8611,
         n8612, n8613, n8614, n8615, n8616, n8617, n8618, n8619, n8620, n8621,
         n8622, n8623, n8624, n8625, n8626, n8627, n8628, n8629, n8630, n8631,
         n8632, n8633, n8634, n8635, n8636, n8637, n8638, n8639, n8640, n8641,
         n8642, n8643, n8644, n8645, n8646, n8647, n8648, n8649, n8650, n8651,
         n8652, n8653, n8654, n8655, n8656, n8657, n8658, n8659, n8660, n8661,
         n8662, n8663, n8664, n8665, n8666, n8667, n8668, n8669, n8670, n8671,
         n8672, n8673, n8674, n8675, n8676, n8677, n8678, n8679, n8680, n8681,
         n8682, n8683, n8684, n8685, n8686, n8687, n8688, n8689, n8690, n8691,
         n8692, n8693, n8694, n8695, n8696, n8697, n8698, n8699, n8700, n8701,
         n8702, n8703, n8704, n8705, n8706, n8707, n8708, n8709, n8710, n8711,
         n8712, n8713, n8714, n8715, n8716, n8717, n8718, n8719, n8720, n8721,
         n8722, n8723, n8724, n8725, n8726, n8727, n8728, n8729, n8730, n8731,
         n8732, n8733, n8734, n8735, n8736, n8737, n8738, n8739, n8740, n8741,
         n8742, n8743, n8744, n8745, n8746, n8747, n8748, n8749, n8750, n8751,
         n8752, n8753, n8754, n8755, n8756, n1, n2, n3, n4, n5, n6, n7, n8, n9,
         n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20010, n21010,
         n22010, n23010, n24010, n25010, n26010, n27010, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n20000, n201, n202, n203, n204, n205, n206, n207, n208, n209, n21000,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n22000, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n23000, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n24000, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n25000, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n26000, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n27000, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n28600, n28700,
         n28800, n28900, n29000, n29100, n29200, n29300, n29400, n29500,
         n29600, n29700, n29800, n29900, n30000, n30100, n302, n303, n304,
         n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315,
         n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326,
         n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337,
         n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348,
         n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
         n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403,
         n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
         n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
         n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
         n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
         n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
         n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634,
         n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645,
         n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656,
         n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667,
         n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678,
         n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689,
         n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700,
         n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711,
         n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722,
         n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733,
         n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744,
         n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755,
         n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766,
         n767, n768, n769, n770, n771, n772, n773, n774, n775, n776, n777,
         n778, n779, n780, n781, n782, n783, n784, n785, n786, n787, n788,
         n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, n799,
         n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810,
         n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, n821,
         n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n832,
         n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, n843,
         n844, n845, n846, n847, n848, n849, n850, n851, n852, n853, n854,
         n855, n856, n857, n858, n859, n860, n861, n862, n863, n864, n865,
         n866, n867, n868, n869, n870, n871, n872, n873, n874, n875, n876,
         n877, n878, n879, n880, n881, n882, n883, n884, n885, n886, n887,
         n888, n889, n890, n891, n892, n893, n894, n895, n896, n897, n898,
         n899, n900, n901, n902, n903, n904, n905, n906, n907, n908, n909,
         n910, n911, n912, n913, n914, n915, n916, n917, n918, n919, n920,
         n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, n931,
         n932, n933, n934, n935, n936, n937, n938, n939, n940, n941, n942,
         n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, n953,
         n954, n955, n956, n957, n958, n959, n960, n961, n962, n963, n964,
         n965, n966, n967, n968, n969, n970, n971, n972, n973, n974, n975,
         n976, n977, n978, n979, n980, n981, n982, n983, n984, n985, n986,
         n987, n988, n989, n990, n991, n992, n993, n994, n995, n996, n997,
         n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007,
         n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017,
         n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027,
         n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037,
         n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047,
         n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057,
         n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067,
         n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077,
         n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087,
         n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097,
         n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107,
         n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117,
         n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127,
         n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137,
         n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147,
         n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157,
         n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167,
         n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177,
         n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187,
         n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197,
         n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207,
         n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217,
         n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227,
         n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237,
         n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247,
         n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257,
         n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267,
         n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277,
         n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287,
         n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297,
         n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307,
         n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317,
         n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327,
         n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337,
         n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347,
         n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357,
         n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367,
         n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377,
         n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387,
         n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397,
         n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407,
         n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417,
         n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427,
         n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437,
         n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447,
         n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457,
         n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467,
         n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477,
         n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487,
         n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497,
         n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507,
         n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517,
         n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527,
         n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537,
         n1538, n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547,
         n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557,
         n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567,
         n1568, n1569, n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577,
         n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587,
         n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597,
         n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606, n1607,
         n1608, n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617,
         n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627,
         n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1637,
         n1638, n1639, n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647,
         n1648, n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657,
         n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667,
         n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677,
         n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686, n1687,
         n1688, n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697,
         n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707,
         n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717,
         n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1726, n1727,
         n1728, n1729, n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1737,
         n1738, n1739, n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747,
         n1748, n1749, n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757,
         n1758, n1759, n1760, n1761, n1762, n1763, n1764, n1765, n1766, n1767,
         n1768, n1769, n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1777,
         n1778, n1779, n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787,
         n1788, n1789, n1790, n1791, n1792, n1793, n1794, n1795, n1796, n1797,
         n1798, n1799, n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807,
         n1808, n1809, n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817,
         n1818, n1819, n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1827,
         n1828, n1829, n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837,
         n1838, n1839, n1840, n1841, n1842, n1843, n1844, n1845, n1846, n1847,
         n1848, n1849, n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857,
         n1858, n1859, n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867,
         n1868, n1869, n1870, n1871, n1872, n1873, n1874, n1875, n1876, n1877,
         n1878, n1879, n1880, n1881, n1882, n1883, n1884, n1885, n1886, n1887,
         n1888, n1889, n1890, n1891, n1892, n1893, n1894, n1895, n1896, n1897,
         n1898, n1899, n1900, n1901, n1902, n1903, n1904, n1905, n1906, n1907,
         n1908, n1909, n1910, n1911, n1912, n1913, n1914, n1915, n1916, n1917,
         n1918, n1919, n1920, n1921, n1922, n1923, n1924, n1925, n1926, n1927,
         n1928, n1929, n1930, n1931, n1932, n1933, n1934, n1935, n1936, n1937,
         n1938, n1939, n1940, n1941, n1942, n1943, n1944, n1945, n1946, n1947,
         n1948, n1949, n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1957,
         n1958, n1959, n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1967,
         n1968, n1969, n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977,
         n1978, n1979, n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987,
         n1988, n1989, n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1997,
         n1998, n1999, n20001, n2001, n2002, n2003, n2004, n2005, n2006, n2007,
         n2008, n2009, n2010, n2011, n2012, n2013, n2014, n2015, n2016, n2017,
         n2018, n2019, n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2027,
         n2028, n2029, n2030, n2031, n2032, n2033, n2034, n2035, n2036, n2037,
         n2038, n2039, n2040, n2041, n2042, n2043, n2044, n2045, n2046, n2047,
         n2048, n2049, n2050, n2051, n2052, n2053, n2054, n2055, n2056, n2057,
         n2058, n2059, n2060, n2061, n2062, n2063, n2064, n2065, n2066, n2067,
         n2068, n2069, n2070, n2071, n2072, n2073, n2074, n2075, n2076, n2077,
         n2078, n2079, n2080, n2081, n2082, n2083, n2084, n2085, n2086, n2087,
         n2088, n2089, n2090, n2091, n2092, n2093, n2094, n2095, n2096, n2097,
         n2098, n2099, n21001, n2101, n2102, n2103, n2104, n2105, n2106, n2107,
         n2108, n2109, n2110, n2111, n2112, n2113, n2114, n2115, n2116, n2117,
         n2118, n2119, n2120, n2121, n2122, n2123, n2124, n2125, n2126, n2127,
         n2128, n2129, n2130, n2131, n2132, n2133, n2134, n2135, n2136, n2137,
         n2138, n2139, n2140, n2141, n2142, n2143, n2144, n2145, n2146, n2147,
         n2148, n2149, n2150, n2151, n2152, n2153, n2154, n2155, n2156, n2157,
         n2158, n2159, n2160, n2161, n2162, n2163, n2164, n2165, n2166, n2167,
         n2168, n2169, n2170, n2171, n2172, n2173, n2174, n2175, n2176, n2177,
         n2178, n2179, n2180, n2181, n2182, n2183, n2184, n2185, n2186, n2187,
         n2188, n2189, n2190, n2191, n2192, n2193, n2194, n2195, n2196, n2197,
         n2198, n2199, n22001, n2201, n2202, n2203, n2204, n2205, n2206, n2207,
         n2208, n2209, n2210, n2211, n2212, n2213, n2214, n2215, n2216, n2217,
         n2218, n2219, n2220, n2221, n2222, n2223, n2224, n2225, n2226, n2227,
         n2228, n2229, n2230, n2231, n2232, n2233, n2234, n2235, n2236, n2237,
         n2238, n2239, n2240, n2241, n2242, n2243, n2244, n2245, n2246, n2247,
         n2248, n2249, n2250, n2251, n2252, n2253, n2254, n2255, n2256, n2257,
         n2258, n2259, n2260, n2261, n2262, n2263, n2264, n2265, n2266, n2267,
         n2268, n2269, n2270, n2271, n2272, n2273, n2274, n2275, n2276, n2277,
         n2278, n2279, n2280, n2281, n2282, n2283, n2284, n2285, n2286, n2287,
         n2288, n2289, n2290, n2291, n2292, n2293, n2294, n2295, n2296, n2297,
         n2298, n2299, n23001, n2301, n2302, n2303, n2304, n2305, n2306, n2307,
         n2308, n2309, n2310, n2311, n2312, n2313, n2314, n2315, n2316, n2317,
         n2318, n2319, n2320, n2321, n2322, n2323, n2324, n2325, n2326, n2327,
         n2328, n2329, n2330, n2331, n2332, n2333, n2334, n2335, n2336, n2337,
         n2338, n2339, n2340, n2341, n2342, n2343, n2344, n2345, n2346, n2347,
         n2348, n2349, n2350, n2351, n2352, n2353, n2354, n2355, n2356, n2357,
         n2358, n2359, n2360, n2361, n2362, n2363, n2364, n2365, n2366, n2367,
         n2368, n2369, n2370, n2371, n2372, n2373, n2374, n2375, n2376, n2377,
         n2378, n2379, n2380, n2381, n2382, n2383, n2384, n2385, n2386, n2387,
         n2388, n2389, n2390, n2391, n2392, n2393, n2394, n2395, n2396, n2397,
         n2398, n2399, n24001, n2401, n2402, n2403, n2404, n2405, n2406, n2407,
         n2408, n2409, n2410, n2411, n2412, n2413, n2414, n2415, n2416, n2417,
         n2418, n2419, n2420, n2421, n2422, n2423, n2424, n2425, n2426, n2427,
         n2428, n2429, n2430, n2431, n2432, n2433, n2434, n2435, n2436, n2437,
         n2438, n2439, n2440, n2441, n2442, n2443, n2444, n2445, n2446, n2447,
         n2448, n2449, n2450, n2451, n2452, n2453, n2454, n2455, n2456, n2457,
         n2458, n2459, n2460, n2461, n2462, n2463, n2464, n2465, n2466, n2467,
         n2468, n2469, n2470, n2471, n2472, n2473, n2474, n2475, n2476, n2477,
         n2478, n2479, n2480, n2481, n2482, n2483, n2484, n2485, n2486, n2487,
         n2488, n2489, n2490, n2491, n2492, n2493, n2494, n2495, n2496, n2497,
         n2498, n2499, n25001, n2501, n2502, n2503, n2504, n2505, n2506, n2507,
         n2508, n2509, n2510, n2511, n2512, n2513, n2514, n2515, n2516, n2517,
         n2518, n2519, n2520, n2521, n2522, n2523, n2524, n2525, n2526, n2527,
         n2528, n2529, n2530, n2531, n2532, n2533, n2534, n2535, n2536, n2537,
         n2538, n2539, n2540, n2541, n2542, n2543, n2544, n2545, n2546, n2547,
         n2548, n2549, n2550, n2551, n2552, n2553, n2554, n2555, n2556, n2557,
         n2558, n2559, n2560, n2561, n2562, n2563, n2564, n2565, n2566, n2567,
         n2568, n2569, n2570, n2571, n2572, n2573, n2574, n2575, n2576, n2577,
         n2578, n2579, n2580, n2581, n2582, n2583, n2584, n2585, n2586, n2587,
         n2588, n2589, n2590, n2591, n2592, n2593, n2594, n2595, n2596, n2597,
         n2598, n2599, n26001, n2601, n2602, n2603, n2604, n2605, n2606, n2607,
         n2608, n2609, n2610, n2611, n2612, n2613, n2614, n2615, n2616, n2617,
         n2618, n2619, n2620, n2621, n2622, n2623, n2624, n2625, n2626, n2627,
         n2628, n2629, n2630, n2631, n2632, n2633, n2634, n2635, n2636, n2637,
         n2638, n2639, n2640, n2641, n2642, n2643, n2644, n2645, n2646, n2647,
         n2648, n2649, n2650, n2651, n2652, n2653, n2654, n2655, n2656, n2657,
         n2658, n2659, n2660, n2661, n2662, n2663, n2664, n2665, n2666, n2667,
         n2668, n2669, n2670, n2671, n2672, n2673, n2674, n2675, n2676, n2677,
         n2678, n2679, n2680, n2681, n2682, n2683, n2684, n2685, n2686, n2687,
         n2688, n2689, n2690, n2691, n2692, n2693, n2694, n2695, n2696, n2697,
         n2698, n2699, n27001, n2701, n2702, n2703, n2704, n2705, n2706, n2707,
         n2708, n2709, n2710, n2711, n2712, n2713, n2714, n2715, n2716, n2717,
         n2718, n2719, n2720, n2721, n2722, n2723, n2724, n2725, n2726, n2727,
         n2728, n2729, n2730, n2731, n2732, n2733, n2734, n2735, n2736, n2737,
         n2738, n2739, n2740, n2741, n2742, n2743, n2744, n2745, n2746, n2747,
         n2748, n2749, n2750, n2751, n2752, n2753, n2754, n2755, n2756, n2757,
         n2758, n2759, n2760, n2761, n2762, n2763, n2764, n2765, n2766, n2767,
         n2768, n2769, n2770, n2771, n2772, n2773, n2774, n2775, n2776, n2777,
         n2778, n2779, n2780, n2781, n2782, n2783, n2784, n2785, n2786, n2787,
         n2788, n2789, n2790, n2791, n2792, n2793, n2794, n2795, n2796, n2797,
         n2798, n2799, n2800, n2801, n2802, n2803, n2804, n2805, n2806, n2807,
         n2808, n2809, n2810, n2811, n2812, n2813, n2814, n2815, n2816, n2817,
         n2818, n2819, n2820, n2821, n2822, n2823, n2824, n2825, n2826, n2827,
         n2828, n2829, n2830, n2831, n2832, n2833, n2834, n2835, n2836, n2837,
         n2838, n2839, n2840, n2841, n2842, n2843, n2844, n2845, n2846, n2847,
         n2848, n2849, n2850, n2851, n2852, n2853, n2854, n2855, n2856, n2857,
         n2858, n2859, n28601, n2861, n2862, n2863, n2864, n2865, n2866, n2867,
         n2868, n2869, n28701, n2871, n2872, n2873, n2874, n2875, n2876, n2877,
         n2878, n2879, n28801, n2881, n2882, n2883, n2884, n2885, n2886, n2887,
         n2888, n2889, n28901, n2891, n2892, n2893, n2894, n2895, n2896, n2897,
         n2898, n2899, n29001, n2901, n2902, n2903, n2904, n2905, n2906, n2907,
         n2908, n2909, n29101, n2911, n2912, n2913, n2914, n2915, n2916, n2917,
         n2918, n2919, n29201, n2921, n2922, n2923, n2924, n2925, n2926, n2927,
         n2928, n2929, n29301, n2931, n2932, n2933, n2934, n2935, n2936, n2937,
         n2938, n2939, n29401, n2941, n2942, n2943, n2944, n2945, n2946, n2947,
         n2948, n2949, n29501, n2951, n2952, n2953, n2954, n2955, n2956, n2957,
         n2958, n2959, n29601, n2961, n2962, n2963, n2964, n2965, n2966, n2967,
         n2968, n2969, n29701, n2971, n2972, n2973, n2974, n2975, n2976, n2977,
         n2978, n2979, n29801, n2981, n2982, n2983, n2984, n2985, n2986, n2987,
         n2988, n2989, n29901, n2991, n2992, n2993, n2994, n2995, n2996, n2997,
         n2998, n2999, n30001, n3001, n3002, n3003, n3004, n3005, n3006, n3007,
         n3008, n3009, n30101, n3011, n3012, n3013, n3014, n3015, n3016, n3017,
         n3018, n3019, n3020, n3021, n3022, n3023, n3024, n3025, n3026, n3027,
         n3028, n3029, n3030, n3031, n3032, n3033, n3034, n3035, n3036, n3037,
         n3038, n3039, n3040, n3041, n3042, n3043, n3044, n3045, n3046, n3047,
         n3048, n3049, n3050, n3051, n3052, n3053, n3054, n3055, n3056, n3057,
         n3058, n3059, n3060, n3061, n3062, n3063, n3064, n3065, n3066, n3067,
         n3068, n3069, n3070, n3071, n3072, n3073, n3074, n3075, n3076, n3077,
         n3078, n3079, n3080, n3081, n3082, n3083, n3084, n3085, n3086, n3087,
         n3088, n3089, n3090, n3091, n3092, n3093, n3094, n3095, n3096, n3097,
         n3098, n3099, n3100, n3101, n3102, n3103, n3104, n3105, n3106, n3107,
         n3108, n3109, n3110, n3111, n3112, n3113, n3114, n3115, n3116, n3117,
         n3118, n3119, n3120, n3121, n3122, n3123, n3124, n3125, n3126, n3127,
         n3128, n3129, n3130, n3131, n3132, n3133, n3134, n3135, n3136, n3137,
         n3138, n3139, n3140, n3141, n3142, n3143, n3144, n3145, n3146, n3147,
         n3148, n3149, n3150, n3151, n3152, n3153, n3154, n3155, n3156, n3157,
         n3158, n3159, n3160, n3161, n3162, n3163, n3164, n3165, n3166, n3167,
         n3168, n3169, n3170, n3171, n3172, n3173, n3174, n3175, n3176, n3177,
         n3178, n3179, n3180, n3181, n3182, n3183, n3184, n3185, n3186, n3187,
         n3188, n3189, n3190, n3191, n3192, n3193, n3194, n3195, n3196, n3197,
         n3198, n3199, n3200, n3201, n3202, n3203, n3204, n3205, n3206, n3207,
         n3208, n3209, n3210, n3211, n3212, n3213, n3214, n3215, n3216, n3217,
         n3218, n3219, n3220, n3221, n3222, n3223, n3224, n3225, n3226, n3227,
         n3228, n3229, n3230, n3231, n3232, n3233, n3234, n3235, n3236, n3237,
         n3238, n3239, n3240, n3241, n3242, n3243, n3244, n3245, n3246, n3247,
         n3248, n3249, n3250, n3251, n3252, n3253, n3254, n3255, n3256, n3257,
         n3258, n3259, n3260, n3261, n3262, n3263, n3264, n3265, n3266, n3267,
         n3268, n3269, n3270, n3271, n3272, n3273, n3274, n3275, n3276, n3277,
         n3278, n3279, n3280, n3281, n3282, n3283, n3284, n3285, n3286, n3287,
         n3288, n3289, n3290, n3291, n3292, n3293, n3294, n3295, n3296, n3297,
         n3298, n3299, n3300, n3301, n3302, n3303, n3304, n3305, n3306, n3307,
         n3308, n3309, n3310, n3311, n3312, n3313, n3314, n3315, n3316, n3317,
         n3318, n3319, n3320, n3321, n3322, n3323, n3324, n3325, n3326, n3327,
         n3328, n3329, n3330, n3331, n3332, n3333, n3334, n3335, n3336, n3337,
         n3338, n3339, n3340, n3341, n3342, n3343, n3344, n3345, n3346, n3347,
         n3348, n3349, n3350, n3351, n3352, n3353, n3354, n3355, n3356, n3357,
         n3358, n3359, n3360, n3361, n3362, n3363, n3364, n3365, n3366, n3367,
         n3368, n3369, n3370, n3371, n3372, n3373, n3374, n3375, n3376, n3377,
         n3378, n3379, n3380, n3381, n3382, n3383, n3384, n3385, n3386, n3387,
         n3388, n3389, n3390, n3391, n3392, n3393, n3394, n3395, n3396, n3397,
         n3398, n3399, n3400, n3401, n3402, n3403, n3404, n3405, n3406, n3407,
         n3408, n3409, n3410, n3411, n3412, n3413, n3414, n3415, n3416, n3417,
         n3418, n3419, n3420, n3421, n3422, n3423, n3424, n3425, n3426, n3427,
         n3428, n3429, n3430, n3431, n3432, n3433, n3434, n3435, n3436, n3437,
         n3438, n3439, n3440, n3441, n3442, n3443, n3444, n3445, n3446, n3447,
         n3448, n3449, n3450, n3451, n3452, n3453, n3454, n3455, n3456, n3457,
         n3458, n3459, n3460, n3461, n3462, n3463, n3464, n3465, n3466, n3467,
         n3468, n3469, n3470, n3471, n3472, n3473, n3474, n3475, n3476, n3477,
         n3478, n3479, n3480, n3481, n3482, n3483, n3484, n3485, n3486, n3487,
         n3488, n3489, n3490, n3491, n3492, n3493, n3494, n3495, n3496, n3497,
         n3498, n3499, n3500, n3501, n3502, n3503, n3504, n3505, n3506, n3507,
         n3508, n3509, n3510, n3511, n3512, n3513, n3514, n3515, n3516, n3517,
         n3518, n3519, n3520, n3521, n3522, n3523, n3524, n3525, n3526, n3527,
         n3528, n3529, n3530, n3531, n3532, n3533, n3534, n3535, n3536, n3537,
         n3538, n3539, n3540, n3541, n3542, n3543, n3544, n3545, n3546, n3547,
         n3548, n3549, n3550, n3551, n3552, n3553, n3554, n3555, n3556, n3557,
         n3558, n3559, n3560, n3561, n3562, n3563, n3564, n3565, n3566, n3567,
         n3568, n3569, n3570, n3571, n3572, n3573, n3574, n3575, n3576, n3577,
         n3578, n3579, n3580, n3581, n3582, n3583, n3584, n3585, n3586, n3587,
         n3588, n3589, n3590, n3591, n3592, n3593, n3594, n3595, n3596, n3597,
         n3598, n3599, n3600, n3601, n3602, n3603, n3604, n3605, n3606, n3607,
         n3608, n3609, n3610, n3611, n3612, n3613, n3614, n3615, n3616, n3617,
         n3618, n3619, n3620, n3621, n3622, n3623, n3624, n3625, n3626, n3627,
         n3628, n3629, n3630, n3631, n3632, n3633, n3634, n3635, n3636, n3637,
         n3638, n3639, n3640, n3641, n3642, n3643, n3644, n3645, n3646, n3647,
         n3648, n3649, n3650, n3651, n3652, n3653, n3654, n3655, n3656, n3657,
         n3658, n3659, n3660, n3661, n3662, n3663, n3664, n3665, n3666, n3667,
         n3668, n3669, n3670, n3671, n3672, n3673, n3674, n3675, n3676, n3677,
         n3678, n3679, n3680, n3681, n3682, n3683, n3684, n3685, n3686, n3687,
         n3688, n3689, n3690, n3691, n3692, n3693, n3694, n3695, n3696, n3697,
         n3698, n3699, n3700, n3701, n3702, n3703, n3704, n3705, n3706, n3707,
         n3708, n3709, n3710, n3711, n3712, n3713, n3714, n3715, n3716, n3717,
         n3718, n3719, n3720, n3721, n3722, n3723, n3724, n3725, n3726, n3727,
         n3728, n3729, n3730, n3731, n3732, n3733, n3734, n3735, n3736, n3737,
         n3738, n3739, n3740, n3741, n3742, n3743, n3744, n3745, n3746, n3747,
         n3748, n3749, n3750, n3751, n3752, n3753, n3754, n3755, n3756, n3757,
         n3758, n3759, n3760, n3761, n3762, n3763, n3764, n3765, n3766, n3767,
         n3768, n3769, n3770, n3771, n3772, n3773, n3774, n3775, n3776, n3777,
         n3778, n3779, n3780, n3781, n3782, n3783, n3784, n3785, n3786, n3787,
         n3788, n3789, n3790, n3791, n3792, n3793, n3794, n3795, n3796, n3797,
         n3798, n3799, n3800, n3801, n3802, n3803, n3804, n3805, n3806, n3807,
         n3808, n3809, n3810, n3811, n3812, n3813, n3814, n3815, n3816, n3817,
         n3818, n3819, n3820, n3821, n3822, n3823, n3824, n3825, n3826, n3827,
         n3828, n3829, n3830, n3831, n3832, n3833, n3834, n3835, n3836, n3837,
         n3838, n3839, n3840, n3841, n3842, n3843, n3844, n3845, n3846, n3847,
         n3848, n3849, n3850, n3851, n3852, n3853, n3854, n3855, n3856, n3857,
         n3858, n3859, n3860, n3861, n3862, n3863, n3864, n3865, n3866, n3867,
         n3868, n3869, n3870, n3871, n3872, n3873, n3874, n3875, n3876, n3877,
         n3878, n3879, n3880, n3881, n3882, n3883, n3884, n3885, n3886, n3887,
         n3888, n3889, n3890, n3891, n3892, n3893, n3894, n3895, n3896, n3897,
         n3898, n3899, n3900, n3901, n3902, n3903, n3904, n3905, n3906, n3907,
         n3908, n3909, n3910, n3911, n3912, n3913, n3914, n3915, n3916, n3917,
         n3918, n3919, n3920, n3921, n3922, n3923, n3924, n3925, n3926, n3927,
         n3928, n3929, n3930, n3931, n3932, n3933, n3934, n3935, n3936, n3937,
         n3938, n3939, n3940, n3941, n3942, n3943, n3944, n3945, n3946, n3947,
         n3948, n3949, n3950, n3951, n3952, n3953, n3954, n3955, n3956, n3957,
         n3958, n3959, n3960, n3961, n3962, n3963, n3964, n3965, n3966, n3967,
         n3968, n3969, n3970, n3971, n3972, n3973, n3974, n3975, n3976, n3977,
         n3978, n3979, n3980, n3981, n3982, n3983, n3984, n3985, n3986, n3987,
         n3988, n3989, n3990, n3991, n3992, n3993, n3994, n3995, n3996, n3997,
         n3998, n3999, n4000, n4001, n4002, n4003, n4004, n4005, n4006, n4007,
         n4008, n4009, n4010, n4011, n4012, n4013, n4014, n4015, n4016, n4017,
         n4018, n4019, n4020, n4021, n4022, n4023, n4024, n4025, n4026, n4027,
         n4028, n4029, n4030, n4031, n4032, n4033, n4034, n4035, n4036, n4037,
         n4038, n4039, n4040, n4041, n4042, n4043, n4044, n4045, n4046, n4047,
         n4048, n4049, n4050, n4051, n4052, n4053, n4054, n4055, n4056, n4057,
         n4058, n4059, n4060, n4061, n4062, n4063, n4064, n4065, n4066, n4067,
         n4068, n4069, n4070, n4071, n4072, n4073, n4074, n4075, n4076, n4077,
         n4078, n4079, n4080, n4081, n4082, n4083, n4084, n4085, n4086, n4087,
         n4088, n4089, n4090, n4091, n4092, n4093, n4094, n4095, n4096, n4097,
         n4098, n4099, n4100, n4101, n4102, n4103, n4104, n4105, n4106, n4107,
         n4108, n4109, n4110, n4111, n4112, n4113, n4114, n4115, n4116, n4117,
         n4118, n4119, n4120, n4121, n4122, n4123, n4124, n4125, n4126, n4127,
         n4128, n4129, n4130, n4131, n4132, n4133, n4134, n4135, n4136, n4137,
         n4138, n4139, n4140, n4141, n4142, n4143, n4144, n4145, n4146, n4147,
         n4148, n4149, n4150, n4151, n4152, n4153, n4154, n4155, n4156, n4157,
         n4158, n4159, n4160, n4161, n4162, n4163, n4164, n4165, n4166, n4167,
         n4168, n4169, n4170, n4171, n4172, n4173, n4174, n4175, n4176, n4177,
         n4178, n4179, n4180, n4181, n4182, n4183, n4184, n4185, n4186, n4187,
         n4188, n4189, n4190, n4191, n4192, n4193, n4194, n4195, n4196, n4197,
         n4198, n4199, n4200, n4201, n4202, n4203, n4204, n4205, n4206, n4207,
         n4208, n4209, n4210, n4211, n4212, n4213, n4214, n4215, n4216, n4217,
         n4218, n4219, n4220, n4221, n4222, n4223, n4224, n4225, n4226, n4227,
         n4228, n4229, n4230, n4231, n4232, n4233, n4234, n4235, n4236, n4237,
         n4238, n4239, n4240, n4241, n4242, n4243, n4244, n4245, n4246, n4247,
         n4248, n4249, n4250, n4251, n4252, n4253, n4254, n4255, n4256, n4257,
         n4258, n4259, n4260, n4261, n4262, n4263, n4264, n4265, n4266, n4267,
         n4268, n4269, n4270, n4271, n4272, n4273, n4274, n4275, n4276, n4277,
         n4278, n4279, n4280, n4281, n4282, n4283, n4284, n4285, n4286, n4287,
         n4288, n4289, n4290, n4291, n4292, n4293, n4294, n4295, n4296, n4297,
         n4298, n4299, n4300, n4301, n4302, n4303, n4304, n4305, n4306, n4307,
         n4308, n4309, n4310, n4311, n4312, n4313, n4314, n4315, n4316, n4317,
         n4318, n4319, n4320, n4321, n4322, n4323, n4324, n4325, n4326, n4327,
         n4328, n4329, n4330, n4331, n4332, n4333, n4334, n4335, n4336, n4337,
         n4338, n4339, n4340, n4341, n4342, n4343, n4344, n4345, n4346, n4347,
         n4348, n4349, n4350, n4351, n4352, n4353, n4354, n4355, n4356, n8757,
         n8758, n8759, n8760, n8761, n8762, n8763, n8764, n8765, n8766, n8767,
         n8768, n8769, n8770, n8771, n8772, n8773, n8774, n8775, n8776, n8777,
         n8778, n8779, n8780, n8781, n8782, n8783, n8784, n8785, n8786, n8787,
         n8788, n8789, n8790, n8791, n8792, n8793, n8794, n8795, n8796, n8797,
         n8798, n8799, n8800, n8801, n8802, n8803, n8804, n8805, n8806, n8807,
         n8808, n8809, n8810, n8811, n8812, n8813, n8814, n8815, n8816, n8817,
         n8818, n8819, n8820, n8821, n8822, n8823, n8824, n8825, n8826, n8827,
         n8828, n8829, n8830, n8831, n8832, n8833, n8834, n8835, n8836, n8837,
         n8838, n8839, n8840, n8841, n8842, n8843, n8844, n8845, n8846, n8847,
         n8848, n8849, n8850, n8851, n8852, n8853, n8854, n8855, n8856, n8857,
         n8858, n8859, n8860, n8861, n8862, n8863, n8864, n8865, n8866, n8867,
         n8868, n8869, n8870, n8871, n8872, n8873, n8874, n8875, n8876, n8877,
         n8878, n8879, n8880, n8881, n8882, n8883, n8884, n8885, n8886, n8887,
         n8888, n8889, n8890, n8891, n8892, n8893, n8894, n8895, n8896, n8897,
         n8898, n8899, n8900, n8901, n8902, n8903, n8904, n8905, n8906, n8907,
         n8908, n8909, n8910, n8911, n8912, n8913, n8914, n8915, n8916, n8917,
         n8918, n8919, n8920, n8921, n8922, n8923, n8924, n8925, n8926, n8927,
         n8928, n8929, n8930, n8931, n8932, n8933, n8934, n8935, n8936, n8937,
         n8938, n8939, n8940, n8941, n8942, n8943, n8944, n8945, n8946, n8947,
         n8948, n8949, n8950, n8951, n8952, n8953, n8954, n8955, n8956, n8957,
         n8958, n8959, n8960, n8961, n8962, n8963, n8964, n8965, n8966, n8967,
         n8968, n8969, n8970, n8971, n8972, n8973, n8974, n8975, n8976, n8977,
         n8978, n8979, n8980, n8981, n8982, n8983, n8984, n8985, n8986, n8987,
         n8988, n8989, n8990, n8991, n8992, n8993, n8994, n8995, n8996, n8997,
         n8998, n8999, n9000, n9001, n9002, n9003, n9004, n9005, n9006, n9007,
         n9008, n9009, n9010, n9011, n9012, n9013, n9014, n9015, n9016, n9017,
         n9018, n9019, n9020, n9021, n9022, n9023, n9024, n9025, n9026, n9027,
         n9028, n9029, n9030, n9031, n9032, n9033, n9034, n9035, n9036, n9037,
         n9038, n9039, n9040, n9041, n9042, n9043, n9044, n9045, n9046, n9047,
         n9048, n9049, n9050, n9051, n9052, n9053, n9054, n9055, n9056, n9057,
         n9058, n9059, n9060, n9061, n9062, n9063, n9064, n9065, n9066, n9067,
         n9068, n9069, n9070, n9071, n9072, n9073, n9074, n9075, n9076, n9077,
         n9078, n9079, n9080, n9081, n9082, n9083, n9084, n9085, n9086, n9087,
         n9088, n9089, n9090, n9091, n9092, n9093, n9094, n9095, n9096, n9097,
         n9098, n9099, n9100, n9101, n9102, n9103, n9104, n9105, n9106, n9107,
         n9108, n9109, n9110, n9111, n9112, n9113, n9114, n9115, n9116, n9117,
         n9118, n9119, n9120, n9121, n9122, n9123, n9124, n9125, n9126, n9127,
         n9128, n9129, n9130, n9131, n9132, n9133, n9134, n9135, n9136, n9137,
         n9138, n9139, n9140, n9141, n9142, n9143, n9144, n9145, n9146, n9147,
         n9148, n9149, n9150, n9151, n9152, n9153, n9154, n9155, n9156, n9157,
         n9158, n9159, n9160, n9161, n9162, n9163, n9164, n9165, n9166, n9167,
         n9168, n9169, n9170, n9171, n9172, n9173, n9174, n9175, n9176, n9177,
         n9178, n9179, n9180, n9181, n9182, n9183, n9184, n9185, n9186, n9187,
         n9188, n9189, n9190, n9191, n9192, n9193, n9194, n9195, n9196, n9197,
         n9198, n9199, n9200, n9201, n9202, n9203, n9204, n9205, n9206, n9207,
         n9208, n9209, n9210, n9211, n9212, n9213, n9214, n9215, n9216, n9217,
         n9218, n9219, n9220, n9221, n9222, n9223, n9224, n9225, n9226, n9227,
         n9228, n9229, n9230, n9231, n9232, n9233, n9234, n9235, n9236, n9237,
         n9238, n9239, n9240, n9241, n9242, n9243, n9244, n9245, n9246, n9247,
         n9248, n9249, n9250, n9251, n9252, n9253, n9254, n9255, n9256, n9257,
         n9258, n9259, n9260, n9261, n9262, n9263, n9264, n9265, n9266, n9267,
         n9268, n9269, n9270, n9271, n9272, n9273, n9274, n9275, n9276, n9277,
         n9278, n9279, n9280, n9281, n9282, n9283, n9284, n9285, n9286, n9287,
         n9288, n9289, n9290, n9291, n9292, n9293, n9294, n9295, n9296, n9297,
         n9298, n9299, n9300, n9301, n9302, n9303, n9304, n9305, n9306, n9307,
         n9308, n9309, n9310, n9311, n9312, n9313, n9314, n9315, n9316, n9317,
         n9318, n9319, n9320, n9321, n9322, n9323, n9324, n9325, n9326, n9327,
         n9328, n9329, n9330, n9331, n9332, n9333, n9334, n9335, n9336, n9337,
         n9338, n9339, n9340, n9341, n9342, n9343, n9344, n9345, n9346, n9347,
         n9348, n9349, n9350, n9351, n9352, n9353, n9354, n9355, n9356, n9357,
         n9358, n9359, n9360, n9361, n9362, n9363, n9364, n9365, n9366, n9367,
         n9368, n9369, n9370, n9371, n9372, n9373, n9374, n9375, n9376, n9377,
         n9378, n9379, n9380, n9381, n9382, n9383, n9384, n9385, n9386, n9387,
         n9388, n9389, n9390, n9391, n9392, n9393, n9394, n9395, n9396, n9397,
         n9398, n9399, n9400, n9401, n9402, n9403, n9404, n9405, n9406, n9407,
         n9408, n9409, n9410, n9411, n9412, n9413, n9414, n9415, n9416, n9417,
         n9418, n9419, n9420, n9421, n9422, n9423, n9424, n9425, n9426, n9427,
         n9428, n9429, n9430, n9431, n9432, n9433, n9434, n9435, n9436, n9437,
         n9438, n9439, n9440, n9441, n9442, n9443, n9444, n9445, n9446, n9447,
         n9448, n9449, n9450, n9451, n9452, n9453, n9454, n9455, n9456, n9457,
         n9458, n9459, n9460, n9461, n9462, n9463, n9464, n9465, n9466, n9467,
         n9468, n9469, n9470, n9471, n9472, n9473, n9474, n9475, n9476, n9477,
         n9478, n9479, n9480, n9481, n9482, n9483, n9484, n9485, n9486, n9487,
         n9488, n9489, n9490, n9491, n9492, n9493, n9494, n9495, n9496, n9497,
         n9498, n9499, n9500, n9501, n9502, n9503, n9504, n9505, n9506, n9507,
         n9508, n9509, n9510, n9511, n9512, n9513, n9514, n9515, n9516, n9517,
         n9518, n9519, n9520, n9521, n9522, n9523, n9524, n9525, n9526, n9527,
         n9528, n9529, n9530, n9531, n9532, n9533, n9534, n9535, n9536, n9537,
         n9538, n9539, n9540, n9541, n9542, n9543, n9544, n9545, n9546, n9547,
         n9548, n9549, n9550, n9551, n9552, n9553, n9554, n9555, n9556, n9557,
         n9558, n9559, n9560, n9561, n9562, n9563, n9564, n9565, n9566, n9567,
         n9568, n9569, n9570, n9571, n9572, n9573, n9574, n9575, n9576, n9577,
         n9578, n9579, n9580, n9581, n9582, n9583, n9584, n9585, n9586, n9587,
         n9588, n9589, n9590, n9591, n9592, n9593, n9594, n9595, n9596, n9597,
         n9598, n9599, n9600, n9601, n9602, n9603, n9604, n9605, n9606, n9607,
         n9608, n9609, n9610, n9611, n9612, n9613, n9614, n9615, n9616, n9617,
         n9618, n9619, n9620, n9621, n9622, n9623, n9624, n9625, n9626, n9627,
         n9628, n9629, n9630, n9631, n9632, n9633, n9634, n9635, n9636, n9637,
         n9638, n9639, n9640, n9641, n9642, n9643, n9644, n9645, n9646, n9647,
         n9648, n9649, n9650, n9651, n9652, n9653, n9654, n9655, n9656, n9657,
         n9658, n9659, n9660, n9661, n9662, n9663, n9664, n9665, n9666, n9667,
         n9668, n9669, n9670, n9671, n9672, n9673, n9674, n9675, n9676, n9677,
         n9678, n9679, n9680, n9681, n9682, n9683, n9684, n9685, n9686, n9687,
         n9688, n9689, n9690, n9691, n9692, n9693, n9694, n9695, n9696, n9697,
         n9698, n9699, n9700, n9701, n9702, n9703, n9704, n9705, n9706, n9707,
         n9708, n9709, n9710, n9711, n9712, n9713, n9714, n9715, n9716, n9717,
         n9718, n9719, n9720, n9721, n9722, n9723, n9724, n9725, n9726, n9727,
         n9728, n9729, n9730, n9731, n9732, n9733, n9734, n9735, n9736, n9737,
         n9738, n9739, n9740, n9741, n9742, n9743, n9744, n9745, n9746, n9747,
         n9748, n9749, n9750, n9751, n9752, n9753, n9754, n9755, n9756, n9757,
         n9758, n9759, n9760, n9761, n9762, n9763, n9764, n9765, n9766, n9767,
         n9768, n9769, n9770, n9771, n9772, n9773, n9774, n9775, n9776, n9777,
         n9778, n9779, n9780, n9781, n9782, n9783, n9784, n9785, n9786, n9787,
         n9788, n9789, n9790, n9791, n9792, n9793, n9794, n9795, n9796, n9797,
         n9798, n9799, n9800, n9801, n9802, n9803, n9804, n9805, n9806, n9807,
         n9808, n9809, n9810, n9811, n9812, n9813, n9814, n9815, n9816, n9817,
         n9818, n9819, n9820, n9821, n9822, n9823, n9824, n9825, n9826, n9827,
         n9828, n9829, n9830, n9831, n9832, n9833, n9834, n9835, n9836, n9837,
         n9838, n9839, n9840, n9841, n9842, n9843, n9844, n9845, n9846, n9847,
         n9848, n9849, n9850, n9851, n9852, n9853, n9854, n9855, n9856, n9857,
         n9858, n9859, n9860, n9861, n9862, n9863, n9864, n9865, n9866, n9867,
         n9868, n9869, n9870, n9871, n9872, n9873, n9874, n9875, n9876, n9877,
         n9878, n9879, n9880, n9881, n9882, n9883, n9884, n9885, n9886, n9887,
         n9888, n9889, n9890, n9891, n9892, n9893, n9894, n9895, n9896, n9897,
         n9898, n9899, n9900, n9901, n9902, n9903, n9904, n9905, n9906, n9907,
         n9908, n9909, n9910, n9911, n9912, n9913, n9914, n9915, n9916, n9917,
         n9918, n9919, n9920, n9921, n9922, n9923, n9924, n9925, n9926, n9927,
         n9928, n9929, n9930, n9931, n9932, n9933, n9934, n9935, n9936, n9937,
         n9938, n9939, n9940, n9941, n9942, n9943, n9944, n9945, n9946, n9947,
         n9948, n9949, n9950, n9951, n9952, n9953, n9954, n9955, n9956, n9957,
         n9958, n9959, n9960, n9961, n9962, n9963, n9964, n9965, n9966, n9967,
         n9968, n9969, n9970, n9971, n9972, n9973, n9974, n9975, n9976, n9977,
         n9978, n9979, n9980, n9981, n9982, n9983, n9984, n9985, n9986, n9987,
         n9988, n9989, n9990, n9991, n9992, n9993, n9994, n9995, n9996, n9997,
         n9998, n9999, n10000, n10001, n10002, n10003, n10004, n10005, n10006,
         n10007, n10008, n10009, n10010, n10011, n10012, n10013, n10014,
         n10015, n10016, n10017, n10018, n10019, n10020, n10021, n10022,
         n10023, n10024, n10025, n10026, n10027, n10028, n10029, n10030,
         n10031, n10032, n10033, n10034, n10035, n10036, n10037, n10038,
         n10039, n10040, n10041, n10042, n10043, n10044, n10045, n10046,
         n10047, n10048, n10049, n10050, n10051, n10052, n10053, n10054,
         n10055, n10056, n10057, n10058, n10059, n10060, n10061, n10062,
         n10063, n10064, n10065, n10066, n10067, n10068, n10069, n10070,
         n10071, n10072, n10073, n10074, n10075, n10076, n10077, n10078,
         n10079, n10080, n10081, n10082, n10083, n10084, n10085, n10086,
         n10087, n10088, n10089, n10090, n10091, n10092, n10093, n10094,
         n10095, n10096, n10097, n10098, n10099, n10100, n10101, n10102,
         n10103, n10104, n10105, n10106, n10107, n10108, n10109, n10110,
         n10111, n10112, n10113, n10114, n10115, n10116, n10117, n10118,
         n10119, n10120, n10121, n10122, n10123, n10124, n10125, n10126,
         n10127, n10128, n10129, n10130, n10131, n10132, n10133, n10134,
         n10135, n10136, n10137, n10138, n10139, n10140, n10141, n10142,
         n10143, n10144, n10145, n10146, n10147, n10148, n10149, n10150,
         n10151, n10152, n10153, n10154, n10155, n10156, n10157, n10158,
         n10159, n10160, n10161, n10162, n10163, n10164, n10165, n10166,
         n10167, n10168, n10169, n10170, n10171, n10172, n10173, n10174,
         n10175, n10176, n10177, n10178, n10179, n10180, n10181, n10182,
         n10183, n10184, n10185, n10186, n10187, n10188, n10189, n10190,
         n10191, n10192, n10193, n10194, n10195, n10196, n10197, n10198,
         n10199, n10200, n10201, n10202, n10203, n10204, n10205, n10206,
         n10207, n10208, n10209, n10210, n10211, n10212, n10213, n10214,
         n10215, n10216, n10217, n10218, n10219, n10220, n10221, n10222,
         n10223, n10224, n10225, n10226, n10227, n10228, n10229, n10230,
         n10231, n10232, n10233, n10234, n10235, n10236, n10237, n10238,
         n10239, n10240, n10241, n10242, n10243, n10244, n10245, n10246,
         n10247, n10248, n10249, n10250, n10251, n10252, n10253, n10254,
         n10255, n10256, n10257, n10258, n10259, n10260, n10261, n10262,
         n10263, n10264, n10265, n10266, n10267, n10268, n10269, n10270,
         n10271, n10272, n10273, n10274, n10275, n10276, n10277, n10278,
         n10279, n10280, n10281, n10282, n10283, n10284, n10285, n10286,
         n10287, n10288, n10289, n10290, n10291, n10292, n10293, n10294,
         n10295, n10296, n10297, n10298, n10299, n10300, n10301, n10302,
         n10303, n10304, n10305, n10306, n10307, n10308, n10309, n10310,
         n10311, n10312, n10313, n10314, n10315, n10316, n10317, n10318,
         n10319, n10320, n10321, n10322, n10323, n10324, n10325, n10326,
         n10327, n10328, n10329, n10330, n10331, n10332, n10333, n10334,
         n10335, n10336, n10337, n10338, n10339, n10340, n10341, n10342,
         n10343, n10344, n10345, n10346, n10347, n10348, n10349, n10350,
         n10351, n10352, n10353, n10354, n10355, n10356, n10357, n10358,
         n10359, n10360, n10361, n10362, n10363, n10364, n10365, n10366,
         n10367, n10368, n10369, n10370, n10371, n10372, n10373, n10374,
         n10375, n10376, n10377, n10378, n10379, n10380, n10381, n10382,
         n10383, n10384, n10385, n10386, n10387, n10388, n10389, n10390,
         n10391, n10392, n10393, n10394, n10395, n10396, n10397, n10398,
         n10399, n10400, n10401, n10402, n10403, n10404, n10405, n10406,
         n10407, n10408, n10409, n10410, n10411, n10412, n10413, n10414,
         n10415, n10416, n10417, n10418, n10419, n10420, n10421, n10422,
         n10423, n10424, n10425, n10426, n10427, n10428, n10429, n10430,
         n10431, n10432, n10433, n10434, n10435, n10436, n10437, n10438,
         n10439, n10440, n10441, n10442, n10443, n10444, n10445, n10446,
         n10447, n10448, n10449, n10450, n10451, n10452, n10453, n10454,
         n10455, n10456, n10457, n10458, n10459, n10460, n10461, n10462,
         n10463, n10464, n10465, n10466, n10467, n10468, n10469, n10470,
         n10471, n10472, n10473, n10474, n10475, n10476, n10477, n10478,
         n10479, n10480, n10481, n10482, n10483, n10484, n10485, n10486,
         n10487, n10488, n10489, n10490, n10491, n10492, n10493, n10494,
         n10495, n10496, n10497, n10498, n10499, n10500, n10501, n10502,
         n10503, n10504, n10505, n10506, n10507, n10508, n10509, n10510,
         n10511, n10512, n10513, n10514, n10515, n10516, n10517, n10518,
         n10519, n10520, n10521, n10522, n10523, n10524, n10525, n10526,
         n10527, n10528, n10529, n10530, n10531, n10532, n10533, n10534,
         n10535, n10536, n10537, n10538, n10539, n10540, n10541, n10542,
         n10543, n10544, n10545, n10546, n10547, n10548, n10549, n10550,
         n10551, n10552, n10553, n10554, n10555, n10556, n10557, n10558,
         n10559, n10560, n10561, n10562, n10563, n10564, n10565, n10566,
         n10567, n10568, n10569, n10570, n10571, n10572, n10573, n10574,
         n10575, n10576, n10577, n10578, n10579, n10580, n10581, n10582,
         n10583, n10584, n10585, n10586, n10587, n10588, n10589, n10590,
         n10591, n10592, n10593, n10594, n10595, n10596, n10597, n10598,
         n10599, n10600, n10601, n10602, n10603, n10604, n10605, n10606,
         n10607, n10608, n10609, n10610, n10611, n10612, n10613, n10614,
         n10615, n10616, n10617, n10618, n10619, n10620, n10621, n10622,
         n10623, n10624, n10625, n10626, n10627, n10628, n10629, n10630,
         n10631, n10632, n10633, n10634, n10635, n10636, n10637, n10638,
         n10639, n10640, n10641, n10642, n10643, n10644, n10645, n10646,
         n10647, n10648, n10649, n10650, n10651, n10652, n10653, n10654,
         n10655, n10656, n10657, n10658, n10659, n10660, n10661, n10662,
         n10663, n10664, n10665, n10666, n10667, n10668, n10669, n10670,
         n10671, n10672, n10673, n10674, n10675, n10676, n10677, n10678,
         n10679, n10680, n10681, n10682, n10683, n10684, n10685, n10686,
         n10687, n10688, n10689, n10690, n10691, n10692, n10693, n10694,
         n10695, n10696, n10697, n10698, n10699, n10700, n10701, n10702,
         n10703, n10704, n10705, n10706, n10707, n10708, n10709, n10710,
         n10711, n10712, n10713, n10714, n10715, n10716, n10717, n10718,
         n10719, n10720, n10721, n10722, n10723, n10724, n10725, n10726,
         n10727, n10728, n10729, n10730, n10731, n10732, n10733, n10734,
         n10735, n10736, n10737, n10738, n10739, n10740, n10741, n10742,
         n10743, n10744, n10745, n10746, n10747, n10748, n10749, n10750,
         n10751, n10752, n10753, n10754, n10755, n10756, n10757, n10758,
         n10759, n10760, n10761, n10762, n10763, n10764, n10765, n10766,
         n10767, n10768, n10769, n10770, n10771, n10772, n10773, n10774,
         n10775, n10776, n10777, n10778, n10779, n10780, n10781, n10782,
         n10783, n10784, n10785, n10786, n10787, n10788, n10789, n10790,
         n10791, n10792, n10793, n10794, n10795, n10796, n10797, n10798,
         n10799, n10800, n10801, n10802, n10803, n10804, n10805, n10806,
         n10807, n10808, n10809, n10810, n10811, n10812, n10813, n10814,
         n10815, n10816, n10817, n10818, n10819, n10820, n10821, n10822,
         n10823, n10824, n10825, n10826, n10827, n10828, n10829, n10830,
         n10831, n10832, n10833, n10834, n10835, n10836, n10837, n10838,
         n10839, n10840, n10841, n10842, n10843, n10844, n10845, n10846,
         n10847, n10848, n10849, n10850, n10851, n10852, n10853, n10854,
         n10855, n10856, n10857, n10858, n10859, n10860, n10861, n10862,
         n10863, n10864, n10865, n10866, n10867, n10868, n10869, n10870,
         n10871, n10872, n10873, n10874, n10875, n10876, n10877, n10878,
         n10879, n10880, n10881, n10882, n10883, n10884, n10885, n10886,
         n10887, n10888, n10889, n10890, n10891, n10892, n10893, n10894,
         n10895, n10896, n10897, n10898, n10899, n10900, n10901, n10902,
         n10903, n10904, n10905, n10906, n10907, n10908, n10909, n10910,
         n10911, n10912, n10913, n10914, n10915, n10916, n10917, n10918,
         n10919, n10920, n10921, n10922, n10923, n10924, n10925, n10926,
         n10927, n10928, n10929, n10930, n10931, n10932, n10933, n10934,
         n10935, n10936, n10937, n10938, n10939, n10940, n10941, n10942,
         n10943, n10944, n10945, n10946, n10947, n10948, n10949, n10950,
         n10951, n10952, n10953, n10954, n10955, n10956, n10957, n10958,
         n10959, n10960, n10961, n10962, n10963, n10964, n10965, n10966,
         n10967, n10968, n10969, n10970, n10971, n10972, n10973, n10974,
         n10975, n10976, n10977, n10978, n10979, n10980, n10981, n10982,
         n10983, n10984, n10985, n10986, n10987, n10988, n10989, n10990,
         n10991, n10992, n10993, n10994, n10995, n10996, n10997, n10998,
         n10999, n11000, n11001, n11002, n11003, n11004, n11005, n11006,
         n11007, n11008, n11009, n11010, n11011, n11012, n11013, n11014,
         n11015, n11016, n11017, n11018, n11019, n11020, n11021, n11022,
         n11023, n11024, n11025, n11026, n11027, n11028, n11029, n11030,
         n11031, n11032, n11033, n11034, n11035, n11036, n11037, n11038,
         n11039, n11040, n11041, n11042, n11043, n11044, n11045, n11046,
         n11047, n11048, n11049, n11050, n11051, n11052, n11053, n11054,
         n11055, n11056, n11057, n11058, n11059, n11060, n11061, n11062,
         n11063, n11064, n11065, n11066, n11067, n11068, n11069, n11070,
         n11071, n11072, n11073, n11074, n11075, n11076, n11077, n11078,
         n11079, n11080, n11081, n11082, n11083, n11084, n11085, n11086,
         n11087, n11088, n11089, n11090, n11091, n11092, n11093, n11094,
         n11095, n11096, n11097, n11098, n11099, n11100, n11101, n11102,
         n11103, n11104, n11105, n11106, n11107, n11108, n11109, n11110,
         n11111, n11112, n11113, n11114, n11115, n11116, n11117, n11118,
         n11119, n11120, n11121, n11122, n11123, n11124, n11125, n11126,
         n11127, n11128, n11129, n11130, n11131, n11132, n11133, n11134,
         n11135, n11136, n11137, n11138, n11139, n11140, n11141, n11142,
         n11143, n11144, n11145, n11146, n11147, n11148, n11149, n11150,
         n11151, n11152, n11153, n11154, n11155, n11156, n11157, n11158,
         n11159, n11160, n11161, n11162, n11163, n11164, n11165, n11166,
         n11167, n11168, n11169, n11170, n11171, n11172, n11173, n11174,
         n11175, n11176, n11177, n11178, n11179, n11180, n11181, n11182,
         n11183, n11184, n11185, n11186, n11187, n11188, n11189, n11190,
         n11191, n11192, n11193, n11194, n11195, n11196, n11197, n11198,
         n11199, n11200, n11201, n11202, n11203, n11204, n11205, n11206,
         n11207, n11208, n11209, n11210, n11211, n11212, n11213, n11214,
         n11215, n11216, n11217, n11218, n11219, n11220, n11221, n11222,
         n11223, n11224, n11225, n11226, n11227, n11228, n11229, n11230,
         n11231, n11232, n11233, n11234, n11235, n11236, n11237, n11238,
         n11239, n11240, n11241, n11242, n11243, n11244, n11245, n11246,
         n11247, n11248, n11249, n11250, n11251, n11252, n11253, n11254,
         n11255, n11256, n11257, n11258, n11259, n11260, n11261, n11262,
         n11263, n11264, n11265, n11266, n11267, n11268, n11269, n11270,
         n11271, n11272, n11273, n11274, n11275, n11276, n11277, n11278,
         n11279, n11280, n11281, n11282, n11283, n11284, n11285, n11286,
         n11287, n11288, n11289, n11290, n11291, n11292, n11293, n11294,
         n11295, n11296, n11297, n11298, n11299, n11300, n11301, n11302,
         n11303, n11304, n11305, n11306, n11307, n11308, n11309, n11310,
         n11311, n11312, n11313, n11314, n11315, n11316, n11317, n11318,
         n11319, n11320, n11321, n11322, n11323, n11324, n11325, n11326,
         n11327, n11328, n11329, n11330, n11331, n11332, n11333, n11334,
         n11335, n11336, n11337, n11338, n11339, n11340, n11341, n11342,
         n11343, n11344, n11345, n11346, n11347, n11348, n11349, n11350,
         n11351, n11352, n11353, n11354, n11355, n11356, n11357, n11358,
         n11359, n11360, n11361, n11362, n11363, n11364, n11365, n11366,
         n11367, n11368, n11369, n11370, n11371, n11372, n11373, n11374,
         n11375, n11376, n11377, n11378, n11379, n11380, n11381, n11382,
         n11383, n11384, n11385, n11386, n11387, n11388, n11389, n11390,
         n11391, n11392, n11393, n11394, n11395, n11396, n11397, n11398,
         n11399, n11400, n11401, n11402, n11403, n11404, n11405, n11406,
         n11407, n11408, n11409, n11410, n11411, n11412, n11413, n11414,
         n11415, n11416, n11417, n11418, n11419, n11420, n11421, n11422,
         n11423, n11424, n11425, n11426, n11427, n11428, n11429, n11430,
         n11431, n11432, n11433, n11434, n11435, n11436, n11437, n11438,
         n11439, n11440, n11441, n11442, n11443, n11444, n11445, n11446,
         n11447, n11448, n11449, n11450, n11451, n11452, n11453, n11454,
         n11455, n11456, n11457, n11458, n11459, n11460, n11461, n11462,
         n11463, n11464, n11465, n11466, n11467, n11468, n11469, n11470,
         n11471, n11472, n11473, n11474, n11475, n11476, n11477, n11478,
         n11479, n11480, n11481, n11482, n11483, n11484, n11485, n11486,
         n11487, n11488, n11489, n11490, n11491, n11492, n11493, n11494,
         n11495, n11496, n11497, n11498, n11499, n11500, n11501, n11502,
         n11503, n11504, n11505, n11506, n11507, n11508, n11509, n11510,
         n11511, n11512, n11513, n11514, n11515, n11516, n11517, n11518,
         n11519, n11520, n11521, n11522, n11523, n11524, n11525, n11526,
         n11527, n11528, n11529, n11530, n11531, n11532, n11533, n11534,
         n11535, n11536, n11537, n11538, n11539, n11540, n11541, n11542,
         n11543, n11544, n11545, n11546, n11547, n11548, n11549, n11550,
         n11551, n11552, n11553, n11554, n11555, n11556, n11557, n11558,
         n11559, n11560, n11561, n11562, n11563, n11564, n11565, n11566,
         n11567, n11568, n11569, n11570, n11571, n11572, n11573, n11574,
         n11575, n11576, n11577, n11578, n11579, n11580, n11581, n11582,
         n11583, n11584, n11585, n11586, n11587, n11588, n11589, n11590,
         n11591, n11592, n11593, n11594, n11595, n11596, n11597, n11598,
         n11599, n11600, n11601, n11602, n11603, n11604, n11605, n11606,
         n11607, n11608, n11609, n11610, n11611, n11612, n11613, n11614,
         n11615, n11616, n11617, n11618, n11619, n11620, n11621, n11622,
         n11623, n11624, n11625, n11626, n11627, n11628, n11629, n11630,
         n11631, n11632, n11633, n11634, n11635, n11636, n11637, n11638,
         n11639, n11640, n11641, n11642, n11643, n11644, n11645, n11646,
         n11647, n11648, n11649, n11650, n11651, n11652, n11653, n11654,
         n11655, n11656, n11657, n11658, n11659, n11660, n11661, n11662,
         n11663, n11664, n11665, n11666, n11667, n11668, n11669, n11670,
         n11671, n11672, n11673, n11674, n11675, n11676, n11677, n11678,
         n11679, n11680, n11681, n11682, n11683, n11684, n11685, n11686,
         n11687, n11688, n11689, n11690, n11691, n11692, n11693, n11694,
         n11695, n11696, n11697, n11698, n11699, n11700, n11701, n11702,
         n11703, n11704, n11705, n11706, n11707, n11708, n11709, n11710,
         n11711, n11712, n11713, n11714, n11715, n11716, n11717, n11718,
         n11719, n11720, n11721, n11722, n11723, n11724, n11725, n11726,
         n11727, n11728, n11729, n11730, n11731, n11732, n11733, n11734,
         n11735, n11736, n11737, n11738, n11739, n11740, n11741, n11742,
         n11743, n11744, n11745, n11746, n11747, n11748, n11749, n11750,
         n11751, n11752, n11753, n11754, n11755, n11756, n11757, n11758,
         n11759, n11760, n11761, n11762, n11763, n11764, n11765, n11766,
         n11767, n11768, n11769, n11770, n11771, n11772, n11773, n11774,
         n11775, n11776, n11777, n11778, n11779, n11780, n11781, n11782,
         n11783, n11784, n11785, n11786, n11787, n11788, n11789, n11790,
         n11791, n11792, n11793, n11794, n11795, n11796, n11797, n11798,
         n11799, n11800, n11801, n11802, n11803, n11804, n11805, n11806,
         n11807, n11808, n11809, n11810, n11811, n11812, n11813, n11814,
         n11815, n11816, n11817, n11818, n11819, n11820, n11821, n11822,
         n11823, n11824, n11825, n11826, n11827, n11828, n11829, n11830,
         n11831, n11832, n11833, n11834, n11835, n11836, n11837, n11838,
         n11839, n11840, n11841, n11842, n11843, n11844, n11845, n11846,
         n11847, n11848, n11849, n11850, n11851, n11852, n11853, n11854,
         n11855, n11856, n11857, n11858, n11859, n11860, n11861, n11862,
         n11863, n11864, n11865, n11866, n11867, n11868, n11869, n11870,
         n11871, n11872, n11873, n11874, n11875, n11876, n11877, n11878,
         n11879, n11880, n11881, n11882, n11883, n11884, n11885, n11886,
         n11887, n11888, n11889, n11890, n11891, n11892, n11893, n11894,
         n11895, n11896, n11897, n11898, n11899, n11900, n11901, n11902,
         n11903, n11904, n11905, n11906, n11907, n11908, n11909, n11910,
         n11911, n11912, n11913, n11914, n11915, n11916, n11917, n11918,
         n11919, n11920, n11921, n11922, n11923, n11924, n11925, n11926,
         n11927, n11928, n11929, n11930, n11931, n11932, n11933, n11934,
         n11935, n11936, n11937, n11938, n11939, n11940, n11941, n11942,
         n11943, n11944, n11945, n11946, n11947, n11948, n11949, n11950,
         n11951, n11952, n11953, n11954, n11955, n11956, n11957, n11958,
         n11959, n11960, n11961, n11962, n11963, n11964, n11965, n11966,
         n11967, n11968, n11969, n11970, n11971, n11972, n11973, n11974,
         n11975, n11976, n11977, n11978, n11979, n11980, n11981, n11982,
         n11983, n11984, n11985, n11986, n11987, n11988, n11989, n11990,
         n11991, n11992, n11993, n11994, n11995, n11996, n11997, n11998,
         n11999, n12000, n12001, n12002, n12003, n12004, n12005, n12006,
         n12007, n12008, n12009, n12010, n12011, n12012, n12013, n12014,
         n12015, n12016, n12017, n12018, n12019, n12020, n12021, n12022,
         n12023, n12024, n12025, n12026, n12027, n12028, n12029, n12030,
         n12031, n12032, n12033, n12034, n12035, n12036, n12037, n12038,
         n12039, n12040, n12041, n12042, n12043, n12044, n12045, n12046,
         n12047, n12048, n12049, n12050, n12051, n12052, n12053, n12054,
         n12055, n12056, n12057, n12058, n12059, n12060, n12061, n12062,
         n12063, n12064, n12065, n12066, n12067, n12068, n12069, n12070,
         n12071, n12072, n12073, n12074, n12075, n12076, n12077, n12078,
         n12079, n12080, n12081, n12082, n12083, n12084, n12085, n12086,
         n12087, n12088, n12089, n12090, n12091, n12092, n12093, n12094,
         n12095, n12096, n12097, n12098, n12099, n12100, n12101, n12102,
         n12103, n12104, n12105, n12106, n12107, n12108, n12109, n12110,
         n12111, n12112, n12113, n12114, n12115, n12116, n12117, n12118,
         n12119, n12120, n12121, n12122, n12123, n12124, n12125, n12126,
         n12127, n12128, n12129, n12130, n12131, n12132, n12133, n12134,
         n12135, n12136, n12137, n12138, n12139, n12140, n12141, n12142,
         n12143, n12144, n12145, n12146, n12147, n12148, n12149, n12150,
         n12151, n12152, n12153, n12154, n12155, n12156, n12157, n12158,
         n12159, n12160, n12161, n12162, n12163, n12164, n12165, n12166,
         n12167, n12168, n12169, n12170, n12171, n12172, n12173, n12174,
         n12175, n12176, n12177, n12178, n12179, n12180, n12181, n12182,
         n12183, n12184, n12185, n12186, n12187, n12188, n12189, n12190,
         n12191, n12192, n12193, n12194, n12195, n12196, n12197, n12198,
         n12199, n12200, n12201, n12202, n12203, n12204, n12205, n12206,
         n12207, n12208, n12209, n12210, n12211, n12212, n12213, n12214,
         n12215, n12216, n12217, n12218, n12219, n12220, n12221, n12222,
         n12223, n12224, n12225, n12226, n12227, n12228, n12229, n12230,
         n12231, n12232, n12233, n12234, n12235, n12236, n12237, n12238,
         n12239, n12240, n12241, n12242, n12243, n12244, n12245, n12246,
         n12247, n12248, n12249, n12250, n12251, n12252, n12253, n12254,
         n12255, n12256, n12257, n12258, n12259, n12260, n12261, n12262,
         n12263, n12264, n12265, n12266, n12267, n12268, n12269, n12270,
         n12271, n12272, n12273, n12274, n12275, n12276, n12277, n12278,
         n12279, n12280, n12281, n12282, n12283, n12284, n12285, n12286,
         n12287, n12288, n12289, n12290, n12291, n12292, n12293, n12294,
         n12295, n12296, n12297, n12298, n12299, n12300, n12301, n12302,
         n12303, n12304, n12305, n12306, n12307, n12308, n12309, n12310,
         n12311, n12312, n12313, n12314, n12315, n12316, n12317, n12318,
         n12319, n12320, n12321, n12322, n12323, n12324, n12325, n12326,
         n12327, n12328, n12329, n12330, n12331, n12332, n12333, n12334,
         n12335, n12336, n12337, n12338, n12339, n12340, n12341, n12342,
         n12343, n12344, n12345, n12346, n12347, n12348, n12349, n12350,
         n12351, n12352, n12353, n12354, n12355, n12356, n12357, n12358,
         n12359, n12360, n12361, n12362, n12363, n12364, n12365, n12366,
         n12367, n12368, n12369, n12370, n12371, n12372, n12373, n12374,
         n12375, n12376, n12377, n12378, n12379, n12380, n12381, n12382,
         n12383, n12384, n12385, n12386, n12387, n12388, n12389, n12390,
         n12391, n12392, n12393, n12394, n12395, n12396, n12397, n12398,
         n12399, n12400, n12401, n12402, n12403, n12404, n12405, n12406,
         n12407, n12408, n12409, n12410, n12411, n12412, n12413, n12414,
         n12415, n12416, n12417, n12418, n12419, n12420, n12421, n12422,
         n12423, n12424, n12425, n12426, n12427, n12428, n12429, n12430,
         n12431, n12432, n12433, n12434, n12435, n12436, n12437, n12438,
         n12439, n12440, n12441, n12442, n12443, n12444, n12445, n12446,
         n12447, n12448, n12449, n12450, n12451, n12452, n12453, n12454,
         n12455, n12456, n12457, n12458, n12459, n12460, n12461, n12462,
         n12463, n12464, n12465, n12466, n12467, n12468, n12469, n12470,
         n12471, n12472, n12473, n12474, n12475, n12476, n12477, n12478,
         n12479, n12480, n12481, n12482, n12483, n12484, n12485, n12486,
         n12487, n12488, n12489, n12490, n12491, n12492, n12493, n12494,
         n12495, n12496, n12497, n12498, n12499, n12500, n12501, n12502,
         n12503, n12504, n12505, n12506, n12507, n12508, n12509, n12510,
         n12511, n12512, n12513, n12514, n12515, n12516, n12517, n12518,
         n12519, n12520, n12521, n12522, n12523, n12524, n12525, n12526,
         n12527, n12528, n12529, n12530, n12531, n12532, n12533, n12534,
         n12535, n12536, n12537, n12538, n12539, n12540, n12541, n12542,
         n12543, n12544, n12545, n12546, n12547, n12548, n12549, n12550,
         n12551, n12552, n12553, n12554, n12555, n12556, n12557, n12558,
         n12559, n12560, n12561, n12562, n12563, n12564, n12565, n12566,
         n12567, n12568, n12569, n12570, n12571, n12572, n12573, n12574,
         n12575, n12576, n12577, n12578, n12579, n12580, n12581, n12582,
         n12583, n12584, n12585, n12586, n12587, n12588, n12589, n12590,
         n12591, n12592, n12593, n12594, n12595, n12596, n12597, n12598,
         n12599, n12600, n12601, n12602, n12603, n12604, n12605, n12606,
         n12607, n12608, n12609, n12610, n12611, n12612, n12613, n12614,
         n12615, n12616, n12617, n12618, n12619, n12620, n12621, n12622,
         n12623, n12624, n12625, n12626, n12627, n12628, n12629, n12630,
         n12631, n12632, n12633, n12634, n12635, n12636, n12637, n12638,
         n12639, n12640, n12641, n12642, n12643, n12644, n12645, n12646,
         n12647, n12648, n12649, n12650, n12651, n12652, n12653, n12654,
         n12655, n12656, n12657, n12658, n12659, n12660, n12661, n12662,
         n12663, n12664, n12665, n12666, n12667, n12668, n12669, n12670,
         n12671, n12672, n12673, n12674, n12675, n12676, n12677, n12678,
         n12679, n12680, n12681, n12682, n12683, n12684, n12685, n12686,
         n12687, n12688, n12689, n12690, n12691, n12692, n12693, n12694,
         n12695, n12696, n12697, n12698, n12699, n12700, n12701, n12702,
         n12703, n12704, n12705, n12706, n12707, n12708, n12709, n12710,
         n12711, n12712, n12713, n12714, n12715, n12716, n12717, n12718,
         n12719, n12720, n12721, n12722, n12723, n12724, n12725, n12726,
         n12727, n12728, n12729, n12730, n12731, n12732, n12733, n12734,
         n12735, n12736, n12737, n12738, n12739, n12740, n12741, n12742,
         n12743, n12744, n12745, n12746, n12747, n12748, n12749, n12750,
         n12751, n12752, n12753, n12754, n12755, n12756, n12757, n12758,
         n12759, n12760, n12761, n12762, n12763, n12764, n12765, n12766,
         n12767, n12768, n12769, n12770, n12771, n12772, n12773, n12774,
         n12775, n12776, n12777, n12778, n12779, n12780, n12781, n12782,
         n12783, n12784, n12785, n12786, n12787, n12788, n12789, n12790,
         n12791, n12792, n12793, n12794, n12795, n12796, n12797, n12798,
         n12799, n12800, n12801, n12802, n12803, n12804, n12805, n12806,
         n12807, n12808, n12809, n12810, n12811, n12812, n12813, n12814,
         n12815, n12816, n12817, n12818, n12819, n12820, n12821, n12822,
         n12823, n12824, n12825, n12826, n12827, n12828, n12829, n12830,
         n12831, n12832, n12833, n12834, n12835, n12836, n12837, n12838,
         n12839, n12840, n12841, n12842, n12843, n12844, n12845, n12846,
         n12847, n12848, n12849, n12850, n12851, n12852, n12853, n12854,
         n12855, n12856, n12857, n12858, n12859, n12860, n12861, n12862,
         n12863, n12864, n12865, n12866, n12867, n12868, n12869, n12870,
         n12871, n12872, n12873, n12874, n12875, n12876, n12877, n12878,
         n12879, n12880, n12881, n12882, n12883, n12884, n12885, n12886,
         n12887, n12888, n12889, n12890, n12891, n12892, n12893, n12894,
         n12895, n12896, n12897, n12898, n12899, n12900, n12901, n12902,
         n12903, n12904, n12905, n12906, n12907, n12908, n12909, n12910,
         n12911, n12912, n12913, n12914, n12915, n12916, n12917, n12918,
         n12919, n12920, n12921, n12922, n12923, n12924, n12925, n12926,
         n12927, n12928, n12929, n12930, n12931, n12932, n12933, n12934,
         n12935, n12936, n12937, n12938, n12939, n12940, n12941, n12942,
         n12943, n12944, n12945, n12946, n12947, n12948, n12949, n12950,
         n12951, n12952, n12953, n12954, n12955, n12956, n12957, n12958,
         n12959, n12960, n12961, n12962, n12963, n12964, n12965, n12966,
         n12967, n12968, n12969, n12970, n12971, n12972, n12973, n12974,
         n12975, n12976, n12977, n12978, n12979, n12980, n12981, n12982,
         n12983, n12984, n12985, n12986, n12987, n12988, n12989, n12990,
         n12991, n12992, n12993, n12994, n12995, n12996, n12997, n12998,
         n12999, n13000, n13001, n13002, n13003, n13004, n13005, n13006,
         n13007, n13008, n13009, n13010, n13011, n13012, n13013, n13014,
         n13015, n13016, n13017, n13018, n13019, n13020, n13021, n13022,
         n13023, n13024, n13025, n13026, n13027, n13028, n13029, n13030,
         n13031, n13032, n13033, n13034, n13035, n13036, n13037, n13038,
         n13039, n13040, n13041, n13042, n13043, n13044, n13045, n13046,
         n13047, n13048, n13049, n13050, n13051, n13052, n13053, n13054,
         n13055, n13056, n13057, n13058, n13059, n13060, n13061, n13062,
         n13063, n13064, n13065, n13066, n13067, n13068, n13069, n13070,
         n13071, n13072, n13073, n13074, n13075, n13076, n13077, n13078,
         n13079, n13080, n13081, n13082, n13083, n13084, n13085, n13086,
         n13087, n13088, n13089, n13090, n13091, n13092, n13093, n13094,
         n13095, n13096, n13097, n13098, n13099, n13100, n13101, n13102,
         n13103, n13104, n13105, n13106, n13107, n13108, n13109, n13110,
         n13111, n13112, n13113, n13114, n13115, n13116, n13117, n13118,
         n13119, n13120, n13121, n13122, n13123, n13124, n13125, n13126,
         n13127, n13128, n13129, n13130, n13131, n13132, n13133, n13134,
         n13135, n13136, n13137, n13138, n13139, n13140, n13141, n13142,
         n13143, n13144, n13145, n13146, n13147, n13148, n13149, n13150,
         n13151, n13152, n13153, n13154, n13155, n13156, n13157, n13158,
         n13159, n13160, n13161, n13162, n13163, n13164, n13165, n13166,
         n13167, n13168, n13169, n13170, n13171, n13172, n13173, n13174,
         n13175, n13176, n13177, n13178, n13179, n13180, n13181, n13182,
         n13183, n13184, n13185, n13186, n13187, n13188, n13189, n13190,
         n13191, n13192, n13193, n13194, n13195, n13196, n13197, n13198,
         n13199, n13200, n13201, n13202, n13203, n13204, n13205, n13206,
         n13207, n13208, n13209, n13210, n13211, n13212, n13213, n13214,
         n13215, n13216, n13217, n13218, n13219, n13220, n13221, n13222,
         n13223, n13224, n13225, n13226, n13227, n13228, n13229, n13230,
         n13231, n13232, n13233, n13234, n13235, n13236, n13237, n13238,
         n13239, n13240, n13241, n13242, n13243, n13244, n13245, n13246,
         n13247, n13248, n13249, n13250, n13251, n13252, n13253, n13254,
         n13255, n13256, n13257, n13258, n13259, n13260, n13261, n13262,
         n13263, n13264, n13265, n13266, n13267, n13268, n13269, n13270,
         n13271, n13272, n13273, n13274, n13275, n13276, n13277, n13278,
         n13279, n13280, n13281, n13282, n13283, n13284, n13285, n13286,
         n13287, n13288, n13289, n13290, n13291, n13292, n13293, n13294,
         n13295, n13296, n13297, n13298, n13299, n13300, n13301, n13302,
         n13303, n13304, n13305, n13306, n13307, n13308, n13309, n13310,
         n13311, n13312, n13313, n13314, n13315, n13316, n13317, n13318,
         n13319, n13320, n13321, n13322, n13323, n13324, n13325, n13326,
         n13327, n13328, n13329, n13330, n13331, n13332, n13333, n13334,
         n13335, n13336, n13337, n13338, n13339, n13340, n13341, n13342,
         n13343, n13344, n13345, n13346, n13347, n13348, n13349, n13350,
         n13351, n13352, n13353, n13354, n13355, n13356, n13357, n13358,
         n13359, n13360, n13361, n13362, n13363, n13364, n13365, n13366,
         n13367, n13368, n13369, n13370, n13371, n13372, n13373, n13374,
         n13375, n13376, n13377, n13378, n13379, n13380, n13381, n13382,
         n13383, n13384, n13385, n13386, n13387, n13388, n13389, n13390,
         n13391, n13392, n13393, n13394, n13395, n13396, n13397, n13398,
         n13399, n13400, n13401, n13402, n13403, n13404, n13405, n13406,
         n13407, n13408, n13409, n13410, n13411, n13412, n13413, n13414,
         n13415, n13416, n13417, n13418, n13419, n13420, n13421, n13422,
         n13423, n13424, n13425, n13426, n13427, n13428, n13429, n13430,
         n13431, n13432, n13433, n13434, n13435, n13436, n13437, n13438,
         n13439, n13440, n13441, n13442, n13443, n13444, n13445, n13446,
         n13447, n13448, n13449, n13450, n13451, n13452, n13453, n13454,
         n13455, n13456, n13457, n13458, n13459, n13460, n13461, n13462,
         n13463, n13464, n13465, n13466, n13467, n13468, n13469, n13470,
         n13471, n13472, n13473, n13474, n13475, n13476, n13477, n13478,
         n13479, n13480, n13481, n13482, n13483, n13484, n13485, n13486,
         n13487, n13488, n13489, n13490, n13491, n13492, n13493, n13494,
         n13495, n13496, n13497, n13498, n13499, n13500, n13501, n13502,
         n13503, n13504, n13505, n13506, n13507, n13508, n13509, n13510,
         n13511, n13512, n13513, n13514, n13515, n13516, n13517, n13518,
         n13519, n13520, n13521, n13522, n13523, n13524, n13525, n13526,
         n13527, n13528, n13529, n13530, n13531, n13532, n13533, n13534,
         n13535, n13536, n13537, n13538, n13539, n13540, n13541, n13542,
         n13543, n13544, n13545, n13546, n13547, n13548, n13549, n13550,
         n13551, n13552, n13553, n13554, n13555, n13556, n13557, n13558,
         n13559, n13560, n13561, n13562, n13563, n13564, n13565, n13566,
         n13567, n13568, n13569, n13570, n13571, n13572, n13573, n13574,
         n13575, n13576, n13577, n13578, n13579, n13580, n13581, n13582,
         n13583, n13584, n13585, n13586, n13587, n13588, n13589, n13590,
         n13591, n13592;
  wire   [4095:0] ram;

  DFF_X1 ram_reg_255__15_ ( .D(n9256), .CK(clk), .Q(ram[4095]) );
  DFF_X1 ram_reg_255__14_ ( .D(n9255), .CK(clk), .Q(ram[4094]) );
  DFF_X1 ram_reg_255__13_ ( .D(n9254), .CK(clk), .Q(ram[4093]) );
  DFF_X1 ram_reg_255__12_ ( .D(n9253), .CK(clk), .Q(ram[4092]) );
  DFF_X1 ram_reg_255__11_ ( .D(n9252), .CK(clk), .Q(ram[4091]) );
  DFF_X1 ram_reg_255__10_ ( .D(n9251), .CK(clk), .Q(ram[4090]) );
  DFF_X1 ram_reg_255__9_ ( .D(n9250), .CK(clk), .Q(ram[4089]) );
  DFF_X1 ram_reg_255__8_ ( .D(n9249), .CK(clk), .Q(ram[4088]) );
  DFF_X1 ram_reg_255__7_ ( .D(n9248), .CK(clk), .Q(ram[4087]) );
  DFF_X1 ram_reg_255__6_ ( .D(n9247), .CK(clk), .Q(ram[4086]) );
  DFF_X1 ram_reg_255__5_ ( .D(n9246), .CK(clk), .Q(ram[4085]) );
  DFF_X1 ram_reg_255__4_ ( .D(n9245), .CK(clk), .Q(ram[4084]) );
  DFF_X1 ram_reg_255__3_ ( .D(n9244), .CK(clk), .Q(ram[4083]) );
  DFF_X1 ram_reg_255__2_ ( .D(n9243), .CK(clk), .Q(ram[4082]) );
  DFF_X1 ram_reg_255__1_ ( .D(n9242), .CK(clk), .Q(ram[4081]) );
  DFF_X1 ram_reg_255__0_ ( .D(n9241), .CK(clk), .Q(ram[4080]) );
  DFF_X1 ram_reg_254__15_ ( .D(n9273), .CK(clk), .Q(ram[4079]) );
  DFF_X1 ram_reg_254__14_ ( .D(n9272), .CK(clk), .Q(ram[4078]) );
  DFF_X1 ram_reg_254__13_ ( .D(n9271), .CK(clk), .Q(ram[4077]) );
  DFF_X1 ram_reg_254__12_ ( .D(n9270), .CK(clk), .Q(ram[4076]) );
  DFF_X1 ram_reg_254__11_ ( .D(n9269), .CK(clk), .Q(ram[4075]) );
  DFF_X1 ram_reg_254__10_ ( .D(n9268), .CK(clk), .Q(ram[4074]) );
  DFF_X1 ram_reg_254__9_ ( .D(n9267), .CK(clk), .Q(ram[4073]) );
  DFF_X1 ram_reg_254__8_ ( .D(n9266), .CK(clk), .Q(ram[4072]) );
  DFF_X1 ram_reg_254__7_ ( .D(n9265), .CK(clk), .Q(ram[4071]) );
  DFF_X1 ram_reg_254__6_ ( .D(n9264), .CK(clk), .Q(ram[4070]) );
  DFF_X1 ram_reg_254__5_ ( .D(n9263), .CK(clk), .Q(ram[4069]) );
  DFF_X1 ram_reg_254__4_ ( .D(n9262), .CK(clk), .Q(ram[4068]) );
  DFF_X1 ram_reg_254__3_ ( .D(n9261), .CK(clk), .Q(ram[4067]) );
  DFF_X1 ram_reg_254__2_ ( .D(n9260), .CK(clk), .Q(ram[4066]) );
  DFF_X1 ram_reg_254__1_ ( .D(n9259), .CK(clk), .Q(ram[4065]) );
  DFF_X1 ram_reg_254__0_ ( .D(n9258), .CK(clk), .Q(ram[4064]) );
  DFF_X1 ram_reg_253__15_ ( .D(n9290), .CK(clk), .Q(ram[4063]) );
  DFF_X1 ram_reg_253__14_ ( .D(n9289), .CK(clk), .Q(ram[4062]) );
  DFF_X1 ram_reg_253__13_ ( .D(n9288), .CK(clk), .Q(ram[4061]) );
  DFF_X1 ram_reg_253__12_ ( .D(n9287), .CK(clk), .Q(ram[4060]) );
  DFF_X1 ram_reg_253__11_ ( .D(n9286), .CK(clk), .Q(ram[4059]) );
  DFF_X1 ram_reg_253__10_ ( .D(n9285), .CK(clk), .Q(ram[4058]) );
  DFF_X1 ram_reg_253__9_ ( .D(n9284), .CK(clk), .Q(ram[4057]) );
  DFF_X1 ram_reg_253__8_ ( .D(n9283), .CK(clk), .Q(ram[4056]) );
  DFF_X1 ram_reg_253__7_ ( .D(n9282), .CK(clk), .Q(ram[4055]) );
  DFF_X1 ram_reg_253__6_ ( .D(n9281), .CK(clk), .Q(ram[4054]) );
  DFF_X1 ram_reg_253__5_ ( .D(n9280), .CK(clk), .Q(ram[4053]) );
  DFF_X1 ram_reg_253__4_ ( .D(n9279), .CK(clk), .Q(ram[4052]) );
  DFF_X1 ram_reg_253__3_ ( .D(n9278), .CK(clk), .Q(ram[4051]) );
  DFF_X1 ram_reg_253__2_ ( .D(n9277), .CK(clk), .Q(ram[4050]) );
  DFF_X1 ram_reg_253__1_ ( .D(n9276), .CK(clk), .Q(ram[4049]) );
  DFF_X1 ram_reg_253__0_ ( .D(n9275), .CK(clk), .Q(ram[4048]) );
  DFF_X1 ram_reg_252__15_ ( .D(n9307), .CK(clk), .Q(ram[4047]) );
  DFF_X1 ram_reg_252__14_ ( .D(n9306), .CK(clk), .Q(ram[4046]) );
  DFF_X1 ram_reg_252__13_ ( .D(n9305), .CK(clk), .Q(ram[4045]) );
  DFF_X1 ram_reg_252__12_ ( .D(n9304), .CK(clk), .Q(ram[4044]) );
  DFF_X1 ram_reg_252__11_ ( .D(n9303), .CK(clk), .Q(ram[4043]) );
  DFF_X1 ram_reg_252__10_ ( .D(n9302), .CK(clk), .Q(ram[4042]) );
  DFF_X1 ram_reg_252__9_ ( .D(n9301), .CK(clk), .Q(ram[4041]) );
  DFF_X1 ram_reg_252__8_ ( .D(n9300), .CK(clk), .Q(ram[4040]) );
  DFF_X1 ram_reg_252__7_ ( .D(n9299), .CK(clk), .Q(ram[4039]) );
  DFF_X1 ram_reg_252__6_ ( .D(n9298), .CK(clk), .Q(ram[4038]) );
  DFF_X1 ram_reg_252__5_ ( .D(n9297), .CK(clk), .Q(ram[4037]) );
  DFF_X1 ram_reg_252__4_ ( .D(n9296), .CK(clk), .Q(ram[4036]) );
  DFF_X1 ram_reg_252__3_ ( .D(n9295), .CK(clk), .Q(ram[4035]) );
  DFF_X1 ram_reg_252__2_ ( .D(n9294), .CK(clk), .Q(ram[4034]) );
  DFF_X1 ram_reg_252__1_ ( .D(n9293), .CK(clk), .Q(ram[4033]) );
  DFF_X1 ram_reg_252__0_ ( .D(n9292), .CK(clk), .Q(ram[4032]) );
  DFF_X1 ram_reg_251__15_ ( .D(n9324), .CK(clk), .Q(ram[4031]) );
  DFF_X1 ram_reg_251__14_ ( .D(n9323), .CK(clk), .Q(ram[4030]) );
  DFF_X1 ram_reg_251__13_ ( .D(n9322), .CK(clk), .Q(ram[4029]) );
  DFF_X1 ram_reg_251__12_ ( .D(n9321), .CK(clk), .Q(ram[4028]) );
  DFF_X1 ram_reg_251__11_ ( .D(n9320), .CK(clk), .Q(ram[4027]) );
  DFF_X1 ram_reg_251__10_ ( .D(n9319), .CK(clk), .Q(ram[4026]) );
  DFF_X1 ram_reg_251__9_ ( .D(n9318), .CK(clk), .Q(ram[4025]) );
  DFF_X1 ram_reg_251__8_ ( .D(n9317), .CK(clk), .Q(ram[4024]) );
  DFF_X1 ram_reg_251__7_ ( .D(n9316), .CK(clk), .Q(ram[4023]) );
  DFF_X1 ram_reg_251__6_ ( .D(n9315), .CK(clk), .Q(ram[4022]) );
  DFF_X1 ram_reg_251__5_ ( .D(n9314), .CK(clk), .Q(ram[4021]) );
  DFF_X1 ram_reg_251__4_ ( .D(n9313), .CK(clk), .Q(ram[4020]) );
  DFF_X1 ram_reg_251__3_ ( .D(n9312), .CK(clk), .Q(ram[4019]) );
  DFF_X1 ram_reg_251__2_ ( .D(n9311), .CK(clk), .Q(ram[4018]) );
  DFF_X1 ram_reg_251__1_ ( .D(n9310), .CK(clk), .Q(ram[4017]) );
  DFF_X1 ram_reg_251__0_ ( .D(n9309), .CK(clk), .Q(ram[4016]) );
  DFF_X1 ram_reg_250__15_ ( .D(n9341), .CK(clk), .Q(ram[4015]) );
  DFF_X1 ram_reg_250__14_ ( .D(n9340), .CK(clk), .Q(ram[4014]) );
  DFF_X1 ram_reg_250__13_ ( .D(n9339), .CK(clk), .Q(ram[4013]) );
  DFF_X1 ram_reg_250__12_ ( .D(n9338), .CK(clk), .Q(ram[4012]) );
  DFF_X1 ram_reg_250__11_ ( .D(n9337), .CK(clk), .Q(ram[4011]) );
  DFF_X1 ram_reg_250__10_ ( .D(n9336), .CK(clk), .Q(ram[4010]) );
  DFF_X1 ram_reg_250__9_ ( .D(n9335), .CK(clk), .Q(ram[4009]) );
  DFF_X1 ram_reg_250__8_ ( .D(n9334), .CK(clk), .Q(ram[4008]) );
  DFF_X1 ram_reg_250__7_ ( .D(n9333), .CK(clk), .Q(ram[4007]) );
  DFF_X1 ram_reg_250__6_ ( .D(n9332), .CK(clk), .Q(ram[4006]) );
  DFF_X1 ram_reg_250__5_ ( .D(n9331), .CK(clk), .Q(ram[4005]) );
  DFF_X1 ram_reg_250__4_ ( .D(n9330), .CK(clk), .Q(ram[4004]) );
  DFF_X1 ram_reg_250__3_ ( .D(n9329), .CK(clk), .Q(ram[4003]) );
  DFF_X1 ram_reg_250__2_ ( .D(n9328), .CK(clk), .Q(ram[4002]) );
  DFF_X1 ram_reg_250__1_ ( .D(n9327), .CK(clk), .Q(ram[4001]) );
  DFF_X1 ram_reg_250__0_ ( .D(n9326), .CK(clk), .Q(ram[4000]) );
  DFF_X1 ram_reg_249__15_ ( .D(n9358), .CK(clk), .Q(ram[3999]) );
  DFF_X1 ram_reg_249__14_ ( .D(n9357), .CK(clk), .Q(ram[3998]) );
  DFF_X1 ram_reg_249__13_ ( .D(n9356), .CK(clk), .Q(ram[3997]) );
  DFF_X1 ram_reg_249__12_ ( .D(n9355), .CK(clk), .Q(ram[3996]) );
  DFF_X1 ram_reg_249__11_ ( .D(n9354), .CK(clk), .Q(ram[3995]) );
  DFF_X1 ram_reg_249__10_ ( .D(n9353), .CK(clk), .Q(ram[3994]) );
  DFF_X1 ram_reg_249__9_ ( .D(n9352), .CK(clk), .Q(ram[3993]) );
  DFF_X1 ram_reg_249__8_ ( .D(n9351), .CK(clk), .Q(ram[3992]) );
  DFF_X1 ram_reg_249__7_ ( .D(n9350), .CK(clk), .Q(ram[3991]) );
  DFF_X1 ram_reg_249__6_ ( .D(n9349), .CK(clk), .Q(ram[3990]) );
  DFF_X1 ram_reg_249__5_ ( .D(n9348), .CK(clk), .Q(ram[3989]) );
  DFF_X1 ram_reg_249__4_ ( .D(n9347), .CK(clk), .Q(ram[3988]) );
  DFF_X1 ram_reg_249__3_ ( .D(n9346), .CK(clk), .Q(ram[3987]) );
  DFF_X1 ram_reg_249__2_ ( .D(n9345), .CK(clk), .Q(ram[3986]) );
  DFF_X1 ram_reg_249__1_ ( .D(n9344), .CK(clk), .Q(ram[3985]) );
  DFF_X1 ram_reg_249__0_ ( .D(n9343), .CK(clk), .Q(ram[3984]) );
  DFF_X1 ram_reg_248__15_ ( .D(n9375), .CK(clk), .Q(ram[3983]) );
  DFF_X1 ram_reg_248__14_ ( .D(n9374), .CK(clk), .Q(ram[3982]) );
  DFF_X1 ram_reg_248__13_ ( .D(n9373), .CK(clk), .Q(ram[3981]) );
  DFF_X1 ram_reg_248__12_ ( .D(n9372), .CK(clk), .Q(ram[3980]) );
  DFF_X1 ram_reg_248__11_ ( .D(n9371), .CK(clk), .Q(ram[3979]) );
  DFF_X1 ram_reg_248__10_ ( .D(n9370), .CK(clk), .Q(ram[3978]) );
  DFF_X1 ram_reg_248__9_ ( .D(n9369), .CK(clk), .Q(ram[3977]) );
  DFF_X1 ram_reg_248__8_ ( .D(n9368), .CK(clk), .Q(ram[3976]) );
  DFF_X1 ram_reg_248__7_ ( .D(n9367), .CK(clk), .Q(ram[3975]) );
  DFF_X1 ram_reg_248__6_ ( .D(n9366), .CK(clk), .Q(ram[3974]) );
  DFF_X1 ram_reg_248__5_ ( .D(n9365), .CK(clk), .Q(ram[3973]) );
  DFF_X1 ram_reg_248__4_ ( .D(n9364), .CK(clk), .Q(ram[3972]) );
  DFF_X1 ram_reg_248__3_ ( .D(n9363), .CK(clk), .Q(ram[3971]) );
  DFF_X1 ram_reg_248__2_ ( .D(n9362), .CK(clk), .Q(ram[3970]) );
  DFF_X1 ram_reg_248__1_ ( .D(n9361), .CK(clk), .Q(ram[3969]) );
  DFF_X1 ram_reg_248__0_ ( .D(n9360), .CK(clk), .Q(ram[3968]) );
  DFF_X1 ram_reg_247__15_ ( .D(n9392), .CK(clk), .Q(ram[3967]) );
  DFF_X1 ram_reg_247__14_ ( .D(n9391), .CK(clk), .Q(ram[3966]) );
  DFF_X1 ram_reg_247__13_ ( .D(n9390), .CK(clk), .Q(ram[3965]) );
  DFF_X1 ram_reg_247__12_ ( .D(n9389), .CK(clk), .Q(ram[3964]) );
  DFF_X1 ram_reg_247__11_ ( .D(n9388), .CK(clk), .Q(ram[3963]) );
  DFF_X1 ram_reg_247__10_ ( .D(n9387), .CK(clk), .Q(ram[3962]) );
  DFF_X1 ram_reg_247__9_ ( .D(n9386), .CK(clk), .Q(ram[3961]) );
  DFF_X1 ram_reg_247__8_ ( .D(n9385), .CK(clk), .Q(ram[3960]) );
  DFF_X1 ram_reg_247__7_ ( .D(n9384), .CK(clk), .Q(ram[3959]) );
  DFF_X1 ram_reg_247__6_ ( .D(n9383), .CK(clk), .Q(ram[3958]) );
  DFF_X1 ram_reg_247__5_ ( .D(n9382), .CK(clk), .Q(ram[3957]) );
  DFF_X1 ram_reg_247__4_ ( .D(n9381), .CK(clk), .Q(ram[3956]) );
  DFF_X1 ram_reg_247__3_ ( .D(n9380), .CK(clk), .Q(ram[3955]) );
  DFF_X1 ram_reg_247__2_ ( .D(n9379), .CK(clk), .Q(ram[3954]) );
  DFF_X1 ram_reg_247__1_ ( .D(n9378), .CK(clk), .Q(ram[3953]) );
  DFF_X1 ram_reg_247__0_ ( .D(n9377), .CK(clk), .Q(ram[3952]) );
  DFF_X1 ram_reg_246__15_ ( .D(n9409), .CK(clk), .Q(ram[3951]) );
  DFF_X1 ram_reg_246__14_ ( .D(n9408), .CK(clk), .Q(ram[3950]) );
  DFF_X1 ram_reg_246__13_ ( .D(n9407), .CK(clk), .Q(ram[3949]) );
  DFF_X1 ram_reg_246__12_ ( .D(n9406), .CK(clk), .Q(ram[3948]) );
  DFF_X1 ram_reg_246__11_ ( .D(n9405), .CK(clk), .Q(ram[3947]) );
  DFF_X1 ram_reg_246__10_ ( .D(n9404), .CK(clk), .Q(ram[3946]) );
  DFF_X1 ram_reg_246__9_ ( .D(n9403), .CK(clk), .Q(ram[3945]) );
  DFF_X1 ram_reg_246__8_ ( .D(n9402), .CK(clk), .Q(ram[3944]) );
  DFF_X1 ram_reg_246__7_ ( .D(n9401), .CK(clk), .Q(ram[3943]) );
  DFF_X1 ram_reg_246__6_ ( .D(n9400), .CK(clk), .Q(ram[3942]) );
  DFF_X1 ram_reg_246__5_ ( .D(n9399), .CK(clk), .Q(ram[3941]) );
  DFF_X1 ram_reg_246__4_ ( .D(n9398), .CK(clk), .Q(ram[3940]) );
  DFF_X1 ram_reg_246__3_ ( .D(n9397), .CK(clk), .Q(ram[3939]) );
  DFF_X1 ram_reg_246__2_ ( .D(n9396), .CK(clk), .Q(ram[3938]) );
  DFF_X1 ram_reg_246__1_ ( .D(n9395), .CK(clk), .Q(ram[3937]) );
  DFF_X1 ram_reg_246__0_ ( .D(n9394), .CK(clk), .Q(ram[3936]) );
  DFF_X1 ram_reg_245__15_ ( .D(n9426), .CK(clk), .Q(ram[3935]) );
  DFF_X1 ram_reg_245__14_ ( .D(n9425), .CK(clk), .Q(ram[3934]) );
  DFF_X1 ram_reg_245__13_ ( .D(n9424), .CK(clk), .Q(ram[3933]) );
  DFF_X1 ram_reg_245__12_ ( .D(n9423), .CK(clk), .Q(ram[3932]) );
  DFF_X1 ram_reg_245__11_ ( .D(n9422), .CK(clk), .Q(ram[3931]) );
  DFF_X1 ram_reg_245__10_ ( .D(n9421), .CK(clk), .Q(ram[3930]) );
  DFF_X1 ram_reg_245__9_ ( .D(n9420), .CK(clk), .Q(ram[3929]) );
  DFF_X1 ram_reg_245__8_ ( .D(n9419), .CK(clk), .Q(ram[3928]) );
  DFF_X1 ram_reg_245__7_ ( .D(n9418), .CK(clk), .Q(ram[3927]) );
  DFF_X1 ram_reg_245__6_ ( .D(n9417), .CK(clk), .Q(ram[3926]) );
  DFF_X1 ram_reg_245__5_ ( .D(n9416), .CK(clk), .Q(ram[3925]) );
  DFF_X1 ram_reg_245__4_ ( .D(n9415), .CK(clk), .Q(ram[3924]) );
  DFF_X1 ram_reg_245__3_ ( .D(n9414), .CK(clk), .Q(ram[3923]) );
  DFF_X1 ram_reg_245__2_ ( .D(n9413), .CK(clk), .Q(ram[3922]) );
  DFF_X1 ram_reg_245__1_ ( .D(n9412), .CK(clk), .Q(ram[3921]) );
  DFF_X1 ram_reg_245__0_ ( .D(n9411), .CK(clk), .Q(ram[3920]) );
  DFF_X1 ram_reg_244__15_ ( .D(n9443), .CK(clk), .Q(ram[3919]) );
  DFF_X1 ram_reg_244__14_ ( .D(n9442), .CK(clk), .Q(ram[3918]) );
  DFF_X1 ram_reg_244__13_ ( .D(n9441), .CK(clk), .Q(ram[3917]) );
  DFF_X1 ram_reg_244__12_ ( .D(n9440), .CK(clk), .Q(ram[3916]) );
  DFF_X1 ram_reg_244__11_ ( .D(n9439), .CK(clk), .Q(ram[3915]) );
  DFF_X1 ram_reg_244__10_ ( .D(n9438), .CK(clk), .Q(ram[3914]) );
  DFF_X1 ram_reg_244__9_ ( .D(n9437), .CK(clk), .Q(ram[3913]) );
  DFF_X1 ram_reg_244__8_ ( .D(n9436), .CK(clk), .Q(ram[3912]) );
  DFF_X1 ram_reg_244__7_ ( .D(n9435), .CK(clk), .Q(ram[3911]) );
  DFF_X1 ram_reg_244__6_ ( .D(n9434), .CK(clk), .Q(ram[3910]) );
  DFF_X1 ram_reg_244__5_ ( .D(n9433), .CK(clk), .Q(ram[3909]) );
  DFF_X1 ram_reg_244__4_ ( .D(n9432), .CK(clk), .Q(ram[3908]) );
  DFF_X1 ram_reg_244__3_ ( .D(n9431), .CK(clk), .Q(ram[3907]) );
  DFF_X1 ram_reg_244__2_ ( .D(n9430), .CK(clk), .Q(ram[3906]) );
  DFF_X1 ram_reg_244__1_ ( .D(n9429), .CK(clk), .Q(ram[3905]) );
  DFF_X1 ram_reg_244__0_ ( .D(n9428), .CK(clk), .Q(ram[3904]) );
  DFF_X1 ram_reg_243__15_ ( .D(n9460), .CK(clk), .Q(ram[3903]) );
  DFF_X1 ram_reg_243__14_ ( .D(n9459), .CK(clk), .Q(ram[3902]) );
  DFF_X1 ram_reg_243__13_ ( .D(n9458), .CK(clk), .Q(ram[3901]) );
  DFF_X1 ram_reg_243__12_ ( .D(n9457), .CK(clk), .Q(ram[3900]) );
  DFF_X1 ram_reg_243__11_ ( .D(n9456), .CK(clk), .Q(ram[3899]) );
  DFF_X1 ram_reg_243__10_ ( .D(n9455), .CK(clk), .Q(ram[3898]) );
  DFF_X1 ram_reg_243__9_ ( .D(n9454), .CK(clk), .Q(ram[3897]) );
  DFF_X1 ram_reg_243__8_ ( .D(n9453), .CK(clk), .Q(ram[3896]) );
  DFF_X1 ram_reg_243__7_ ( .D(n9452), .CK(clk), .Q(ram[3895]) );
  DFF_X1 ram_reg_243__6_ ( .D(n9451), .CK(clk), .Q(ram[3894]) );
  DFF_X1 ram_reg_243__5_ ( .D(n9450), .CK(clk), .Q(ram[3893]) );
  DFF_X1 ram_reg_243__4_ ( .D(n9449), .CK(clk), .Q(ram[3892]) );
  DFF_X1 ram_reg_243__3_ ( .D(n9448), .CK(clk), .Q(ram[3891]) );
  DFF_X1 ram_reg_243__2_ ( .D(n9447), .CK(clk), .Q(ram[3890]) );
  DFF_X1 ram_reg_243__1_ ( .D(n9446), .CK(clk), .Q(ram[3889]) );
  DFF_X1 ram_reg_243__0_ ( .D(n9445), .CK(clk), .Q(ram[3888]) );
  DFF_X1 ram_reg_242__15_ ( .D(n9477), .CK(clk), .Q(ram[3887]) );
  DFF_X1 ram_reg_242__14_ ( .D(n9476), .CK(clk), .Q(ram[3886]) );
  DFF_X1 ram_reg_242__13_ ( .D(n9475), .CK(clk), .Q(ram[3885]) );
  DFF_X1 ram_reg_242__12_ ( .D(n9474), .CK(clk), .Q(ram[3884]) );
  DFF_X1 ram_reg_242__11_ ( .D(n9473), .CK(clk), .Q(ram[3883]) );
  DFF_X1 ram_reg_242__10_ ( .D(n9472), .CK(clk), .Q(ram[3882]) );
  DFF_X1 ram_reg_242__9_ ( .D(n9471), .CK(clk), .Q(ram[3881]) );
  DFF_X1 ram_reg_242__8_ ( .D(n9470), .CK(clk), .Q(ram[3880]) );
  DFF_X1 ram_reg_242__7_ ( .D(n9469), .CK(clk), .Q(ram[3879]) );
  DFF_X1 ram_reg_242__6_ ( .D(n9468), .CK(clk), .Q(ram[3878]) );
  DFF_X1 ram_reg_242__5_ ( .D(n9467), .CK(clk), .Q(ram[3877]) );
  DFF_X1 ram_reg_242__4_ ( .D(n9466), .CK(clk), .Q(ram[3876]) );
  DFF_X1 ram_reg_242__3_ ( .D(n9465), .CK(clk), .Q(ram[3875]) );
  DFF_X1 ram_reg_242__2_ ( .D(n9464), .CK(clk), .Q(ram[3874]) );
  DFF_X1 ram_reg_242__1_ ( .D(n9463), .CK(clk), .Q(ram[3873]) );
  DFF_X1 ram_reg_242__0_ ( .D(n9462), .CK(clk), .Q(ram[3872]) );
  DFF_X1 ram_reg_241__15_ ( .D(n9494), .CK(clk), .Q(ram[3871]) );
  DFF_X1 ram_reg_241__14_ ( .D(n9493), .CK(clk), .Q(ram[3870]) );
  DFF_X1 ram_reg_241__13_ ( .D(n9492), .CK(clk), .Q(ram[3869]) );
  DFF_X1 ram_reg_241__12_ ( .D(n9491), .CK(clk), .Q(ram[3868]) );
  DFF_X1 ram_reg_241__11_ ( .D(n9490), .CK(clk), .Q(ram[3867]) );
  DFF_X1 ram_reg_241__10_ ( .D(n9489), .CK(clk), .Q(ram[3866]) );
  DFF_X1 ram_reg_241__9_ ( .D(n9488), .CK(clk), .Q(ram[3865]) );
  DFF_X1 ram_reg_241__8_ ( .D(n9487), .CK(clk), .Q(ram[3864]) );
  DFF_X1 ram_reg_241__7_ ( .D(n9486), .CK(clk), .Q(ram[3863]) );
  DFF_X1 ram_reg_241__6_ ( .D(n9485), .CK(clk), .Q(ram[3862]) );
  DFF_X1 ram_reg_241__5_ ( .D(n9484), .CK(clk), .Q(ram[3861]) );
  DFF_X1 ram_reg_241__4_ ( .D(n9483), .CK(clk), .Q(ram[3860]) );
  DFF_X1 ram_reg_241__3_ ( .D(n9482), .CK(clk), .Q(ram[3859]) );
  DFF_X1 ram_reg_241__2_ ( .D(n9481), .CK(clk), .Q(ram[3858]) );
  DFF_X1 ram_reg_241__1_ ( .D(n9480), .CK(clk), .Q(ram[3857]) );
  DFF_X1 ram_reg_241__0_ ( .D(n9479), .CK(clk), .Q(ram[3856]) );
  DFF_X1 ram_reg_240__15_ ( .D(n9511), .CK(clk), .Q(ram[3855]) );
  DFF_X1 ram_reg_240__14_ ( .D(n9510), .CK(clk), .Q(ram[3854]) );
  DFF_X1 ram_reg_240__13_ ( .D(n9509), .CK(clk), .Q(ram[3853]) );
  DFF_X1 ram_reg_240__12_ ( .D(n9508), .CK(clk), .Q(ram[3852]) );
  DFF_X1 ram_reg_240__11_ ( .D(n9507), .CK(clk), .Q(ram[3851]) );
  DFF_X1 ram_reg_240__10_ ( .D(n9506), .CK(clk), .Q(ram[3850]) );
  DFF_X1 ram_reg_240__9_ ( .D(n9505), .CK(clk), .Q(ram[3849]) );
  DFF_X1 ram_reg_240__8_ ( .D(n9504), .CK(clk), .Q(ram[3848]) );
  DFF_X1 ram_reg_240__7_ ( .D(n9503), .CK(clk), .Q(ram[3847]) );
  DFF_X1 ram_reg_240__6_ ( .D(n9502), .CK(clk), .Q(ram[3846]) );
  DFF_X1 ram_reg_240__5_ ( .D(n9501), .CK(clk), .Q(ram[3845]) );
  DFF_X1 ram_reg_240__4_ ( .D(n9500), .CK(clk), .Q(ram[3844]) );
  DFF_X1 ram_reg_240__3_ ( .D(n9499), .CK(clk), .Q(ram[3843]) );
  DFF_X1 ram_reg_240__2_ ( .D(n9498), .CK(clk), .Q(ram[3842]) );
  DFF_X1 ram_reg_240__1_ ( .D(n9497), .CK(clk), .Q(ram[3841]) );
  DFF_X1 ram_reg_240__0_ ( .D(n9496), .CK(clk), .Q(ram[3840]) );
  DFF_X1 ram_reg_239__15_ ( .D(n9528), .CK(clk), .Q(ram[3839]) );
  DFF_X1 ram_reg_239__14_ ( .D(n9527), .CK(clk), .Q(ram[3838]) );
  DFF_X1 ram_reg_239__13_ ( .D(n9526), .CK(clk), .Q(ram[3837]) );
  DFF_X1 ram_reg_239__12_ ( .D(n9525), .CK(clk), .Q(ram[3836]) );
  DFF_X1 ram_reg_239__11_ ( .D(n9524), .CK(clk), .Q(ram[3835]) );
  DFF_X1 ram_reg_239__10_ ( .D(n9523), .CK(clk), .Q(ram[3834]) );
  DFF_X1 ram_reg_239__9_ ( .D(n9522), .CK(clk), .Q(ram[3833]) );
  DFF_X1 ram_reg_239__8_ ( .D(n9521), .CK(clk), .Q(ram[3832]) );
  DFF_X1 ram_reg_239__7_ ( .D(n9520), .CK(clk), .Q(ram[3831]) );
  DFF_X1 ram_reg_239__6_ ( .D(n9519), .CK(clk), .Q(ram[3830]) );
  DFF_X1 ram_reg_239__5_ ( .D(n9518), .CK(clk), .Q(ram[3829]) );
  DFF_X1 ram_reg_239__4_ ( .D(n9517), .CK(clk), .Q(ram[3828]) );
  DFF_X1 ram_reg_239__3_ ( .D(n9516), .CK(clk), .Q(ram[3827]) );
  DFF_X1 ram_reg_239__2_ ( .D(n9515), .CK(clk), .Q(ram[3826]) );
  DFF_X1 ram_reg_239__1_ ( .D(n9514), .CK(clk), .Q(ram[3825]) );
  DFF_X1 ram_reg_239__0_ ( .D(n9513), .CK(clk), .Q(ram[3824]) );
  DFF_X1 ram_reg_238__15_ ( .D(n9545), .CK(clk), .Q(ram[3823]) );
  DFF_X1 ram_reg_238__14_ ( .D(n9544), .CK(clk), .Q(ram[3822]) );
  DFF_X1 ram_reg_238__13_ ( .D(n9543), .CK(clk), .Q(ram[3821]) );
  DFF_X1 ram_reg_238__12_ ( .D(n9542), .CK(clk), .Q(ram[3820]) );
  DFF_X1 ram_reg_238__11_ ( .D(n9541), .CK(clk), .Q(ram[3819]) );
  DFF_X1 ram_reg_238__10_ ( .D(n9540), .CK(clk), .Q(ram[3818]) );
  DFF_X1 ram_reg_238__9_ ( .D(n9539), .CK(clk), .Q(ram[3817]) );
  DFF_X1 ram_reg_238__8_ ( .D(n9538), .CK(clk), .Q(ram[3816]) );
  DFF_X1 ram_reg_238__7_ ( .D(n9537), .CK(clk), .Q(ram[3815]) );
  DFF_X1 ram_reg_238__6_ ( .D(n9536), .CK(clk), .Q(ram[3814]) );
  DFF_X1 ram_reg_238__5_ ( .D(n9535), .CK(clk), .Q(ram[3813]) );
  DFF_X1 ram_reg_238__4_ ( .D(n9534), .CK(clk), .Q(ram[3812]) );
  DFF_X1 ram_reg_238__3_ ( .D(n9533), .CK(clk), .Q(ram[3811]) );
  DFF_X1 ram_reg_238__2_ ( .D(n9532), .CK(clk), .Q(ram[3810]) );
  DFF_X1 ram_reg_238__1_ ( .D(n9531), .CK(clk), .Q(ram[3809]) );
  DFF_X1 ram_reg_238__0_ ( .D(n9530), .CK(clk), .Q(ram[3808]) );
  DFF_X1 ram_reg_237__15_ ( .D(n9562), .CK(clk), .Q(ram[3807]) );
  DFF_X1 ram_reg_237__14_ ( .D(n9561), .CK(clk), .Q(ram[3806]) );
  DFF_X1 ram_reg_237__13_ ( .D(n9560), .CK(clk), .Q(ram[3805]) );
  DFF_X1 ram_reg_237__12_ ( .D(n9559), .CK(clk), .Q(ram[3804]) );
  DFF_X1 ram_reg_237__11_ ( .D(n9558), .CK(clk), .Q(ram[3803]) );
  DFF_X1 ram_reg_237__10_ ( .D(n9557), .CK(clk), .Q(ram[3802]) );
  DFF_X1 ram_reg_237__9_ ( .D(n9556), .CK(clk), .Q(ram[3801]) );
  DFF_X1 ram_reg_237__8_ ( .D(n9555), .CK(clk), .Q(ram[3800]) );
  DFF_X1 ram_reg_237__7_ ( .D(n9554), .CK(clk), .Q(ram[3799]) );
  DFF_X1 ram_reg_237__6_ ( .D(n9553), .CK(clk), .Q(ram[3798]) );
  DFF_X1 ram_reg_237__5_ ( .D(n9552), .CK(clk), .Q(ram[3797]) );
  DFF_X1 ram_reg_237__4_ ( .D(n9551), .CK(clk), .Q(ram[3796]) );
  DFF_X1 ram_reg_237__3_ ( .D(n9550), .CK(clk), .Q(ram[3795]) );
  DFF_X1 ram_reg_237__2_ ( .D(n9549), .CK(clk), .Q(ram[3794]) );
  DFF_X1 ram_reg_237__1_ ( .D(n9548), .CK(clk), .Q(ram[3793]) );
  DFF_X1 ram_reg_237__0_ ( .D(n9547), .CK(clk), .Q(ram[3792]) );
  DFF_X1 ram_reg_236__15_ ( .D(n9579), .CK(clk), .Q(ram[3791]) );
  DFF_X1 ram_reg_236__14_ ( .D(n9578), .CK(clk), .Q(ram[3790]) );
  DFF_X1 ram_reg_236__13_ ( .D(n9577), .CK(clk), .Q(ram[3789]) );
  DFF_X1 ram_reg_236__12_ ( .D(n9576), .CK(clk), .Q(ram[3788]) );
  DFF_X1 ram_reg_236__11_ ( .D(n9575), .CK(clk), .Q(ram[3787]) );
  DFF_X1 ram_reg_236__10_ ( .D(n9574), .CK(clk), .Q(ram[3786]) );
  DFF_X1 ram_reg_236__9_ ( .D(n9573), .CK(clk), .Q(ram[3785]) );
  DFF_X1 ram_reg_236__8_ ( .D(n9572), .CK(clk), .Q(ram[3784]) );
  DFF_X1 ram_reg_236__7_ ( .D(n9571), .CK(clk), .Q(ram[3783]) );
  DFF_X1 ram_reg_236__6_ ( .D(n9570), .CK(clk), .Q(ram[3782]) );
  DFF_X1 ram_reg_236__5_ ( .D(n9569), .CK(clk), .Q(ram[3781]) );
  DFF_X1 ram_reg_236__4_ ( .D(n9568), .CK(clk), .Q(ram[3780]) );
  DFF_X1 ram_reg_236__3_ ( .D(n9567), .CK(clk), .Q(ram[3779]) );
  DFF_X1 ram_reg_236__2_ ( .D(n9566), .CK(clk), .Q(ram[3778]) );
  DFF_X1 ram_reg_236__1_ ( .D(n9565), .CK(clk), .Q(ram[3777]) );
  DFF_X1 ram_reg_236__0_ ( .D(n9564), .CK(clk), .Q(ram[3776]) );
  DFF_X1 ram_reg_235__15_ ( .D(n9596), .CK(clk), .Q(ram[3775]) );
  DFF_X1 ram_reg_235__14_ ( .D(n9595), .CK(clk), .Q(ram[3774]) );
  DFF_X1 ram_reg_235__13_ ( .D(n9594), .CK(clk), .Q(ram[3773]) );
  DFF_X1 ram_reg_235__12_ ( .D(n9593), .CK(clk), .Q(ram[3772]) );
  DFF_X1 ram_reg_235__11_ ( .D(n9592), .CK(clk), .Q(ram[3771]) );
  DFF_X1 ram_reg_235__10_ ( .D(n9591), .CK(clk), .Q(ram[3770]) );
  DFF_X1 ram_reg_235__9_ ( .D(n9590), .CK(clk), .Q(ram[3769]) );
  DFF_X1 ram_reg_235__8_ ( .D(n9589), .CK(clk), .Q(ram[3768]) );
  DFF_X1 ram_reg_235__7_ ( .D(n9588), .CK(clk), .Q(ram[3767]) );
  DFF_X1 ram_reg_235__6_ ( .D(n9587), .CK(clk), .Q(ram[3766]) );
  DFF_X1 ram_reg_235__5_ ( .D(n9586), .CK(clk), .Q(ram[3765]) );
  DFF_X1 ram_reg_235__4_ ( .D(n9585), .CK(clk), .Q(ram[3764]) );
  DFF_X1 ram_reg_235__3_ ( .D(n9584), .CK(clk), .Q(ram[3763]) );
  DFF_X1 ram_reg_235__2_ ( .D(n9583), .CK(clk), .Q(ram[3762]) );
  DFF_X1 ram_reg_235__1_ ( .D(n9582), .CK(clk), .Q(ram[3761]) );
  DFF_X1 ram_reg_235__0_ ( .D(n9581), .CK(clk), .Q(ram[3760]) );
  DFF_X1 ram_reg_234__15_ ( .D(n9613), .CK(clk), .Q(ram[3759]) );
  DFF_X1 ram_reg_234__14_ ( .D(n9612), .CK(clk), .Q(ram[3758]) );
  DFF_X1 ram_reg_234__13_ ( .D(n9611), .CK(clk), .Q(ram[3757]) );
  DFF_X1 ram_reg_234__12_ ( .D(n9610), .CK(clk), .Q(ram[3756]) );
  DFF_X1 ram_reg_234__11_ ( .D(n9609), .CK(clk), .Q(ram[3755]) );
  DFF_X1 ram_reg_234__10_ ( .D(n9608), .CK(clk), .Q(ram[3754]) );
  DFF_X1 ram_reg_234__9_ ( .D(n9607), .CK(clk), .Q(ram[3753]) );
  DFF_X1 ram_reg_234__8_ ( .D(n9606), .CK(clk), .Q(ram[3752]) );
  DFF_X1 ram_reg_234__7_ ( .D(n9605), .CK(clk), .Q(ram[3751]) );
  DFF_X1 ram_reg_234__6_ ( .D(n9604), .CK(clk), .Q(ram[3750]) );
  DFF_X1 ram_reg_234__5_ ( .D(n9603), .CK(clk), .Q(ram[3749]) );
  DFF_X1 ram_reg_234__4_ ( .D(n9602), .CK(clk), .Q(ram[3748]) );
  DFF_X1 ram_reg_234__3_ ( .D(n9601), .CK(clk), .Q(ram[3747]) );
  DFF_X1 ram_reg_234__2_ ( .D(n9600), .CK(clk), .Q(ram[3746]) );
  DFF_X1 ram_reg_234__1_ ( .D(n9599), .CK(clk), .Q(ram[3745]) );
  DFF_X1 ram_reg_234__0_ ( .D(n9598), .CK(clk), .Q(ram[3744]) );
  DFF_X1 ram_reg_233__15_ ( .D(n9630), .CK(clk), .Q(ram[3743]) );
  DFF_X1 ram_reg_233__14_ ( .D(n9629), .CK(clk), .Q(ram[3742]) );
  DFF_X1 ram_reg_233__13_ ( .D(n9628), .CK(clk), .Q(ram[3741]) );
  DFF_X1 ram_reg_233__12_ ( .D(n9627), .CK(clk), .Q(ram[3740]) );
  DFF_X1 ram_reg_233__11_ ( .D(n9626), .CK(clk), .Q(ram[3739]) );
  DFF_X1 ram_reg_233__10_ ( .D(n9625), .CK(clk), .Q(ram[3738]) );
  DFF_X1 ram_reg_233__9_ ( .D(n9624), .CK(clk), .Q(ram[3737]) );
  DFF_X1 ram_reg_233__8_ ( .D(n9623), .CK(clk), .Q(ram[3736]) );
  DFF_X1 ram_reg_233__7_ ( .D(n9622), .CK(clk), .Q(ram[3735]) );
  DFF_X1 ram_reg_233__6_ ( .D(n9621), .CK(clk), .Q(ram[3734]) );
  DFF_X1 ram_reg_233__5_ ( .D(n9620), .CK(clk), .Q(ram[3733]) );
  DFF_X1 ram_reg_233__4_ ( .D(n9619), .CK(clk), .Q(ram[3732]) );
  DFF_X1 ram_reg_233__3_ ( .D(n9618), .CK(clk), .Q(ram[3731]) );
  DFF_X1 ram_reg_233__2_ ( .D(n9617), .CK(clk), .Q(ram[3730]) );
  DFF_X1 ram_reg_233__1_ ( .D(n9616), .CK(clk), .Q(ram[3729]) );
  DFF_X1 ram_reg_233__0_ ( .D(n9615), .CK(clk), .Q(ram[3728]) );
  DFF_X1 ram_reg_232__15_ ( .D(n9647), .CK(clk), .Q(ram[3727]) );
  DFF_X1 ram_reg_232__14_ ( .D(n9646), .CK(clk), .Q(ram[3726]) );
  DFF_X1 ram_reg_232__13_ ( .D(n9645), .CK(clk), .Q(ram[3725]) );
  DFF_X1 ram_reg_232__12_ ( .D(n9644), .CK(clk), .Q(ram[3724]) );
  DFF_X1 ram_reg_232__11_ ( .D(n9643), .CK(clk), .Q(ram[3723]) );
  DFF_X1 ram_reg_232__10_ ( .D(n9642), .CK(clk), .Q(ram[3722]) );
  DFF_X1 ram_reg_232__9_ ( .D(n9641), .CK(clk), .Q(ram[3721]) );
  DFF_X1 ram_reg_232__8_ ( .D(n9640), .CK(clk), .Q(ram[3720]) );
  DFF_X1 ram_reg_232__7_ ( .D(n9639), .CK(clk), .Q(ram[3719]) );
  DFF_X1 ram_reg_232__6_ ( .D(n9638), .CK(clk), .Q(ram[3718]) );
  DFF_X1 ram_reg_232__5_ ( .D(n9637), .CK(clk), .Q(ram[3717]) );
  DFF_X1 ram_reg_232__4_ ( .D(n9636), .CK(clk), .Q(ram[3716]) );
  DFF_X1 ram_reg_232__3_ ( .D(n9635), .CK(clk), .Q(ram[3715]) );
  DFF_X1 ram_reg_232__2_ ( .D(n9634), .CK(clk), .Q(ram[3714]) );
  DFF_X1 ram_reg_232__1_ ( .D(n9633), .CK(clk), .Q(ram[3713]) );
  DFF_X1 ram_reg_232__0_ ( .D(n9632), .CK(clk), .Q(ram[3712]) );
  DFF_X1 ram_reg_231__15_ ( .D(n9664), .CK(clk), .Q(ram[3711]) );
  DFF_X1 ram_reg_231__14_ ( .D(n9663), .CK(clk), .Q(ram[3710]) );
  DFF_X1 ram_reg_231__13_ ( .D(n9662), .CK(clk), .Q(ram[3709]) );
  DFF_X1 ram_reg_231__12_ ( .D(n9661), .CK(clk), .Q(ram[3708]) );
  DFF_X1 ram_reg_231__11_ ( .D(n9660), .CK(clk), .Q(ram[3707]) );
  DFF_X1 ram_reg_231__10_ ( .D(n9659), .CK(clk), .Q(ram[3706]) );
  DFF_X1 ram_reg_231__9_ ( .D(n9658), .CK(clk), .Q(ram[3705]) );
  DFF_X1 ram_reg_231__8_ ( .D(n9657), .CK(clk), .Q(ram[3704]) );
  DFF_X1 ram_reg_231__7_ ( .D(n9656), .CK(clk), .Q(ram[3703]) );
  DFF_X1 ram_reg_231__6_ ( .D(n9655), .CK(clk), .Q(ram[3702]) );
  DFF_X1 ram_reg_231__5_ ( .D(n9654), .CK(clk), .Q(ram[3701]) );
  DFF_X1 ram_reg_231__4_ ( .D(n9653), .CK(clk), .Q(ram[3700]) );
  DFF_X1 ram_reg_231__3_ ( .D(n9652), .CK(clk), .Q(ram[3699]) );
  DFF_X1 ram_reg_231__2_ ( .D(n9651), .CK(clk), .Q(ram[3698]) );
  DFF_X1 ram_reg_231__1_ ( .D(n9650), .CK(clk), .Q(ram[3697]) );
  DFF_X1 ram_reg_231__0_ ( .D(n9649), .CK(clk), .Q(ram[3696]) );
  DFF_X1 ram_reg_230__15_ ( .D(n9681), .CK(clk), .Q(ram[3695]) );
  DFF_X1 ram_reg_230__14_ ( .D(n9680), .CK(clk), .Q(ram[3694]) );
  DFF_X1 ram_reg_230__13_ ( .D(n9679), .CK(clk), .Q(ram[3693]) );
  DFF_X1 ram_reg_230__12_ ( .D(n9678), .CK(clk), .Q(ram[3692]) );
  DFF_X1 ram_reg_230__11_ ( .D(n9677), .CK(clk), .Q(ram[3691]) );
  DFF_X1 ram_reg_230__10_ ( .D(n9676), .CK(clk), .Q(ram[3690]) );
  DFF_X1 ram_reg_230__9_ ( .D(n9675), .CK(clk), .Q(ram[3689]) );
  DFF_X1 ram_reg_230__8_ ( .D(n9674), .CK(clk), .Q(ram[3688]) );
  DFF_X1 ram_reg_230__7_ ( .D(n9673), .CK(clk), .Q(ram[3687]) );
  DFF_X1 ram_reg_230__6_ ( .D(n9672), .CK(clk), .Q(ram[3686]) );
  DFF_X1 ram_reg_230__5_ ( .D(n9671), .CK(clk), .Q(ram[3685]) );
  DFF_X1 ram_reg_230__4_ ( .D(n9670), .CK(clk), .Q(ram[3684]) );
  DFF_X1 ram_reg_230__3_ ( .D(n9669), .CK(clk), .Q(ram[3683]) );
  DFF_X1 ram_reg_230__2_ ( .D(n9668), .CK(clk), .Q(ram[3682]) );
  DFF_X1 ram_reg_230__1_ ( .D(n9667), .CK(clk), .Q(ram[3681]) );
  DFF_X1 ram_reg_230__0_ ( .D(n9666), .CK(clk), .Q(ram[3680]) );
  DFF_X1 ram_reg_229__15_ ( .D(n9698), .CK(clk), .Q(ram[3679]) );
  DFF_X1 ram_reg_229__14_ ( .D(n9697), .CK(clk), .Q(ram[3678]) );
  DFF_X1 ram_reg_229__13_ ( .D(n9696), .CK(clk), .Q(ram[3677]) );
  DFF_X1 ram_reg_229__12_ ( .D(n9695), .CK(clk), .Q(ram[3676]) );
  DFF_X1 ram_reg_229__11_ ( .D(n9694), .CK(clk), .Q(ram[3675]) );
  DFF_X1 ram_reg_229__10_ ( .D(n9693), .CK(clk), .Q(ram[3674]) );
  DFF_X1 ram_reg_229__9_ ( .D(n9692), .CK(clk), .Q(ram[3673]) );
  DFF_X1 ram_reg_229__8_ ( .D(n9691), .CK(clk), .Q(ram[3672]) );
  DFF_X1 ram_reg_229__7_ ( .D(n9690), .CK(clk), .Q(ram[3671]) );
  DFF_X1 ram_reg_229__6_ ( .D(n9689), .CK(clk), .Q(ram[3670]) );
  DFF_X1 ram_reg_229__5_ ( .D(n9688), .CK(clk), .Q(ram[3669]) );
  DFF_X1 ram_reg_229__4_ ( .D(n9687), .CK(clk), .Q(ram[3668]) );
  DFF_X1 ram_reg_229__3_ ( .D(n9686), .CK(clk), .Q(ram[3667]) );
  DFF_X1 ram_reg_229__2_ ( .D(n9685), .CK(clk), .Q(ram[3666]) );
  DFF_X1 ram_reg_229__1_ ( .D(n9684), .CK(clk), .Q(ram[3665]) );
  DFF_X1 ram_reg_229__0_ ( .D(n9683), .CK(clk), .Q(ram[3664]) );
  DFF_X1 ram_reg_228__15_ ( .D(n9715), .CK(clk), .Q(ram[3663]) );
  DFF_X1 ram_reg_228__14_ ( .D(n9714), .CK(clk), .Q(ram[3662]) );
  DFF_X1 ram_reg_228__13_ ( .D(n9713), .CK(clk), .Q(ram[3661]) );
  DFF_X1 ram_reg_228__12_ ( .D(n9712), .CK(clk), .Q(ram[3660]) );
  DFF_X1 ram_reg_228__11_ ( .D(n9711), .CK(clk), .Q(ram[3659]) );
  DFF_X1 ram_reg_228__10_ ( .D(n9710), .CK(clk), .Q(ram[3658]) );
  DFF_X1 ram_reg_228__9_ ( .D(n9709), .CK(clk), .Q(ram[3657]) );
  DFF_X1 ram_reg_228__8_ ( .D(n9708), .CK(clk), .Q(ram[3656]) );
  DFF_X1 ram_reg_228__7_ ( .D(n9707), .CK(clk), .Q(ram[3655]) );
  DFF_X1 ram_reg_228__6_ ( .D(n9706), .CK(clk), .Q(ram[3654]) );
  DFF_X1 ram_reg_228__5_ ( .D(n9705), .CK(clk), .Q(ram[3653]) );
  DFF_X1 ram_reg_228__4_ ( .D(n9704), .CK(clk), .Q(ram[3652]) );
  DFF_X1 ram_reg_228__3_ ( .D(n9703), .CK(clk), .Q(ram[3651]) );
  DFF_X1 ram_reg_228__2_ ( .D(n9702), .CK(clk), .Q(ram[3650]) );
  DFF_X1 ram_reg_228__1_ ( .D(n9701), .CK(clk), .Q(ram[3649]) );
  DFF_X1 ram_reg_228__0_ ( .D(n9700), .CK(clk), .Q(ram[3648]) );
  DFF_X1 ram_reg_227__15_ ( .D(n9732), .CK(clk), .Q(ram[3647]) );
  DFF_X1 ram_reg_227__14_ ( .D(n9731), .CK(clk), .Q(ram[3646]) );
  DFF_X1 ram_reg_227__13_ ( .D(n9730), .CK(clk), .Q(ram[3645]) );
  DFF_X1 ram_reg_227__12_ ( .D(n9729), .CK(clk), .Q(ram[3644]) );
  DFF_X1 ram_reg_227__11_ ( .D(n9728), .CK(clk), .Q(ram[3643]) );
  DFF_X1 ram_reg_227__10_ ( .D(n9727), .CK(clk), .Q(ram[3642]) );
  DFF_X1 ram_reg_227__9_ ( .D(n9726), .CK(clk), .Q(ram[3641]) );
  DFF_X1 ram_reg_227__8_ ( .D(n9725), .CK(clk), .Q(ram[3640]) );
  DFF_X1 ram_reg_227__7_ ( .D(n9724), .CK(clk), .Q(ram[3639]) );
  DFF_X1 ram_reg_227__6_ ( .D(n9723), .CK(clk), .Q(ram[3638]) );
  DFF_X1 ram_reg_227__5_ ( .D(n9722), .CK(clk), .Q(ram[3637]) );
  DFF_X1 ram_reg_227__4_ ( .D(n9721), .CK(clk), .Q(ram[3636]) );
  DFF_X1 ram_reg_227__3_ ( .D(n9720), .CK(clk), .Q(ram[3635]) );
  DFF_X1 ram_reg_227__2_ ( .D(n9719), .CK(clk), .Q(ram[3634]) );
  DFF_X1 ram_reg_227__1_ ( .D(n9718), .CK(clk), .Q(ram[3633]) );
  DFF_X1 ram_reg_227__0_ ( .D(n9717), .CK(clk), .Q(ram[3632]) );
  DFF_X1 ram_reg_226__15_ ( .D(n9749), .CK(clk), .Q(ram[3631]) );
  DFF_X1 ram_reg_226__14_ ( .D(n9748), .CK(clk), .Q(ram[3630]) );
  DFF_X1 ram_reg_226__13_ ( .D(n9747), .CK(clk), .Q(ram[3629]) );
  DFF_X1 ram_reg_226__12_ ( .D(n9746), .CK(clk), .Q(ram[3628]) );
  DFF_X1 ram_reg_226__11_ ( .D(n9745), .CK(clk), .Q(ram[3627]) );
  DFF_X1 ram_reg_226__10_ ( .D(n9744), .CK(clk), .Q(ram[3626]) );
  DFF_X1 ram_reg_226__9_ ( .D(n9743), .CK(clk), .Q(ram[3625]) );
  DFF_X1 ram_reg_226__8_ ( .D(n9742), .CK(clk), .Q(ram[3624]) );
  DFF_X1 ram_reg_226__7_ ( .D(n9741), .CK(clk), .Q(ram[3623]) );
  DFF_X1 ram_reg_226__6_ ( .D(n9740), .CK(clk), .Q(ram[3622]) );
  DFF_X1 ram_reg_226__5_ ( .D(n9739), .CK(clk), .Q(ram[3621]) );
  DFF_X1 ram_reg_226__4_ ( .D(n9738), .CK(clk), .Q(ram[3620]) );
  DFF_X1 ram_reg_226__3_ ( .D(n9737), .CK(clk), .Q(ram[3619]) );
  DFF_X1 ram_reg_226__2_ ( .D(n9736), .CK(clk), .Q(ram[3618]) );
  DFF_X1 ram_reg_226__1_ ( .D(n9735), .CK(clk), .Q(ram[3617]) );
  DFF_X1 ram_reg_226__0_ ( .D(n9734), .CK(clk), .Q(ram[3616]) );
  DFF_X1 ram_reg_225__15_ ( .D(n9766), .CK(clk), .Q(ram[3615]) );
  DFF_X1 ram_reg_225__14_ ( .D(n9765), .CK(clk), .Q(ram[3614]) );
  DFF_X1 ram_reg_225__13_ ( .D(n9764), .CK(clk), .Q(ram[3613]) );
  DFF_X1 ram_reg_225__12_ ( .D(n9763), .CK(clk), .Q(ram[3612]) );
  DFF_X1 ram_reg_225__11_ ( .D(n9762), .CK(clk), .Q(ram[3611]) );
  DFF_X1 ram_reg_225__10_ ( .D(n9761), .CK(clk), .Q(ram[3610]) );
  DFF_X1 ram_reg_225__9_ ( .D(n9760), .CK(clk), .Q(ram[3609]) );
  DFF_X1 ram_reg_225__8_ ( .D(n9759), .CK(clk), .Q(ram[3608]) );
  DFF_X1 ram_reg_225__7_ ( .D(n9758), .CK(clk), .Q(ram[3607]) );
  DFF_X1 ram_reg_225__6_ ( .D(n9757), .CK(clk), .Q(ram[3606]) );
  DFF_X1 ram_reg_225__5_ ( .D(n9756), .CK(clk), .Q(ram[3605]) );
  DFF_X1 ram_reg_225__4_ ( .D(n9755), .CK(clk), .Q(ram[3604]) );
  DFF_X1 ram_reg_225__3_ ( .D(n9754), .CK(clk), .Q(ram[3603]) );
  DFF_X1 ram_reg_225__2_ ( .D(n9753), .CK(clk), .Q(ram[3602]) );
  DFF_X1 ram_reg_225__1_ ( .D(n9752), .CK(clk), .Q(ram[3601]) );
  DFF_X1 ram_reg_225__0_ ( .D(n9751), .CK(clk), .Q(ram[3600]) );
  DFF_X1 ram_reg_224__15_ ( .D(n9783), .CK(clk), .Q(ram[3599]) );
  DFF_X1 ram_reg_224__14_ ( .D(n9782), .CK(clk), .Q(ram[3598]) );
  DFF_X1 ram_reg_224__13_ ( .D(n9781), .CK(clk), .Q(ram[3597]) );
  DFF_X1 ram_reg_224__12_ ( .D(n9780), .CK(clk), .Q(ram[3596]) );
  DFF_X1 ram_reg_224__11_ ( .D(n9779), .CK(clk), .Q(ram[3595]) );
  DFF_X1 ram_reg_224__10_ ( .D(n9778), .CK(clk), .Q(ram[3594]) );
  DFF_X1 ram_reg_224__9_ ( .D(n9777), .CK(clk), .Q(ram[3593]) );
  DFF_X1 ram_reg_224__8_ ( .D(n9776), .CK(clk), .Q(ram[3592]) );
  DFF_X1 ram_reg_224__7_ ( .D(n9775), .CK(clk), .Q(ram[3591]) );
  DFF_X1 ram_reg_224__6_ ( .D(n9774), .CK(clk), .Q(ram[3590]) );
  DFF_X1 ram_reg_224__5_ ( .D(n9773), .CK(clk), .Q(ram[3589]) );
  DFF_X1 ram_reg_224__4_ ( .D(n9772), .CK(clk), .Q(ram[3588]) );
  DFF_X1 ram_reg_224__3_ ( .D(n9771), .CK(clk), .Q(ram[3587]) );
  DFF_X1 ram_reg_224__2_ ( .D(n9770), .CK(clk), .Q(ram[3586]) );
  DFF_X1 ram_reg_224__1_ ( .D(n9769), .CK(clk), .Q(ram[3585]) );
  DFF_X1 ram_reg_224__0_ ( .D(n9768), .CK(clk), .Q(ram[3584]) );
  DFF_X1 ram_reg_223__15_ ( .D(n9800), .CK(clk), .Q(ram[3583]) );
  DFF_X1 ram_reg_223__14_ ( .D(n9799), .CK(clk), .Q(ram[3582]) );
  DFF_X1 ram_reg_223__13_ ( .D(n9798), .CK(clk), .Q(ram[3581]) );
  DFF_X1 ram_reg_223__12_ ( .D(n9797), .CK(clk), .Q(ram[3580]) );
  DFF_X1 ram_reg_223__11_ ( .D(n9796), .CK(clk), .Q(ram[3579]) );
  DFF_X1 ram_reg_223__10_ ( .D(n9795), .CK(clk), .Q(ram[3578]) );
  DFF_X1 ram_reg_223__9_ ( .D(n9794), .CK(clk), .Q(ram[3577]) );
  DFF_X1 ram_reg_223__8_ ( .D(n9793), .CK(clk), .Q(ram[3576]) );
  DFF_X1 ram_reg_223__7_ ( .D(n9792), .CK(clk), .Q(ram[3575]) );
  DFF_X1 ram_reg_223__6_ ( .D(n9791), .CK(clk), .Q(ram[3574]) );
  DFF_X1 ram_reg_223__5_ ( .D(n9790), .CK(clk), .Q(ram[3573]) );
  DFF_X1 ram_reg_223__4_ ( .D(n9789), .CK(clk), .Q(ram[3572]) );
  DFF_X1 ram_reg_223__3_ ( .D(n9788), .CK(clk), .Q(ram[3571]) );
  DFF_X1 ram_reg_223__2_ ( .D(n9787), .CK(clk), .Q(ram[3570]) );
  DFF_X1 ram_reg_223__1_ ( .D(n9786), .CK(clk), .Q(ram[3569]) );
  DFF_X1 ram_reg_223__0_ ( .D(n9785), .CK(clk), .Q(ram[3568]) );
  DFF_X1 ram_reg_222__15_ ( .D(n9817), .CK(clk), .Q(ram[3567]) );
  DFF_X1 ram_reg_222__14_ ( .D(n9816), .CK(clk), .Q(ram[3566]) );
  DFF_X1 ram_reg_222__13_ ( .D(n9815), .CK(clk), .Q(ram[3565]) );
  DFF_X1 ram_reg_222__12_ ( .D(n9814), .CK(clk), .Q(ram[3564]) );
  DFF_X1 ram_reg_222__11_ ( .D(n9813), .CK(clk), .Q(ram[3563]) );
  DFF_X1 ram_reg_222__10_ ( .D(n9812), .CK(clk), .Q(ram[3562]) );
  DFF_X1 ram_reg_222__9_ ( .D(n9811), .CK(clk), .Q(ram[3561]) );
  DFF_X1 ram_reg_222__8_ ( .D(n9810), .CK(clk), .Q(ram[3560]) );
  DFF_X1 ram_reg_222__7_ ( .D(n9809), .CK(clk), .Q(ram[3559]) );
  DFF_X1 ram_reg_222__6_ ( .D(n9808), .CK(clk), .Q(ram[3558]) );
  DFF_X1 ram_reg_222__5_ ( .D(n9807), .CK(clk), .Q(ram[3557]) );
  DFF_X1 ram_reg_222__4_ ( .D(n9806), .CK(clk), .Q(ram[3556]) );
  DFF_X1 ram_reg_222__3_ ( .D(n9805), .CK(clk), .Q(ram[3555]) );
  DFF_X1 ram_reg_222__2_ ( .D(n9804), .CK(clk), .Q(ram[3554]) );
  DFF_X1 ram_reg_222__1_ ( .D(n9803), .CK(clk), .Q(ram[3553]) );
  DFF_X1 ram_reg_222__0_ ( .D(n9802), .CK(clk), .Q(ram[3552]) );
  DFF_X1 ram_reg_221__15_ ( .D(n9834), .CK(clk), .Q(ram[3551]) );
  DFF_X1 ram_reg_221__14_ ( .D(n9833), .CK(clk), .Q(ram[3550]) );
  DFF_X1 ram_reg_221__13_ ( .D(n9832), .CK(clk), .Q(ram[3549]) );
  DFF_X1 ram_reg_221__12_ ( .D(n9831), .CK(clk), .Q(ram[3548]) );
  DFF_X1 ram_reg_221__11_ ( .D(n9830), .CK(clk), .Q(ram[3547]) );
  DFF_X1 ram_reg_221__10_ ( .D(n9829), .CK(clk), .Q(ram[3546]) );
  DFF_X1 ram_reg_221__9_ ( .D(n9828), .CK(clk), .Q(ram[3545]) );
  DFF_X1 ram_reg_221__8_ ( .D(n9827), .CK(clk), .Q(ram[3544]) );
  DFF_X1 ram_reg_221__7_ ( .D(n9826), .CK(clk), .Q(ram[3543]) );
  DFF_X1 ram_reg_221__6_ ( .D(n9825), .CK(clk), .Q(ram[3542]) );
  DFF_X1 ram_reg_221__5_ ( .D(n9824), .CK(clk), .Q(ram[3541]) );
  DFF_X1 ram_reg_221__4_ ( .D(n9823), .CK(clk), .Q(ram[3540]) );
  DFF_X1 ram_reg_221__3_ ( .D(n9822), .CK(clk), .Q(ram[3539]) );
  DFF_X1 ram_reg_221__2_ ( .D(n9821), .CK(clk), .Q(ram[3538]) );
  DFF_X1 ram_reg_221__1_ ( .D(n9820), .CK(clk), .Q(ram[3537]) );
  DFF_X1 ram_reg_221__0_ ( .D(n9819), .CK(clk), .Q(ram[3536]) );
  DFF_X1 ram_reg_220__15_ ( .D(n9851), .CK(clk), .Q(ram[3535]) );
  DFF_X1 ram_reg_220__14_ ( .D(n9850), .CK(clk), .Q(ram[3534]) );
  DFF_X1 ram_reg_220__13_ ( .D(n9849), .CK(clk), .Q(ram[3533]) );
  DFF_X1 ram_reg_220__12_ ( .D(n9848), .CK(clk), .Q(ram[3532]) );
  DFF_X1 ram_reg_220__11_ ( .D(n9847), .CK(clk), .Q(ram[3531]) );
  DFF_X1 ram_reg_220__10_ ( .D(n9846), .CK(clk), .Q(ram[3530]) );
  DFF_X1 ram_reg_220__9_ ( .D(n9845), .CK(clk), .Q(ram[3529]) );
  DFF_X1 ram_reg_220__8_ ( .D(n9844), .CK(clk), .Q(ram[3528]) );
  DFF_X1 ram_reg_220__7_ ( .D(n9843), .CK(clk), .Q(ram[3527]) );
  DFF_X1 ram_reg_220__6_ ( .D(n9842), .CK(clk), .Q(ram[3526]) );
  DFF_X1 ram_reg_220__5_ ( .D(n9841), .CK(clk), .Q(ram[3525]) );
  DFF_X1 ram_reg_220__4_ ( .D(n9840), .CK(clk), .Q(ram[3524]) );
  DFF_X1 ram_reg_220__3_ ( .D(n9839), .CK(clk), .Q(ram[3523]) );
  DFF_X1 ram_reg_220__2_ ( .D(n9838), .CK(clk), .Q(ram[3522]) );
  DFF_X1 ram_reg_220__1_ ( .D(n9837), .CK(clk), .Q(ram[3521]) );
  DFF_X1 ram_reg_220__0_ ( .D(n9836), .CK(clk), .Q(ram[3520]) );
  DFF_X1 ram_reg_219__15_ ( .D(n9868), .CK(clk), .Q(ram[3519]) );
  DFF_X1 ram_reg_219__14_ ( .D(n9867), .CK(clk), .Q(ram[3518]) );
  DFF_X1 ram_reg_219__13_ ( .D(n9866), .CK(clk), .Q(ram[3517]) );
  DFF_X1 ram_reg_219__12_ ( .D(n9865), .CK(clk), .Q(ram[3516]) );
  DFF_X1 ram_reg_219__11_ ( .D(n9864), .CK(clk), .Q(ram[3515]) );
  DFF_X1 ram_reg_219__10_ ( .D(n9863), .CK(clk), .Q(ram[3514]) );
  DFF_X1 ram_reg_219__9_ ( .D(n9862), .CK(clk), .Q(ram[3513]) );
  DFF_X1 ram_reg_219__8_ ( .D(n9861), .CK(clk), .Q(ram[3512]) );
  DFF_X1 ram_reg_219__7_ ( .D(n9860), .CK(clk), .Q(ram[3511]) );
  DFF_X1 ram_reg_219__6_ ( .D(n9859), .CK(clk), .Q(ram[3510]) );
  DFF_X1 ram_reg_219__5_ ( .D(n9858), .CK(clk), .Q(ram[3509]) );
  DFF_X1 ram_reg_219__4_ ( .D(n9857), .CK(clk), .Q(ram[3508]) );
  DFF_X1 ram_reg_219__3_ ( .D(n9856), .CK(clk), .Q(ram[3507]) );
  DFF_X1 ram_reg_219__2_ ( .D(n9855), .CK(clk), .Q(ram[3506]) );
  DFF_X1 ram_reg_219__1_ ( .D(n9854), .CK(clk), .Q(ram[3505]) );
  DFF_X1 ram_reg_219__0_ ( .D(n9853), .CK(clk), .Q(ram[3504]) );
  DFF_X1 ram_reg_218__15_ ( .D(n9885), .CK(clk), .Q(ram[3503]) );
  DFF_X1 ram_reg_218__14_ ( .D(n9884), .CK(clk), .Q(ram[3502]) );
  DFF_X1 ram_reg_218__13_ ( .D(n9883), .CK(clk), .Q(ram[3501]) );
  DFF_X1 ram_reg_218__12_ ( .D(n9882), .CK(clk), .Q(ram[3500]) );
  DFF_X1 ram_reg_218__11_ ( .D(n9881), .CK(clk), .Q(ram[3499]) );
  DFF_X1 ram_reg_218__10_ ( .D(n9880), .CK(clk), .Q(ram[3498]) );
  DFF_X1 ram_reg_218__9_ ( .D(n9879), .CK(clk), .Q(ram[3497]) );
  DFF_X1 ram_reg_218__8_ ( .D(n9878), .CK(clk), .Q(ram[3496]) );
  DFF_X1 ram_reg_218__7_ ( .D(n9877), .CK(clk), .Q(ram[3495]) );
  DFF_X1 ram_reg_218__6_ ( .D(n9876), .CK(clk), .Q(ram[3494]) );
  DFF_X1 ram_reg_218__5_ ( .D(n9875), .CK(clk), .Q(ram[3493]) );
  DFF_X1 ram_reg_218__4_ ( .D(n9874), .CK(clk), .Q(ram[3492]) );
  DFF_X1 ram_reg_218__3_ ( .D(n9873), .CK(clk), .Q(ram[3491]) );
  DFF_X1 ram_reg_218__2_ ( .D(n9872), .CK(clk), .Q(ram[3490]) );
  DFF_X1 ram_reg_218__1_ ( .D(n9871), .CK(clk), .Q(ram[3489]) );
  DFF_X1 ram_reg_218__0_ ( .D(n9870), .CK(clk), .Q(ram[3488]) );
  DFF_X1 ram_reg_217__15_ ( .D(n9902), .CK(clk), .Q(ram[3487]) );
  DFF_X1 ram_reg_217__14_ ( .D(n9901), .CK(clk), .Q(ram[3486]) );
  DFF_X1 ram_reg_217__13_ ( .D(n9900), .CK(clk), .Q(ram[3485]) );
  DFF_X1 ram_reg_217__12_ ( .D(n9899), .CK(clk), .Q(ram[3484]) );
  DFF_X1 ram_reg_217__11_ ( .D(n9898), .CK(clk), .Q(ram[3483]) );
  DFF_X1 ram_reg_217__10_ ( .D(n9897), .CK(clk), .Q(ram[3482]) );
  DFF_X1 ram_reg_217__9_ ( .D(n9896), .CK(clk), .Q(ram[3481]) );
  DFF_X1 ram_reg_217__8_ ( .D(n9895), .CK(clk), .Q(ram[3480]) );
  DFF_X1 ram_reg_217__7_ ( .D(n9894), .CK(clk), .Q(ram[3479]) );
  DFF_X1 ram_reg_217__6_ ( .D(n9893), .CK(clk), .Q(ram[3478]) );
  DFF_X1 ram_reg_217__5_ ( .D(n9892), .CK(clk), .Q(ram[3477]) );
  DFF_X1 ram_reg_217__4_ ( .D(n9891), .CK(clk), .Q(ram[3476]) );
  DFF_X1 ram_reg_217__3_ ( .D(n9890), .CK(clk), .Q(ram[3475]) );
  DFF_X1 ram_reg_217__2_ ( .D(n9889), .CK(clk), .Q(ram[3474]) );
  DFF_X1 ram_reg_217__1_ ( .D(n9888), .CK(clk), .Q(ram[3473]) );
  DFF_X1 ram_reg_217__0_ ( .D(n9887), .CK(clk), .Q(ram[3472]) );
  DFF_X1 ram_reg_216__15_ ( .D(n9919), .CK(clk), .Q(ram[3471]) );
  DFF_X1 ram_reg_216__14_ ( .D(n9918), .CK(clk), .Q(ram[3470]) );
  DFF_X1 ram_reg_216__13_ ( .D(n9917), .CK(clk), .Q(ram[3469]) );
  DFF_X1 ram_reg_216__12_ ( .D(n9916), .CK(clk), .Q(ram[3468]) );
  DFF_X1 ram_reg_216__11_ ( .D(n9915), .CK(clk), .Q(ram[3467]) );
  DFF_X1 ram_reg_216__10_ ( .D(n9914), .CK(clk), .Q(ram[3466]) );
  DFF_X1 ram_reg_216__9_ ( .D(n9913), .CK(clk), .Q(ram[3465]) );
  DFF_X1 ram_reg_216__8_ ( .D(n9912), .CK(clk), .Q(ram[3464]) );
  DFF_X1 ram_reg_216__7_ ( .D(n9911), .CK(clk), .Q(ram[3463]) );
  DFF_X1 ram_reg_216__6_ ( .D(n9910), .CK(clk), .Q(ram[3462]) );
  DFF_X1 ram_reg_216__5_ ( .D(n9909), .CK(clk), .Q(ram[3461]) );
  DFF_X1 ram_reg_216__4_ ( .D(n9908), .CK(clk), .Q(ram[3460]) );
  DFF_X1 ram_reg_216__3_ ( .D(n9907), .CK(clk), .Q(ram[3459]) );
  DFF_X1 ram_reg_216__2_ ( .D(n9906), .CK(clk), .Q(ram[3458]) );
  DFF_X1 ram_reg_216__1_ ( .D(n9905), .CK(clk), .Q(ram[3457]) );
  DFF_X1 ram_reg_216__0_ ( .D(n9904), .CK(clk), .Q(ram[3456]) );
  DFF_X1 ram_reg_215__15_ ( .D(n9936), .CK(clk), .Q(ram[3455]) );
  DFF_X1 ram_reg_215__14_ ( .D(n9935), .CK(clk), .Q(ram[3454]) );
  DFF_X1 ram_reg_215__13_ ( .D(n9934), .CK(clk), .Q(ram[3453]) );
  DFF_X1 ram_reg_215__12_ ( .D(n9933), .CK(clk), .Q(ram[3452]) );
  DFF_X1 ram_reg_215__11_ ( .D(n9932), .CK(clk), .Q(ram[3451]) );
  DFF_X1 ram_reg_215__10_ ( .D(n9931), .CK(clk), .Q(ram[3450]) );
  DFF_X1 ram_reg_215__9_ ( .D(n9930), .CK(clk), .Q(ram[3449]) );
  DFF_X1 ram_reg_215__8_ ( .D(n9929), .CK(clk), .Q(ram[3448]) );
  DFF_X1 ram_reg_215__7_ ( .D(n9928), .CK(clk), .Q(ram[3447]) );
  DFF_X1 ram_reg_215__6_ ( .D(n9927), .CK(clk), .Q(ram[3446]) );
  DFF_X1 ram_reg_215__5_ ( .D(n9926), .CK(clk), .Q(ram[3445]) );
  DFF_X1 ram_reg_215__4_ ( .D(n9925), .CK(clk), .Q(ram[3444]) );
  DFF_X1 ram_reg_215__3_ ( .D(n9924), .CK(clk), .Q(ram[3443]) );
  DFF_X1 ram_reg_215__2_ ( .D(n9923), .CK(clk), .Q(ram[3442]) );
  DFF_X1 ram_reg_215__1_ ( .D(n9922), .CK(clk), .Q(ram[3441]) );
  DFF_X1 ram_reg_215__0_ ( .D(n9921), .CK(clk), .Q(ram[3440]) );
  DFF_X1 ram_reg_214__15_ ( .D(n9953), .CK(clk), .Q(ram[3439]) );
  DFF_X1 ram_reg_214__14_ ( .D(n9952), .CK(clk), .Q(ram[3438]) );
  DFF_X1 ram_reg_214__13_ ( .D(n9951), .CK(clk), .Q(ram[3437]) );
  DFF_X1 ram_reg_214__12_ ( .D(n9950), .CK(clk), .Q(ram[3436]) );
  DFF_X1 ram_reg_214__11_ ( .D(n9949), .CK(clk), .Q(ram[3435]) );
  DFF_X1 ram_reg_214__10_ ( .D(n9948), .CK(clk), .Q(ram[3434]) );
  DFF_X1 ram_reg_214__9_ ( .D(n9947), .CK(clk), .Q(ram[3433]) );
  DFF_X1 ram_reg_214__8_ ( .D(n9946), .CK(clk), .Q(ram[3432]) );
  DFF_X1 ram_reg_214__7_ ( .D(n9945), .CK(clk), .Q(ram[3431]) );
  DFF_X1 ram_reg_214__6_ ( .D(n9944), .CK(clk), .Q(ram[3430]) );
  DFF_X1 ram_reg_214__5_ ( .D(n9943), .CK(clk), .Q(ram[3429]) );
  DFF_X1 ram_reg_214__4_ ( .D(n9942), .CK(clk), .Q(ram[3428]) );
  DFF_X1 ram_reg_214__3_ ( .D(n9941), .CK(clk), .Q(ram[3427]) );
  DFF_X1 ram_reg_214__2_ ( .D(n9940), .CK(clk), .Q(ram[3426]) );
  DFF_X1 ram_reg_214__1_ ( .D(n9939), .CK(clk), .Q(ram[3425]) );
  DFF_X1 ram_reg_214__0_ ( .D(n9938), .CK(clk), .Q(ram[3424]) );
  DFF_X1 ram_reg_213__15_ ( .D(n9970), .CK(clk), .Q(ram[3423]) );
  DFF_X1 ram_reg_213__14_ ( .D(n9969), .CK(clk), .Q(ram[3422]) );
  DFF_X1 ram_reg_213__13_ ( .D(n9968), .CK(clk), .Q(ram[3421]) );
  DFF_X1 ram_reg_213__12_ ( .D(n9967), .CK(clk), .Q(ram[3420]) );
  DFF_X1 ram_reg_213__11_ ( .D(n9966), .CK(clk), .Q(ram[3419]) );
  DFF_X1 ram_reg_213__10_ ( .D(n9965), .CK(clk), .Q(ram[3418]) );
  DFF_X1 ram_reg_213__9_ ( .D(n9964), .CK(clk), .Q(ram[3417]) );
  DFF_X1 ram_reg_213__8_ ( .D(n9963), .CK(clk), .Q(ram[3416]) );
  DFF_X1 ram_reg_213__7_ ( .D(n9962), .CK(clk), .Q(ram[3415]) );
  DFF_X1 ram_reg_213__6_ ( .D(n9961), .CK(clk), .Q(ram[3414]) );
  DFF_X1 ram_reg_213__5_ ( .D(n9960), .CK(clk), .Q(ram[3413]) );
  DFF_X1 ram_reg_213__4_ ( .D(n9959), .CK(clk), .Q(ram[3412]) );
  DFF_X1 ram_reg_213__3_ ( .D(n9958), .CK(clk), .Q(ram[3411]) );
  DFF_X1 ram_reg_213__2_ ( .D(n9957), .CK(clk), .Q(ram[3410]) );
  DFF_X1 ram_reg_213__1_ ( .D(n9956), .CK(clk), .Q(ram[3409]) );
  DFF_X1 ram_reg_213__0_ ( .D(n9955), .CK(clk), .Q(ram[3408]) );
  DFF_X1 ram_reg_212__15_ ( .D(n9987), .CK(clk), .Q(ram[3407]) );
  DFF_X1 ram_reg_212__14_ ( .D(n9986), .CK(clk), .Q(ram[3406]) );
  DFF_X1 ram_reg_212__13_ ( .D(n9985), .CK(clk), .Q(ram[3405]) );
  DFF_X1 ram_reg_212__12_ ( .D(n9984), .CK(clk), .Q(ram[3404]) );
  DFF_X1 ram_reg_212__11_ ( .D(n9983), .CK(clk), .Q(ram[3403]) );
  DFF_X1 ram_reg_212__10_ ( .D(n9982), .CK(clk), .Q(ram[3402]) );
  DFF_X1 ram_reg_212__9_ ( .D(n9981), .CK(clk), .Q(ram[3401]) );
  DFF_X1 ram_reg_212__8_ ( .D(n9980), .CK(clk), .Q(ram[3400]) );
  DFF_X1 ram_reg_212__7_ ( .D(n9979), .CK(clk), .Q(ram[3399]) );
  DFF_X1 ram_reg_212__6_ ( .D(n9978), .CK(clk), .Q(ram[3398]) );
  DFF_X1 ram_reg_212__5_ ( .D(n9977), .CK(clk), .Q(ram[3397]) );
  DFF_X1 ram_reg_212__4_ ( .D(n9976), .CK(clk), .Q(ram[3396]) );
  DFF_X1 ram_reg_212__3_ ( .D(n9975), .CK(clk), .Q(ram[3395]) );
  DFF_X1 ram_reg_212__2_ ( .D(n9974), .CK(clk), .Q(ram[3394]) );
  DFF_X1 ram_reg_212__1_ ( .D(n9973), .CK(clk), .Q(ram[3393]) );
  DFF_X1 ram_reg_212__0_ ( .D(n9972), .CK(clk), .Q(ram[3392]) );
  DFF_X1 ram_reg_211__15_ ( .D(n10004), .CK(clk), .Q(ram[3391]) );
  DFF_X1 ram_reg_211__14_ ( .D(n10003), .CK(clk), .Q(ram[3390]) );
  DFF_X1 ram_reg_211__13_ ( .D(n10002), .CK(clk), .Q(ram[3389]) );
  DFF_X1 ram_reg_211__12_ ( .D(n10001), .CK(clk), .Q(ram[3388]) );
  DFF_X1 ram_reg_211__11_ ( .D(n10000), .CK(clk), .Q(ram[3387]) );
  DFF_X1 ram_reg_211__10_ ( .D(n9999), .CK(clk), .Q(ram[3386]) );
  DFF_X1 ram_reg_211__9_ ( .D(n9998), .CK(clk), .Q(ram[3385]) );
  DFF_X1 ram_reg_211__8_ ( .D(n9997), .CK(clk), .Q(ram[3384]) );
  DFF_X1 ram_reg_211__7_ ( .D(n9996), .CK(clk), .Q(ram[3383]) );
  DFF_X1 ram_reg_211__6_ ( .D(n9995), .CK(clk), .Q(ram[3382]) );
  DFF_X1 ram_reg_211__5_ ( .D(n9994), .CK(clk), .Q(ram[3381]) );
  DFF_X1 ram_reg_211__4_ ( .D(n9993), .CK(clk), .Q(ram[3380]) );
  DFF_X1 ram_reg_211__3_ ( .D(n9992), .CK(clk), .Q(ram[3379]) );
  DFF_X1 ram_reg_211__2_ ( .D(n9991), .CK(clk), .Q(ram[3378]) );
  DFF_X1 ram_reg_211__1_ ( .D(n9990), .CK(clk), .Q(ram[3377]) );
  DFF_X1 ram_reg_211__0_ ( .D(n9989), .CK(clk), .Q(ram[3376]) );
  DFF_X1 ram_reg_210__15_ ( .D(n10021), .CK(clk), .Q(ram[3375]) );
  DFF_X1 ram_reg_210__14_ ( .D(n10020), .CK(clk), .Q(ram[3374]) );
  DFF_X1 ram_reg_210__13_ ( .D(n10019), .CK(clk), .Q(ram[3373]) );
  DFF_X1 ram_reg_210__12_ ( .D(n10018), .CK(clk), .Q(ram[3372]) );
  DFF_X1 ram_reg_210__11_ ( .D(n10017), .CK(clk), .Q(ram[3371]) );
  DFF_X1 ram_reg_210__10_ ( .D(n10016), .CK(clk), .Q(ram[3370]) );
  DFF_X1 ram_reg_210__9_ ( .D(n10015), .CK(clk), .Q(ram[3369]) );
  DFF_X1 ram_reg_210__8_ ( .D(n10014), .CK(clk), .Q(ram[3368]) );
  DFF_X1 ram_reg_210__7_ ( .D(n10013), .CK(clk), .Q(ram[3367]) );
  DFF_X1 ram_reg_210__6_ ( .D(n10012), .CK(clk), .Q(ram[3366]) );
  DFF_X1 ram_reg_210__5_ ( .D(n10011), .CK(clk), .Q(ram[3365]) );
  DFF_X1 ram_reg_210__4_ ( .D(n10010), .CK(clk), .Q(ram[3364]) );
  DFF_X1 ram_reg_210__3_ ( .D(n10009), .CK(clk), .Q(ram[3363]) );
  DFF_X1 ram_reg_210__2_ ( .D(n10008), .CK(clk), .Q(ram[3362]) );
  DFF_X1 ram_reg_210__1_ ( .D(n10007), .CK(clk), .Q(ram[3361]) );
  DFF_X1 ram_reg_210__0_ ( .D(n10006), .CK(clk), .Q(ram[3360]) );
  DFF_X1 ram_reg_209__15_ ( .D(n10038), .CK(clk), .Q(ram[3359]) );
  DFF_X1 ram_reg_209__14_ ( .D(n10037), .CK(clk), .Q(ram[3358]) );
  DFF_X1 ram_reg_209__13_ ( .D(n10036), .CK(clk), .Q(ram[3357]) );
  DFF_X1 ram_reg_209__12_ ( .D(n10035), .CK(clk), .Q(ram[3356]) );
  DFF_X1 ram_reg_209__11_ ( .D(n10034), .CK(clk), .Q(ram[3355]) );
  DFF_X1 ram_reg_209__10_ ( .D(n10033), .CK(clk), .Q(ram[3354]) );
  DFF_X1 ram_reg_209__9_ ( .D(n10032), .CK(clk), .Q(ram[3353]) );
  DFF_X1 ram_reg_209__8_ ( .D(n10031), .CK(clk), .Q(ram[3352]) );
  DFF_X1 ram_reg_209__7_ ( .D(n10030), .CK(clk), .Q(ram[3351]) );
  DFF_X1 ram_reg_209__6_ ( .D(n10029), .CK(clk), .Q(ram[3350]) );
  DFF_X1 ram_reg_209__5_ ( .D(n10028), .CK(clk), .Q(ram[3349]) );
  DFF_X1 ram_reg_209__4_ ( .D(n10027), .CK(clk), .Q(ram[3348]) );
  DFF_X1 ram_reg_209__3_ ( .D(n10026), .CK(clk), .Q(ram[3347]) );
  DFF_X1 ram_reg_209__2_ ( .D(n10025), .CK(clk), .Q(ram[3346]) );
  DFF_X1 ram_reg_209__1_ ( .D(n10024), .CK(clk), .Q(ram[3345]) );
  DFF_X1 ram_reg_209__0_ ( .D(n10023), .CK(clk), .Q(ram[3344]) );
  DFF_X1 ram_reg_208__15_ ( .D(n10055), .CK(clk), .Q(ram[3343]) );
  DFF_X1 ram_reg_208__14_ ( .D(n10054), .CK(clk), .Q(ram[3342]) );
  DFF_X1 ram_reg_208__13_ ( .D(n10053), .CK(clk), .Q(ram[3341]) );
  DFF_X1 ram_reg_208__12_ ( .D(n10052), .CK(clk), .Q(ram[3340]) );
  DFF_X1 ram_reg_208__11_ ( .D(n10051), .CK(clk), .Q(ram[3339]) );
  DFF_X1 ram_reg_208__10_ ( .D(n10050), .CK(clk), .Q(ram[3338]) );
  DFF_X1 ram_reg_208__9_ ( .D(n10049), .CK(clk), .Q(ram[3337]) );
  DFF_X1 ram_reg_208__8_ ( .D(n10048), .CK(clk), .Q(ram[3336]) );
  DFF_X1 ram_reg_208__7_ ( .D(n10047), .CK(clk), .Q(ram[3335]) );
  DFF_X1 ram_reg_208__6_ ( .D(n10046), .CK(clk), .Q(ram[3334]) );
  DFF_X1 ram_reg_208__5_ ( .D(n10045), .CK(clk), .Q(ram[3333]) );
  DFF_X1 ram_reg_208__4_ ( .D(n10044), .CK(clk), .Q(ram[3332]) );
  DFF_X1 ram_reg_208__3_ ( .D(n10043), .CK(clk), .Q(ram[3331]) );
  DFF_X1 ram_reg_208__2_ ( .D(n10042), .CK(clk), .Q(ram[3330]) );
  DFF_X1 ram_reg_208__1_ ( .D(n10041), .CK(clk), .Q(ram[3329]) );
  DFF_X1 ram_reg_208__0_ ( .D(n10040), .CK(clk), .Q(ram[3328]) );
  DFF_X1 ram_reg_207__15_ ( .D(n10072), .CK(clk), .Q(ram[3327]) );
  DFF_X1 ram_reg_207__14_ ( .D(n10071), .CK(clk), .Q(ram[3326]) );
  DFF_X1 ram_reg_207__13_ ( .D(n10070), .CK(clk), .Q(ram[3325]) );
  DFF_X1 ram_reg_207__12_ ( .D(n10069), .CK(clk), .Q(ram[3324]) );
  DFF_X1 ram_reg_207__11_ ( .D(n10068), .CK(clk), .Q(ram[3323]) );
  DFF_X1 ram_reg_207__10_ ( .D(n10067), .CK(clk), .Q(ram[3322]) );
  DFF_X1 ram_reg_207__9_ ( .D(n10066), .CK(clk), .Q(ram[3321]) );
  DFF_X1 ram_reg_207__8_ ( .D(n10065), .CK(clk), .Q(ram[3320]) );
  DFF_X1 ram_reg_207__7_ ( .D(n10064), .CK(clk), .Q(ram[3319]) );
  DFF_X1 ram_reg_207__6_ ( .D(n10063), .CK(clk), .Q(ram[3318]) );
  DFF_X1 ram_reg_207__5_ ( .D(n10062), .CK(clk), .Q(ram[3317]) );
  DFF_X1 ram_reg_207__4_ ( .D(n10061), .CK(clk), .Q(ram[3316]) );
  DFF_X1 ram_reg_207__3_ ( .D(n10060), .CK(clk), .Q(ram[3315]) );
  DFF_X1 ram_reg_207__2_ ( .D(n10059), .CK(clk), .Q(ram[3314]) );
  DFF_X1 ram_reg_207__1_ ( .D(n10058), .CK(clk), .Q(ram[3313]) );
  DFF_X1 ram_reg_207__0_ ( .D(n10057), .CK(clk), .Q(ram[3312]) );
  DFF_X1 ram_reg_206__15_ ( .D(n10089), .CK(clk), .Q(ram[3311]) );
  DFF_X1 ram_reg_206__14_ ( .D(n10088), .CK(clk), .Q(ram[3310]) );
  DFF_X1 ram_reg_206__13_ ( .D(n10087), .CK(clk), .Q(ram[3309]) );
  DFF_X1 ram_reg_206__12_ ( .D(n10086), .CK(clk), .Q(ram[3308]) );
  DFF_X1 ram_reg_206__11_ ( .D(n10085), .CK(clk), .Q(ram[3307]) );
  DFF_X1 ram_reg_206__10_ ( .D(n10084), .CK(clk), .Q(ram[3306]) );
  DFF_X1 ram_reg_206__9_ ( .D(n10083), .CK(clk), .Q(ram[3305]) );
  DFF_X1 ram_reg_206__8_ ( .D(n10082), .CK(clk), .Q(ram[3304]) );
  DFF_X1 ram_reg_206__7_ ( .D(n10081), .CK(clk), .Q(ram[3303]) );
  DFF_X1 ram_reg_206__6_ ( .D(n10080), .CK(clk), .Q(ram[3302]) );
  DFF_X1 ram_reg_206__5_ ( .D(n10079), .CK(clk), .Q(ram[3301]) );
  DFF_X1 ram_reg_206__4_ ( .D(n10078), .CK(clk), .Q(ram[3300]) );
  DFF_X1 ram_reg_206__3_ ( .D(n10077), .CK(clk), .Q(ram[3299]) );
  DFF_X1 ram_reg_206__2_ ( .D(n10076), .CK(clk), .Q(ram[3298]) );
  DFF_X1 ram_reg_206__1_ ( .D(n10075), .CK(clk), .Q(ram[3297]) );
  DFF_X1 ram_reg_206__0_ ( .D(n10074), .CK(clk), .Q(ram[3296]) );
  DFF_X1 ram_reg_205__15_ ( .D(n10106), .CK(clk), .Q(ram[3295]) );
  DFF_X1 ram_reg_205__14_ ( .D(n10105), .CK(clk), .Q(ram[3294]) );
  DFF_X1 ram_reg_205__13_ ( .D(n10104), .CK(clk), .Q(ram[3293]) );
  DFF_X1 ram_reg_205__12_ ( .D(n10103), .CK(clk), .Q(ram[3292]) );
  DFF_X1 ram_reg_205__11_ ( .D(n10102), .CK(clk), .Q(ram[3291]) );
  DFF_X1 ram_reg_205__10_ ( .D(n10101), .CK(clk), .Q(ram[3290]) );
  DFF_X1 ram_reg_205__9_ ( .D(n10100), .CK(clk), .Q(ram[3289]) );
  DFF_X1 ram_reg_205__8_ ( .D(n10099), .CK(clk), .Q(ram[3288]) );
  DFF_X1 ram_reg_205__7_ ( .D(n10098), .CK(clk), .Q(ram[3287]) );
  DFF_X1 ram_reg_205__6_ ( .D(n10097), .CK(clk), .Q(ram[3286]) );
  DFF_X1 ram_reg_205__5_ ( .D(n10096), .CK(clk), .Q(ram[3285]) );
  DFF_X1 ram_reg_205__4_ ( .D(n10095), .CK(clk), .Q(ram[3284]) );
  DFF_X1 ram_reg_205__3_ ( .D(n10094), .CK(clk), .Q(ram[3283]) );
  DFF_X1 ram_reg_205__2_ ( .D(n10093), .CK(clk), .Q(ram[3282]) );
  DFF_X1 ram_reg_205__1_ ( .D(n10092), .CK(clk), .Q(ram[3281]) );
  DFF_X1 ram_reg_205__0_ ( .D(n10091), .CK(clk), .Q(ram[3280]) );
  DFF_X1 ram_reg_204__15_ ( .D(n10123), .CK(clk), .Q(ram[3279]) );
  DFF_X1 ram_reg_204__14_ ( .D(n10122), .CK(clk), .Q(ram[3278]) );
  DFF_X1 ram_reg_204__13_ ( .D(n10121), .CK(clk), .Q(ram[3277]) );
  DFF_X1 ram_reg_204__12_ ( .D(n10120), .CK(clk), .Q(ram[3276]) );
  DFF_X1 ram_reg_204__11_ ( .D(n10119), .CK(clk), .Q(ram[3275]) );
  DFF_X1 ram_reg_204__10_ ( .D(n10118), .CK(clk), .Q(ram[3274]) );
  DFF_X1 ram_reg_204__9_ ( .D(n10117), .CK(clk), .Q(ram[3273]) );
  DFF_X1 ram_reg_204__8_ ( .D(n10116), .CK(clk), .Q(ram[3272]) );
  DFF_X1 ram_reg_204__7_ ( .D(n10115), .CK(clk), .Q(ram[3271]) );
  DFF_X1 ram_reg_204__6_ ( .D(n10114), .CK(clk), .Q(ram[3270]) );
  DFF_X1 ram_reg_204__5_ ( .D(n10113), .CK(clk), .Q(ram[3269]) );
  DFF_X1 ram_reg_204__4_ ( .D(n10112), .CK(clk), .Q(ram[3268]) );
  DFF_X1 ram_reg_204__3_ ( .D(n10111), .CK(clk), .Q(ram[3267]) );
  DFF_X1 ram_reg_204__2_ ( .D(n10110), .CK(clk), .Q(ram[3266]) );
  DFF_X1 ram_reg_204__1_ ( .D(n10109), .CK(clk), .Q(ram[3265]) );
  DFF_X1 ram_reg_204__0_ ( .D(n10108), .CK(clk), .Q(ram[3264]) );
  DFF_X1 ram_reg_203__15_ ( .D(n10140), .CK(clk), .Q(ram[3263]) );
  DFF_X1 ram_reg_203__14_ ( .D(n10139), .CK(clk), .Q(ram[3262]) );
  DFF_X1 ram_reg_203__13_ ( .D(n10138), .CK(clk), .Q(ram[3261]) );
  DFF_X1 ram_reg_203__12_ ( .D(n10137), .CK(clk), .Q(ram[3260]) );
  DFF_X1 ram_reg_203__11_ ( .D(n10136), .CK(clk), .Q(ram[3259]) );
  DFF_X1 ram_reg_203__10_ ( .D(n10135), .CK(clk), .Q(ram[3258]) );
  DFF_X1 ram_reg_203__9_ ( .D(n10134), .CK(clk), .Q(ram[3257]) );
  DFF_X1 ram_reg_203__8_ ( .D(n10133), .CK(clk), .Q(ram[3256]) );
  DFF_X1 ram_reg_203__7_ ( .D(n10132), .CK(clk), .Q(ram[3255]) );
  DFF_X1 ram_reg_203__6_ ( .D(n10131), .CK(clk), .Q(ram[3254]) );
  DFF_X1 ram_reg_203__5_ ( .D(n10130), .CK(clk), .Q(ram[3253]) );
  DFF_X1 ram_reg_203__4_ ( .D(n10129), .CK(clk), .Q(ram[3252]) );
  DFF_X1 ram_reg_203__3_ ( .D(n10128), .CK(clk), .Q(ram[3251]) );
  DFF_X1 ram_reg_203__2_ ( .D(n10127), .CK(clk), .Q(ram[3250]) );
  DFF_X1 ram_reg_203__1_ ( .D(n10126), .CK(clk), .Q(ram[3249]) );
  DFF_X1 ram_reg_203__0_ ( .D(n10125), .CK(clk), .Q(ram[3248]) );
  DFF_X1 ram_reg_202__15_ ( .D(n10157), .CK(clk), .Q(ram[3247]) );
  DFF_X1 ram_reg_202__14_ ( .D(n10156), .CK(clk), .Q(ram[3246]) );
  DFF_X1 ram_reg_202__13_ ( .D(n10155), .CK(clk), .Q(ram[3245]) );
  DFF_X1 ram_reg_202__12_ ( .D(n10154), .CK(clk), .Q(ram[3244]) );
  DFF_X1 ram_reg_202__11_ ( .D(n10153), .CK(clk), .Q(ram[3243]) );
  DFF_X1 ram_reg_202__10_ ( .D(n10152), .CK(clk), .Q(ram[3242]) );
  DFF_X1 ram_reg_202__9_ ( .D(n10151), .CK(clk), .Q(ram[3241]) );
  DFF_X1 ram_reg_202__8_ ( .D(n10150), .CK(clk), .Q(ram[3240]) );
  DFF_X1 ram_reg_202__7_ ( .D(n10149), .CK(clk), .Q(ram[3239]) );
  DFF_X1 ram_reg_202__6_ ( .D(n10148), .CK(clk), .Q(ram[3238]) );
  DFF_X1 ram_reg_202__5_ ( .D(n10147), .CK(clk), .Q(ram[3237]) );
  DFF_X1 ram_reg_202__4_ ( .D(n10146), .CK(clk), .Q(ram[3236]) );
  DFF_X1 ram_reg_202__3_ ( .D(n10145), .CK(clk), .Q(ram[3235]) );
  DFF_X1 ram_reg_202__2_ ( .D(n10144), .CK(clk), .Q(ram[3234]) );
  DFF_X1 ram_reg_202__1_ ( .D(n10143), .CK(clk), .Q(ram[3233]) );
  DFF_X1 ram_reg_202__0_ ( .D(n10142), .CK(clk), .Q(ram[3232]) );
  DFF_X1 ram_reg_201__15_ ( .D(n10174), .CK(clk), .Q(ram[3231]) );
  DFF_X1 ram_reg_201__14_ ( .D(n10173), .CK(clk), .Q(ram[3230]) );
  DFF_X1 ram_reg_201__13_ ( .D(n10172), .CK(clk), .Q(ram[3229]) );
  DFF_X1 ram_reg_201__12_ ( .D(n10171), .CK(clk), .Q(ram[3228]) );
  DFF_X1 ram_reg_201__11_ ( .D(n10170), .CK(clk), .Q(ram[3227]) );
  DFF_X1 ram_reg_201__10_ ( .D(n10169), .CK(clk), .Q(ram[3226]) );
  DFF_X1 ram_reg_201__9_ ( .D(n10168), .CK(clk), .Q(ram[3225]) );
  DFF_X1 ram_reg_201__8_ ( .D(n10167), .CK(clk), .Q(ram[3224]) );
  DFF_X1 ram_reg_201__7_ ( .D(n10166), .CK(clk), .Q(ram[3223]) );
  DFF_X1 ram_reg_201__6_ ( .D(n10165), .CK(clk), .Q(ram[3222]) );
  DFF_X1 ram_reg_201__5_ ( .D(n10164), .CK(clk), .Q(ram[3221]) );
  DFF_X1 ram_reg_201__4_ ( .D(n10163), .CK(clk), .Q(ram[3220]) );
  DFF_X1 ram_reg_201__3_ ( .D(n10162), .CK(clk), .Q(ram[3219]) );
  DFF_X1 ram_reg_201__2_ ( .D(n10161), .CK(clk), .Q(ram[3218]) );
  DFF_X1 ram_reg_201__1_ ( .D(n10160), .CK(clk), .Q(ram[3217]) );
  DFF_X1 ram_reg_201__0_ ( .D(n10159), .CK(clk), .Q(ram[3216]) );
  DFF_X1 ram_reg_200__15_ ( .D(n10191), .CK(clk), .Q(ram[3215]) );
  DFF_X1 ram_reg_200__14_ ( .D(n10190), .CK(clk), .Q(ram[3214]) );
  DFF_X1 ram_reg_200__13_ ( .D(n10189), .CK(clk), .Q(ram[3213]) );
  DFF_X1 ram_reg_200__12_ ( .D(n10188), .CK(clk), .Q(ram[3212]) );
  DFF_X1 ram_reg_200__11_ ( .D(n10187), .CK(clk), .Q(ram[3211]) );
  DFF_X1 ram_reg_200__10_ ( .D(n10186), .CK(clk), .Q(ram[3210]) );
  DFF_X1 ram_reg_200__9_ ( .D(n10185), .CK(clk), .Q(ram[3209]) );
  DFF_X1 ram_reg_200__8_ ( .D(n10184), .CK(clk), .Q(ram[3208]) );
  DFF_X1 ram_reg_200__7_ ( .D(n10183), .CK(clk), .Q(ram[3207]) );
  DFF_X1 ram_reg_200__6_ ( .D(n10182), .CK(clk), .Q(ram[3206]) );
  DFF_X1 ram_reg_200__5_ ( .D(n10181), .CK(clk), .Q(ram[3205]) );
  DFF_X1 ram_reg_200__4_ ( .D(n10180), .CK(clk), .Q(ram[3204]) );
  DFF_X1 ram_reg_200__3_ ( .D(n10179), .CK(clk), .Q(ram[3203]) );
  DFF_X1 ram_reg_200__2_ ( .D(n10178), .CK(clk), .Q(ram[3202]) );
  DFF_X1 ram_reg_200__1_ ( .D(n10177), .CK(clk), .Q(ram[3201]) );
  DFF_X1 ram_reg_200__0_ ( .D(n10176), .CK(clk), .Q(ram[3200]) );
  DFF_X1 ram_reg_199__15_ ( .D(n10208), .CK(clk), .Q(ram[3199]) );
  DFF_X1 ram_reg_199__14_ ( .D(n10207), .CK(clk), .Q(ram[3198]) );
  DFF_X1 ram_reg_199__13_ ( .D(n10206), .CK(clk), .Q(ram[3197]) );
  DFF_X1 ram_reg_199__12_ ( .D(n10205), .CK(clk), .Q(ram[3196]) );
  DFF_X1 ram_reg_199__11_ ( .D(n10204), .CK(clk), .Q(ram[3195]) );
  DFF_X1 ram_reg_199__10_ ( .D(n10203), .CK(clk), .Q(ram[3194]) );
  DFF_X1 ram_reg_199__9_ ( .D(n10202), .CK(clk), .Q(ram[3193]) );
  DFF_X1 ram_reg_199__8_ ( .D(n10201), .CK(clk), .Q(ram[3192]) );
  DFF_X1 ram_reg_199__7_ ( .D(n10200), .CK(clk), .Q(ram[3191]) );
  DFF_X1 ram_reg_199__6_ ( .D(n10199), .CK(clk), .Q(ram[3190]) );
  DFF_X1 ram_reg_199__5_ ( .D(n10198), .CK(clk), .Q(ram[3189]) );
  DFF_X1 ram_reg_199__4_ ( .D(n10197), .CK(clk), .Q(ram[3188]) );
  DFF_X1 ram_reg_199__3_ ( .D(n10196), .CK(clk), .Q(ram[3187]) );
  DFF_X1 ram_reg_199__2_ ( .D(n10195), .CK(clk), .Q(ram[3186]) );
  DFF_X1 ram_reg_199__1_ ( .D(n10194), .CK(clk), .Q(ram[3185]) );
  DFF_X1 ram_reg_199__0_ ( .D(n10193), .CK(clk), .Q(ram[3184]) );
  DFF_X1 ram_reg_198__15_ ( .D(n10225), .CK(clk), .Q(ram[3183]) );
  DFF_X1 ram_reg_198__14_ ( .D(n10224), .CK(clk), .Q(ram[3182]) );
  DFF_X1 ram_reg_198__13_ ( .D(n10223), .CK(clk), .Q(ram[3181]) );
  DFF_X1 ram_reg_198__12_ ( .D(n10222), .CK(clk), .Q(ram[3180]) );
  DFF_X1 ram_reg_198__11_ ( .D(n10221), .CK(clk), .Q(ram[3179]) );
  DFF_X1 ram_reg_198__10_ ( .D(n10220), .CK(clk), .Q(ram[3178]) );
  DFF_X1 ram_reg_198__9_ ( .D(n10219), .CK(clk), .Q(ram[3177]) );
  DFF_X1 ram_reg_198__8_ ( .D(n10218), .CK(clk), .Q(ram[3176]) );
  DFF_X1 ram_reg_198__7_ ( .D(n10217), .CK(clk), .Q(ram[3175]) );
  DFF_X1 ram_reg_198__6_ ( .D(n10216), .CK(clk), .Q(ram[3174]) );
  DFF_X1 ram_reg_198__5_ ( .D(n10215), .CK(clk), .Q(ram[3173]) );
  DFF_X1 ram_reg_198__4_ ( .D(n10214), .CK(clk), .Q(ram[3172]) );
  DFF_X1 ram_reg_198__3_ ( .D(n10213), .CK(clk), .Q(ram[3171]) );
  DFF_X1 ram_reg_198__2_ ( .D(n10212), .CK(clk), .Q(ram[3170]) );
  DFF_X1 ram_reg_198__1_ ( .D(n10211), .CK(clk), .Q(ram[3169]) );
  DFF_X1 ram_reg_198__0_ ( .D(n10210), .CK(clk), .Q(ram[3168]) );
  DFF_X1 ram_reg_197__15_ ( .D(n10242), .CK(clk), .Q(ram[3167]) );
  DFF_X1 ram_reg_197__14_ ( .D(n10241), .CK(clk), .Q(ram[3166]) );
  DFF_X1 ram_reg_197__13_ ( .D(n10240), .CK(clk), .Q(ram[3165]) );
  DFF_X1 ram_reg_197__12_ ( .D(n10239), .CK(clk), .Q(ram[3164]) );
  DFF_X1 ram_reg_197__11_ ( .D(n10238), .CK(clk), .Q(ram[3163]) );
  DFF_X1 ram_reg_197__10_ ( .D(n10237), .CK(clk), .Q(ram[3162]) );
  DFF_X1 ram_reg_197__9_ ( .D(n10236), .CK(clk), .Q(ram[3161]) );
  DFF_X1 ram_reg_197__8_ ( .D(n10235), .CK(clk), .Q(ram[3160]) );
  DFF_X1 ram_reg_197__7_ ( .D(n10234), .CK(clk), .Q(ram[3159]) );
  DFF_X1 ram_reg_197__6_ ( .D(n10233), .CK(clk), .Q(ram[3158]) );
  DFF_X1 ram_reg_197__5_ ( .D(n10232), .CK(clk), .Q(ram[3157]) );
  DFF_X1 ram_reg_197__4_ ( .D(n10231), .CK(clk), .Q(ram[3156]) );
  DFF_X1 ram_reg_197__3_ ( .D(n10230), .CK(clk), .Q(ram[3155]) );
  DFF_X1 ram_reg_197__2_ ( .D(n10229), .CK(clk), .Q(ram[3154]) );
  DFF_X1 ram_reg_197__1_ ( .D(n10228), .CK(clk), .Q(ram[3153]) );
  DFF_X1 ram_reg_197__0_ ( .D(n10227), .CK(clk), .Q(ram[3152]) );
  DFF_X1 ram_reg_196__15_ ( .D(n10259), .CK(clk), .Q(ram[3151]) );
  DFF_X1 ram_reg_196__14_ ( .D(n10258), .CK(clk), .Q(ram[3150]) );
  DFF_X1 ram_reg_196__13_ ( .D(n10257), .CK(clk), .Q(ram[3149]) );
  DFF_X1 ram_reg_196__12_ ( .D(n10256), .CK(clk), .Q(ram[3148]) );
  DFF_X1 ram_reg_196__11_ ( .D(n10255), .CK(clk), .Q(ram[3147]) );
  DFF_X1 ram_reg_196__10_ ( .D(n10254), .CK(clk), .Q(ram[3146]) );
  DFF_X1 ram_reg_196__9_ ( .D(n10253), .CK(clk), .Q(ram[3145]) );
  DFF_X1 ram_reg_196__8_ ( .D(n10252), .CK(clk), .Q(ram[3144]) );
  DFF_X1 ram_reg_196__7_ ( .D(n10251), .CK(clk), .Q(ram[3143]) );
  DFF_X1 ram_reg_196__6_ ( .D(n10250), .CK(clk), .Q(ram[3142]) );
  DFF_X1 ram_reg_196__5_ ( .D(n10249), .CK(clk), .Q(ram[3141]) );
  DFF_X1 ram_reg_196__4_ ( .D(n10248), .CK(clk), .Q(ram[3140]) );
  DFF_X1 ram_reg_196__3_ ( .D(n10247), .CK(clk), .Q(ram[3139]) );
  DFF_X1 ram_reg_196__2_ ( .D(n10246), .CK(clk), .Q(ram[3138]) );
  DFF_X1 ram_reg_196__1_ ( .D(n10245), .CK(clk), .Q(ram[3137]) );
  DFF_X1 ram_reg_196__0_ ( .D(n10244), .CK(clk), .Q(ram[3136]) );
  DFF_X1 ram_reg_195__15_ ( .D(n10276), .CK(clk), .Q(ram[3135]) );
  DFF_X1 ram_reg_195__14_ ( .D(n10275), .CK(clk), .Q(ram[3134]) );
  DFF_X1 ram_reg_195__13_ ( .D(n10274), .CK(clk), .Q(ram[3133]) );
  DFF_X1 ram_reg_195__12_ ( .D(n10273), .CK(clk), .Q(ram[3132]) );
  DFF_X1 ram_reg_195__11_ ( .D(n10272), .CK(clk), .Q(ram[3131]) );
  DFF_X1 ram_reg_195__10_ ( .D(n10271), .CK(clk), .Q(ram[3130]) );
  DFF_X1 ram_reg_195__9_ ( .D(n10270), .CK(clk), .Q(ram[3129]) );
  DFF_X1 ram_reg_195__8_ ( .D(n10269), .CK(clk), .Q(ram[3128]) );
  DFF_X1 ram_reg_195__7_ ( .D(n10268), .CK(clk), .Q(ram[3127]) );
  DFF_X1 ram_reg_195__6_ ( .D(n10267), .CK(clk), .Q(ram[3126]) );
  DFF_X1 ram_reg_195__5_ ( .D(n10266), .CK(clk), .Q(ram[3125]) );
  DFF_X1 ram_reg_195__4_ ( .D(n10265), .CK(clk), .Q(ram[3124]) );
  DFF_X1 ram_reg_195__3_ ( .D(n10264), .CK(clk), .Q(ram[3123]) );
  DFF_X1 ram_reg_195__2_ ( .D(n10263), .CK(clk), .Q(ram[3122]) );
  DFF_X1 ram_reg_195__1_ ( .D(n10262), .CK(clk), .Q(ram[3121]) );
  DFF_X1 ram_reg_195__0_ ( .D(n10261), .CK(clk), .Q(ram[3120]) );
  DFF_X1 ram_reg_194__15_ ( .D(n10293), .CK(clk), .Q(ram[3119]) );
  DFF_X1 ram_reg_194__14_ ( .D(n10292), .CK(clk), .Q(ram[3118]) );
  DFF_X1 ram_reg_194__13_ ( .D(n10291), .CK(clk), .Q(ram[3117]) );
  DFF_X1 ram_reg_194__12_ ( .D(n10290), .CK(clk), .Q(ram[3116]) );
  DFF_X1 ram_reg_194__11_ ( .D(n10289), .CK(clk), .Q(ram[3115]) );
  DFF_X1 ram_reg_194__10_ ( .D(n10288), .CK(clk), .Q(ram[3114]) );
  DFF_X1 ram_reg_194__9_ ( .D(n10287), .CK(clk), .Q(ram[3113]) );
  DFF_X1 ram_reg_194__8_ ( .D(n10286), .CK(clk), .Q(ram[3112]) );
  DFF_X1 ram_reg_194__7_ ( .D(n10285), .CK(clk), .Q(ram[3111]) );
  DFF_X1 ram_reg_194__6_ ( .D(n10284), .CK(clk), .Q(ram[3110]) );
  DFF_X1 ram_reg_194__5_ ( .D(n10283), .CK(clk), .Q(ram[3109]) );
  DFF_X1 ram_reg_194__4_ ( .D(n10282), .CK(clk), .Q(ram[3108]) );
  DFF_X1 ram_reg_194__3_ ( .D(n10281), .CK(clk), .Q(ram[3107]) );
  DFF_X1 ram_reg_194__2_ ( .D(n10280), .CK(clk), .Q(ram[3106]) );
  DFF_X1 ram_reg_194__1_ ( .D(n10279), .CK(clk), .Q(ram[3105]) );
  DFF_X1 ram_reg_194__0_ ( .D(n10278), .CK(clk), .Q(ram[3104]) );
  DFF_X1 ram_reg_193__15_ ( .D(n10310), .CK(clk), .Q(ram[3103]) );
  DFF_X1 ram_reg_193__14_ ( .D(n10309), .CK(clk), .Q(ram[3102]) );
  DFF_X1 ram_reg_193__13_ ( .D(n10308), .CK(clk), .Q(ram[3101]) );
  DFF_X1 ram_reg_193__12_ ( .D(n10307), .CK(clk), .Q(ram[3100]) );
  DFF_X1 ram_reg_193__11_ ( .D(n10306), .CK(clk), .Q(ram[3099]) );
  DFF_X1 ram_reg_193__10_ ( .D(n10305), .CK(clk), .Q(ram[3098]) );
  DFF_X1 ram_reg_193__9_ ( .D(n10304), .CK(clk), .Q(ram[3097]) );
  DFF_X1 ram_reg_193__8_ ( .D(n10303), .CK(clk), .Q(ram[3096]) );
  DFF_X1 ram_reg_193__7_ ( .D(n10302), .CK(clk), .Q(ram[3095]) );
  DFF_X1 ram_reg_193__6_ ( .D(n10301), .CK(clk), .Q(ram[3094]) );
  DFF_X1 ram_reg_193__5_ ( .D(n10300), .CK(clk), .Q(ram[3093]) );
  DFF_X1 ram_reg_193__4_ ( .D(n10299), .CK(clk), .Q(ram[3092]) );
  DFF_X1 ram_reg_193__3_ ( .D(n10298), .CK(clk), .Q(ram[3091]) );
  DFF_X1 ram_reg_193__2_ ( .D(n10297), .CK(clk), .Q(ram[3090]) );
  DFF_X1 ram_reg_193__1_ ( .D(n10296), .CK(clk), .Q(ram[3089]) );
  DFF_X1 ram_reg_193__0_ ( .D(n10295), .CK(clk), .Q(ram[3088]) );
  DFF_X1 ram_reg_192__15_ ( .D(n10327), .CK(clk), .Q(ram[3087]) );
  DFF_X1 ram_reg_192__14_ ( .D(n10326), .CK(clk), .Q(ram[3086]) );
  DFF_X1 ram_reg_192__13_ ( .D(n10325), .CK(clk), .Q(ram[3085]) );
  DFF_X1 ram_reg_192__12_ ( .D(n10324), .CK(clk), .Q(ram[3084]) );
  DFF_X1 ram_reg_192__11_ ( .D(n10323), .CK(clk), .Q(ram[3083]) );
  DFF_X1 ram_reg_192__10_ ( .D(n10322), .CK(clk), .Q(ram[3082]) );
  DFF_X1 ram_reg_192__9_ ( .D(n10321), .CK(clk), .Q(ram[3081]) );
  DFF_X1 ram_reg_192__8_ ( .D(n10320), .CK(clk), .Q(ram[3080]) );
  DFF_X1 ram_reg_192__7_ ( .D(n10319), .CK(clk), .Q(ram[3079]) );
  DFF_X1 ram_reg_192__6_ ( .D(n10318), .CK(clk), .Q(ram[3078]) );
  DFF_X1 ram_reg_192__5_ ( .D(n10317), .CK(clk), .Q(ram[3077]) );
  DFF_X1 ram_reg_192__4_ ( .D(n10316), .CK(clk), .Q(ram[3076]) );
  DFF_X1 ram_reg_192__3_ ( .D(n10315), .CK(clk), .Q(ram[3075]) );
  DFF_X1 ram_reg_192__2_ ( .D(n10314), .CK(clk), .Q(ram[3074]) );
  DFF_X1 ram_reg_192__1_ ( .D(n10313), .CK(clk), .Q(ram[3073]) );
  DFF_X1 ram_reg_192__0_ ( .D(n10312), .CK(clk), .Q(ram[3072]) );
  DFF_X1 ram_reg_191__15_ ( .D(n10344), .CK(clk), .Q(ram[3071]) );
  DFF_X1 ram_reg_191__14_ ( .D(n10343), .CK(clk), .Q(ram[3070]) );
  DFF_X1 ram_reg_191__13_ ( .D(n10342), .CK(clk), .Q(ram[3069]) );
  DFF_X1 ram_reg_191__12_ ( .D(n10341), .CK(clk), .Q(ram[3068]) );
  DFF_X1 ram_reg_191__11_ ( .D(n10340), .CK(clk), .Q(ram[3067]) );
  DFF_X1 ram_reg_191__10_ ( .D(n10339), .CK(clk), .Q(ram[3066]) );
  DFF_X1 ram_reg_191__9_ ( .D(n10338), .CK(clk), .Q(ram[3065]) );
  DFF_X1 ram_reg_191__8_ ( .D(n10337), .CK(clk), .Q(ram[3064]) );
  DFF_X1 ram_reg_191__7_ ( .D(n10336), .CK(clk), .Q(ram[3063]) );
  DFF_X1 ram_reg_191__6_ ( .D(n10335), .CK(clk), .Q(ram[3062]) );
  DFF_X1 ram_reg_191__5_ ( .D(n10334), .CK(clk), .Q(ram[3061]) );
  DFF_X1 ram_reg_191__4_ ( .D(n10333), .CK(clk), .Q(ram[3060]) );
  DFF_X1 ram_reg_191__3_ ( .D(n10332), .CK(clk), .Q(ram[3059]) );
  DFF_X1 ram_reg_191__2_ ( .D(n10331), .CK(clk), .Q(ram[3058]) );
  DFF_X1 ram_reg_191__1_ ( .D(n10330), .CK(clk), .Q(ram[3057]) );
  DFF_X1 ram_reg_191__0_ ( .D(n10329), .CK(clk), .Q(ram[3056]) );
  DFF_X1 ram_reg_190__15_ ( .D(n10361), .CK(clk), .Q(ram[3055]) );
  DFF_X1 ram_reg_190__14_ ( .D(n10360), .CK(clk), .Q(ram[3054]) );
  DFF_X1 ram_reg_190__13_ ( .D(n10359), .CK(clk), .Q(ram[3053]) );
  DFF_X1 ram_reg_190__12_ ( .D(n10358), .CK(clk), .Q(ram[3052]) );
  DFF_X1 ram_reg_190__11_ ( .D(n10357), .CK(clk), .Q(ram[3051]) );
  DFF_X1 ram_reg_190__10_ ( .D(n10356), .CK(clk), .Q(ram[3050]) );
  DFF_X1 ram_reg_190__9_ ( .D(n10355), .CK(clk), .Q(ram[3049]) );
  DFF_X1 ram_reg_190__8_ ( .D(n10354), .CK(clk), .Q(ram[3048]) );
  DFF_X1 ram_reg_190__7_ ( .D(n10353), .CK(clk), .Q(ram[3047]) );
  DFF_X1 ram_reg_190__6_ ( .D(n10352), .CK(clk), .Q(ram[3046]) );
  DFF_X1 ram_reg_190__5_ ( .D(n10351), .CK(clk), .Q(ram[3045]) );
  DFF_X1 ram_reg_190__4_ ( .D(n10350), .CK(clk), .Q(ram[3044]) );
  DFF_X1 ram_reg_190__3_ ( .D(n10349), .CK(clk), .Q(ram[3043]) );
  DFF_X1 ram_reg_190__2_ ( .D(n10348), .CK(clk), .Q(ram[3042]) );
  DFF_X1 ram_reg_190__1_ ( .D(n10347), .CK(clk), .Q(ram[3041]) );
  DFF_X1 ram_reg_190__0_ ( .D(n10346), .CK(clk), .Q(ram[3040]) );
  DFF_X1 ram_reg_189__15_ ( .D(n10378), .CK(clk), .Q(ram[3039]) );
  DFF_X1 ram_reg_189__14_ ( .D(n10377), .CK(clk), .Q(ram[3038]) );
  DFF_X1 ram_reg_189__13_ ( .D(n10376), .CK(clk), .Q(ram[3037]) );
  DFF_X1 ram_reg_189__12_ ( .D(n10375), .CK(clk), .Q(ram[3036]) );
  DFF_X1 ram_reg_189__11_ ( .D(n10374), .CK(clk), .Q(ram[3035]) );
  DFF_X1 ram_reg_189__10_ ( .D(n10373), .CK(clk), .Q(ram[3034]) );
  DFF_X1 ram_reg_189__9_ ( .D(n10372), .CK(clk), .Q(ram[3033]) );
  DFF_X1 ram_reg_189__8_ ( .D(n10371), .CK(clk), .Q(ram[3032]) );
  DFF_X1 ram_reg_189__7_ ( .D(n10370), .CK(clk), .Q(ram[3031]) );
  DFF_X1 ram_reg_189__6_ ( .D(n10369), .CK(clk), .Q(ram[3030]) );
  DFF_X1 ram_reg_189__5_ ( .D(n10368), .CK(clk), .Q(ram[3029]) );
  DFF_X1 ram_reg_189__4_ ( .D(n10367), .CK(clk), .Q(ram[3028]) );
  DFF_X1 ram_reg_189__3_ ( .D(n10366), .CK(clk), .Q(ram[3027]) );
  DFF_X1 ram_reg_189__2_ ( .D(n10365), .CK(clk), .Q(ram[3026]) );
  DFF_X1 ram_reg_189__1_ ( .D(n10364), .CK(clk), .Q(ram[3025]) );
  DFF_X1 ram_reg_189__0_ ( .D(n10363), .CK(clk), .Q(ram[3024]) );
  DFF_X1 ram_reg_188__15_ ( .D(n10395), .CK(clk), .Q(ram[3023]) );
  DFF_X1 ram_reg_188__14_ ( .D(n10394), .CK(clk), .Q(ram[3022]) );
  DFF_X1 ram_reg_188__13_ ( .D(n10393), .CK(clk), .Q(ram[3021]) );
  DFF_X1 ram_reg_188__12_ ( .D(n10392), .CK(clk), .Q(ram[3020]) );
  DFF_X1 ram_reg_188__11_ ( .D(n10391), .CK(clk), .Q(ram[3019]) );
  DFF_X1 ram_reg_188__10_ ( .D(n10390), .CK(clk), .Q(ram[3018]) );
  DFF_X1 ram_reg_188__9_ ( .D(n10389), .CK(clk), .Q(ram[3017]) );
  DFF_X1 ram_reg_188__8_ ( .D(n10388), .CK(clk), .Q(ram[3016]) );
  DFF_X1 ram_reg_188__7_ ( .D(n10387), .CK(clk), .Q(ram[3015]) );
  DFF_X1 ram_reg_188__6_ ( .D(n10386), .CK(clk), .Q(ram[3014]) );
  DFF_X1 ram_reg_188__5_ ( .D(n10385), .CK(clk), .Q(ram[3013]) );
  DFF_X1 ram_reg_188__4_ ( .D(n10384), .CK(clk), .Q(ram[3012]) );
  DFF_X1 ram_reg_188__3_ ( .D(n10383), .CK(clk), .Q(ram[3011]) );
  DFF_X1 ram_reg_188__2_ ( .D(n10382), .CK(clk), .Q(ram[3010]) );
  DFF_X1 ram_reg_188__1_ ( .D(n10381), .CK(clk), .Q(ram[3009]) );
  DFF_X1 ram_reg_188__0_ ( .D(n10380), .CK(clk), .Q(ram[3008]) );
  DFF_X1 ram_reg_187__15_ ( .D(n10412), .CK(clk), .Q(ram[3007]) );
  DFF_X1 ram_reg_187__14_ ( .D(n10411), .CK(clk), .Q(ram[3006]) );
  DFF_X1 ram_reg_187__13_ ( .D(n10410), .CK(clk), .Q(ram[3005]) );
  DFF_X1 ram_reg_187__12_ ( .D(n10409), .CK(clk), .Q(ram[3004]) );
  DFF_X1 ram_reg_187__11_ ( .D(n10408), .CK(clk), .Q(ram[3003]) );
  DFF_X1 ram_reg_187__10_ ( .D(n10407), .CK(clk), .Q(ram[3002]) );
  DFF_X1 ram_reg_187__9_ ( .D(n10406), .CK(clk), .Q(ram[3001]) );
  DFF_X1 ram_reg_187__8_ ( .D(n10405), .CK(clk), .Q(ram[3000]) );
  DFF_X1 ram_reg_187__7_ ( .D(n10404), .CK(clk), .Q(ram[2999]) );
  DFF_X1 ram_reg_187__6_ ( .D(n10403), .CK(clk), .Q(ram[2998]) );
  DFF_X1 ram_reg_187__5_ ( .D(n10402), .CK(clk), .Q(ram[2997]) );
  DFF_X1 ram_reg_187__4_ ( .D(n10401), .CK(clk), .Q(ram[2996]) );
  DFF_X1 ram_reg_187__3_ ( .D(n10400), .CK(clk), .Q(ram[2995]) );
  DFF_X1 ram_reg_187__2_ ( .D(n10399), .CK(clk), .Q(ram[2994]) );
  DFF_X1 ram_reg_187__1_ ( .D(n10398), .CK(clk), .Q(ram[2993]) );
  DFF_X1 ram_reg_187__0_ ( .D(n10397), .CK(clk), .Q(ram[2992]) );
  DFF_X1 ram_reg_186__15_ ( .D(n10429), .CK(clk), .Q(ram[2991]) );
  DFF_X1 ram_reg_186__14_ ( .D(n10428), .CK(clk), .Q(ram[2990]) );
  DFF_X1 ram_reg_186__13_ ( .D(n10427), .CK(clk), .Q(ram[2989]) );
  DFF_X1 ram_reg_186__12_ ( .D(n10426), .CK(clk), .Q(ram[2988]) );
  DFF_X1 ram_reg_186__11_ ( .D(n10425), .CK(clk), .Q(ram[2987]) );
  DFF_X1 ram_reg_186__10_ ( .D(n10424), .CK(clk), .Q(ram[2986]) );
  DFF_X1 ram_reg_186__9_ ( .D(n10423), .CK(clk), .Q(ram[2985]) );
  DFF_X1 ram_reg_186__8_ ( .D(n10422), .CK(clk), .Q(ram[2984]) );
  DFF_X1 ram_reg_186__7_ ( .D(n10421), .CK(clk), .Q(ram[2983]) );
  DFF_X1 ram_reg_186__6_ ( .D(n10420), .CK(clk), .Q(ram[2982]) );
  DFF_X1 ram_reg_186__5_ ( .D(n10419), .CK(clk), .Q(ram[2981]) );
  DFF_X1 ram_reg_186__4_ ( .D(n10418), .CK(clk), .Q(ram[2980]) );
  DFF_X1 ram_reg_186__3_ ( .D(n10417), .CK(clk), .Q(ram[2979]) );
  DFF_X1 ram_reg_186__2_ ( .D(n10416), .CK(clk), .Q(ram[2978]) );
  DFF_X1 ram_reg_186__1_ ( .D(n10415), .CK(clk), .Q(ram[2977]) );
  DFF_X1 ram_reg_186__0_ ( .D(n10414), .CK(clk), .Q(ram[2976]) );
  DFF_X1 ram_reg_185__15_ ( .D(n10446), .CK(clk), .Q(ram[2975]) );
  DFF_X1 ram_reg_185__14_ ( .D(n10445), .CK(clk), .Q(ram[2974]) );
  DFF_X1 ram_reg_185__13_ ( .D(n10444), .CK(clk), .Q(ram[2973]) );
  DFF_X1 ram_reg_185__12_ ( .D(n10443), .CK(clk), .Q(ram[2972]) );
  DFF_X1 ram_reg_185__11_ ( .D(n10442), .CK(clk), .Q(ram[2971]) );
  DFF_X1 ram_reg_185__10_ ( .D(n10441), .CK(clk), .Q(ram[2970]) );
  DFF_X1 ram_reg_185__9_ ( .D(n10440), .CK(clk), .Q(ram[2969]) );
  DFF_X1 ram_reg_185__8_ ( .D(n10439), .CK(clk), .Q(ram[2968]) );
  DFF_X1 ram_reg_185__7_ ( .D(n10438), .CK(clk), .Q(ram[2967]) );
  DFF_X1 ram_reg_185__6_ ( .D(n10437), .CK(clk), .Q(ram[2966]) );
  DFF_X1 ram_reg_185__5_ ( .D(n10436), .CK(clk), .Q(ram[2965]) );
  DFF_X1 ram_reg_185__4_ ( .D(n10435), .CK(clk), .Q(ram[2964]) );
  DFF_X1 ram_reg_185__3_ ( .D(n10434), .CK(clk), .Q(ram[2963]) );
  DFF_X1 ram_reg_185__2_ ( .D(n10433), .CK(clk), .Q(ram[2962]) );
  DFF_X1 ram_reg_185__1_ ( .D(n10432), .CK(clk), .Q(ram[2961]) );
  DFF_X1 ram_reg_185__0_ ( .D(n10431), .CK(clk), .Q(ram[2960]) );
  DFF_X1 ram_reg_184__15_ ( .D(n10463), .CK(clk), .Q(ram[2959]) );
  DFF_X1 ram_reg_184__14_ ( .D(n10462), .CK(clk), .Q(ram[2958]) );
  DFF_X1 ram_reg_184__13_ ( .D(n10461), .CK(clk), .Q(ram[2957]) );
  DFF_X1 ram_reg_184__12_ ( .D(n10460), .CK(clk), .Q(ram[2956]) );
  DFF_X1 ram_reg_184__11_ ( .D(n10459), .CK(clk), .Q(ram[2955]) );
  DFF_X1 ram_reg_184__10_ ( .D(n10458), .CK(clk), .Q(ram[2954]) );
  DFF_X1 ram_reg_184__9_ ( .D(n10457), .CK(clk), .Q(ram[2953]) );
  DFF_X1 ram_reg_184__8_ ( .D(n10456), .CK(clk), .Q(ram[2952]) );
  DFF_X1 ram_reg_184__7_ ( .D(n10455), .CK(clk), .Q(ram[2951]) );
  DFF_X1 ram_reg_184__6_ ( .D(n10454), .CK(clk), .Q(ram[2950]) );
  DFF_X1 ram_reg_184__5_ ( .D(n10453), .CK(clk), .Q(ram[2949]) );
  DFF_X1 ram_reg_184__4_ ( .D(n10452), .CK(clk), .Q(ram[2948]) );
  DFF_X1 ram_reg_184__3_ ( .D(n10451), .CK(clk), .Q(ram[2947]) );
  DFF_X1 ram_reg_184__2_ ( .D(n10450), .CK(clk), .Q(ram[2946]) );
  DFF_X1 ram_reg_184__1_ ( .D(n10449), .CK(clk), .Q(ram[2945]) );
  DFF_X1 ram_reg_184__0_ ( .D(n10448), .CK(clk), .Q(ram[2944]) );
  DFF_X1 ram_reg_183__15_ ( .D(n10480), .CK(clk), .Q(ram[2943]) );
  DFF_X1 ram_reg_183__14_ ( .D(n10479), .CK(clk), .Q(ram[2942]) );
  DFF_X1 ram_reg_183__13_ ( .D(n10478), .CK(clk), .Q(ram[2941]) );
  DFF_X1 ram_reg_183__12_ ( .D(n10477), .CK(clk), .Q(ram[2940]) );
  DFF_X1 ram_reg_183__11_ ( .D(n10476), .CK(clk), .Q(ram[2939]) );
  DFF_X1 ram_reg_183__10_ ( .D(n10475), .CK(clk), .Q(ram[2938]) );
  DFF_X1 ram_reg_183__9_ ( .D(n10474), .CK(clk), .Q(ram[2937]) );
  DFF_X1 ram_reg_183__8_ ( .D(n10473), .CK(clk), .Q(ram[2936]) );
  DFF_X1 ram_reg_183__7_ ( .D(n10472), .CK(clk), .Q(ram[2935]) );
  DFF_X1 ram_reg_183__6_ ( .D(n10471), .CK(clk), .Q(ram[2934]) );
  DFF_X1 ram_reg_183__5_ ( .D(n10470), .CK(clk), .Q(ram[2933]) );
  DFF_X1 ram_reg_183__4_ ( .D(n10469), .CK(clk), .Q(ram[2932]) );
  DFF_X1 ram_reg_183__3_ ( .D(n10468), .CK(clk), .Q(ram[2931]) );
  DFF_X1 ram_reg_183__2_ ( .D(n10467), .CK(clk), .Q(ram[2930]) );
  DFF_X1 ram_reg_183__1_ ( .D(n10466), .CK(clk), .Q(ram[2929]) );
  DFF_X1 ram_reg_183__0_ ( .D(n10465), .CK(clk), .Q(ram[2928]) );
  DFF_X1 ram_reg_182__15_ ( .D(n10497), .CK(clk), .Q(ram[2927]) );
  DFF_X1 ram_reg_182__14_ ( .D(n10496), .CK(clk), .Q(ram[2926]) );
  DFF_X1 ram_reg_182__13_ ( .D(n10495), .CK(clk), .Q(ram[2925]) );
  DFF_X1 ram_reg_182__12_ ( .D(n10494), .CK(clk), .Q(ram[2924]) );
  DFF_X1 ram_reg_182__11_ ( .D(n10493), .CK(clk), .Q(ram[2923]) );
  DFF_X1 ram_reg_182__10_ ( .D(n10492), .CK(clk), .Q(ram[2922]) );
  DFF_X1 ram_reg_182__9_ ( .D(n10491), .CK(clk), .Q(ram[2921]) );
  DFF_X1 ram_reg_182__8_ ( .D(n10490), .CK(clk), .Q(ram[2920]) );
  DFF_X1 ram_reg_182__7_ ( .D(n10489), .CK(clk), .Q(ram[2919]) );
  DFF_X1 ram_reg_182__6_ ( .D(n10488), .CK(clk), .Q(ram[2918]) );
  DFF_X1 ram_reg_182__5_ ( .D(n10487), .CK(clk), .Q(ram[2917]) );
  DFF_X1 ram_reg_182__4_ ( .D(n10486), .CK(clk), .Q(ram[2916]) );
  DFF_X1 ram_reg_182__3_ ( .D(n10485), .CK(clk), .Q(ram[2915]) );
  DFF_X1 ram_reg_182__2_ ( .D(n10484), .CK(clk), .Q(ram[2914]) );
  DFF_X1 ram_reg_182__1_ ( .D(n10483), .CK(clk), .Q(ram[2913]) );
  DFF_X1 ram_reg_182__0_ ( .D(n10482), .CK(clk), .Q(ram[2912]) );
  DFF_X1 ram_reg_181__15_ ( .D(n10514), .CK(clk), .Q(ram[2911]) );
  DFF_X1 ram_reg_181__14_ ( .D(n10513), .CK(clk), .Q(ram[2910]) );
  DFF_X1 ram_reg_181__13_ ( .D(n10512), .CK(clk), .Q(ram[2909]) );
  DFF_X1 ram_reg_181__12_ ( .D(n10511), .CK(clk), .Q(ram[2908]) );
  DFF_X1 ram_reg_181__11_ ( .D(n10510), .CK(clk), .Q(ram[2907]) );
  DFF_X1 ram_reg_181__10_ ( .D(n10509), .CK(clk), .Q(ram[2906]) );
  DFF_X1 ram_reg_181__9_ ( .D(n10508), .CK(clk), .Q(ram[2905]) );
  DFF_X1 ram_reg_181__8_ ( .D(n10507), .CK(clk), .Q(ram[2904]) );
  DFF_X1 ram_reg_181__7_ ( .D(n10506), .CK(clk), .Q(ram[2903]) );
  DFF_X1 ram_reg_181__6_ ( .D(n10505), .CK(clk), .Q(ram[2902]) );
  DFF_X1 ram_reg_181__5_ ( .D(n10504), .CK(clk), .Q(ram[2901]) );
  DFF_X1 ram_reg_181__4_ ( .D(n10503), .CK(clk), .Q(ram[2900]) );
  DFF_X1 ram_reg_181__3_ ( .D(n10502), .CK(clk), .Q(ram[2899]) );
  DFF_X1 ram_reg_181__2_ ( .D(n10501), .CK(clk), .Q(ram[2898]) );
  DFF_X1 ram_reg_181__1_ ( .D(n10500), .CK(clk), .Q(ram[2897]) );
  DFF_X1 ram_reg_181__0_ ( .D(n10499), .CK(clk), .Q(ram[2896]) );
  DFF_X1 ram_reg_180__15_ ( .D(n10531), .CK(clk), .Q(ram[2895]) );
  DFF_X1 ram_reg_180__14_ ( .D(n10530), .CK(clk), .Q(ram[2894]) );
  DFF_X1 ram_reg_180__13_ ( .D(n10529), .CK(clk), .Q(ram[2893]) );
  DFF_X1 ram_reg_180__12_ ( .D(n10528), .CK(clk), .Q(ram[2892]) );
  DFF_X1 ram_reg_180__11_ ( .D(n10527), .CK(clk), .Q(ram[2891]) );
  DFF_X1 ram_reg_180__10_ ( .D(n10526), .CK(clk), .Q(ram[2890]) );
  DFF_X1 ram_reg_180__9_ ( .D(n10525), .CK(clk), .Q(ram[2889]) );
  DFF_X1 ram_reg_180__8_ ( .D(n10524), .CK(clk), .Q(ram[2888]) );
  DFF_X1 ram_reg_180__7_ ( .D(n10523), .CK(clk), .Q(ram[2887]) );
  DFF_X1 ram_reg_180__6_ ( .D(n10522), .CK(clk), .Q(ram[2886]) );
  DFF_X1 ram_reg_180__5_ ( .D(n10521), .CK(clk), .Q(ram[2885]) );
  DFF_X1 ram_reg_180__4_ ( .D(n10520), .CK(clk), .Q(ram[2884]) );
  DFF_X1 ram_reg_180__3_ ( .D(n10519), .CK(clk), .Q(ram[2883]) );
  DFF_X1 ram_reg_180__2_ ( .D(n10518), .CK(clk), .Q(ram[2882]) );
  DFF_X1 ram_reg_180__1_ ( .D(n10517), .CK(clk), .Q(ram[2881]) );
  DFF_X1 ram_reg_180__0_ ( .D(n10516), .CK(clk), .Q(ram[2880]) );
  DFF_X1 ram_reg_179__15_ ( .D(n10548), .CK(clk), .Q(ram[2879]) );
  DFF_X1 ram_reg_179__14_ ( .D(n10547), .CK(clk), .Q(ram[2878]) );
  DFF_X1 ram_reg_179__13_ ( .D(n10546), .CK(clk), .Q(ram[2877]) );
  DFF_X1 ram_reg_179__12_ ( .D(n10545), .CK(clk), .Q(ram[2876]) );
  DFF_X1 ram_reg_179__11_ ( .D(n10544), .CK(clk), .Q(ram[2875]) );
  DFF_X1 ram_reg_179__10_ ( .D(n10543), .CK(clk), .Q(ram[2874]) );
  DFF_X1 ram_reg_179__9_ ( .D(n10542), .CK(clk), .Q(ram[2873]) );
  DFF_X1 ram_reg_179__8_ ( .D(n10541), .CK(clk), .Q(ram[2872]) );
  DFF_X1 ram_reg_179__7_ ( .D(n10540), .CK(clk), .Q(ram[2871]) );
  DFF_X1 ram_reg_179__6_ ( .D(n10539), .CK(clk), .Q(ram[2870]) );
  DFF_X1 ram_reg_179__5_ ( .D(n10538), .CK(clk), .Q(ram[2869]) );
  DFF_X1 ram_reg_179__4_ ( .D(n10537), .CK(clk), .Q(ram[2868]) );
  DFF_X1 ram_reg_179__3_ ( .D(n10536), .CK(clk), .Q(ram[2867]) );
  DFF_X1 ram_reg_179__2_ ( .D(n10535), .CK(clk), .Q(ram[2866]) );
  DFF_X1 ram_reg_179__1_ ( .D(n10534), .CK(clk), .Q(ram[2865]) );
  DFF_X1 ram_reg_179__0_ ( .D(n10533), .CK(clk), .Q(ram[2864]) );
  DFF_X1 ram_reg_178__15_ ( .D(n10565), .CK(clk), .Q(ram[2863]) );
  DFF_X1 ram_reg_178__14_ ( .D(n10564), .CK(clk), .Q(ram[2862]) );
  DFF_X1 ram_reg_178__13_ ( .D(n10563), .CK(clk), .Q(ram[2861]) );
  DFF_X1 ram_reg_178__12_ ( .D(n10562), .CK(clk), .Q(ram[2860]) );
  DFF_X1 ram_reg_178__11_ ( .D(n10561), .CK(clk), .Q(ram[2859]) );
  DFF_X1 ram_reg_178__10_ ( .D(n10560), .CK(clk), .Q(ram[2858]) );
  DFF_X1 ram_reg_178__9_ ( .D(n10559), .CK(clk), .Q(ram[2857]) );
  DFF_X1 ram_reg_178__8_ ( .D(n10558), .CK(clk), .Q(ram[2856]) );
  DFF_X1 ram_reg_178__7_ ( .D(n10557), .CK(clk), .Q(ram[2855]) );
  DFF_X1 ram_reg_178__6_ ( .D(n10556), .CK(clk), .Q(ram[2854]) );
  DFF_X1 ram_reg_178__5_ ( .D(n10555), .CK(clk), .Q(ram[2853]) );
  DFF_X1 ram_reg_178__4_ ( .D(n10554), .CK(clk), .Q(ram[2852]) );
  DFF_X1 ram_reg_178__3_ ( .D(n10553), .CK(clk), .Q(ram[2851]) );
  DFF_X1 ram_reg_178__2_ ( .D(n10552), .CK(clk), .Q(ram[2850]) );
  DFF_X1 ram_reg_178__1_ ( .D(n10551), .CK(clk), .Q(ram[2849]) );
  DFF_X1 ram_reg_178__0_ ( .D(n10550), .CK(clk), .Q(ram[2848]) );
  DFF_X1 ram_reg_177__15_ ( .D(n10582), .CK(clk), .Q(ram[2847]) );
  DFF_X1 ram_reg_177__14_ ( .D(n10581), .CK(clk), .Q(ram[2846]) );
  DFF_X1 ram_reg_177__13_ ( .D(n10580), .CK(clk), .Q(ram[2845]) );
  DFF_X1 ram_reg_177__12_ ( .D(n10579), .CK(clk), .Q(ram[2844]) );
  DFF_X1 ram_reg_177__11_ ( .D(n10578), .CK(clk), .Q(ram[2843]) );
  DFF_X1 ram_reg_177__10_ ( .D(n10577), .CK(clk), .Q(ram[2842]) );
  DFF_X1 ram_reg_177__9_ ( .D(n10576), .CK(clk), .Q(ram[2841]) );
  DFF_X1 ram_reg_177__8_ ( .D(n10575), .CK(clk), .Q(ram[2840]) );
  DFF_X1 ram_reg_177__7_ ( .D(n10574), .CK(clk), .Q(ram[2839]) );
  DFF_X1 ram_reg_177__6_ ( .D(n10573), .CK(clk), .Q(ram[2838]) );
  DFF_X1 ram_reg_177__5_ ( .D(n10572), .CK(clk), .Q(ram[2837]) );
  DFF_X1 ram_reg_177__4_ ( .D(n10571), .CK(clk), .Q(ram[2836]) );
  DFF_X1 ram_reg_177__3_ ( .D(n10570), .CK(clk), .Q(ram[2835]) );
  DFF_X1 ram_reg_177__2_ ( .D(n10569), .CK(clk), .Q(ram[2834]) );
  DFF_X1 ram_reg_177__1_ ( .D(n10568), .CK(clk), .Q(ram[2833]) );
  DFF_X1 ram_reg_177__0_ ( .D(n10567), .CK(clk), .Q(ram[2832]) );
  DFF_X1 ram_reg_176__15_ ( .D(n10599), .CK(clk), .Q(ram[2831]) );
  DFF_X1 ram_reg_176__14_ ( .D(n10598), .CK(clk), .Q(ram[2830]) );
  DFF_X1 ram_reg_176__13_ ( .D(n10597), .CK(clk), .Q(ram[2829]) );
  DFF_X1 ram_reg_176__12_ ( .D(n10596), .CK(clk), .Q(ram[2828]) );
  DFF_X1 ram_reg_176__11_ ( .D(n10595), .CK(clk), .Q(ram[2827]) );
  DFF_X1 ram_reg_176__10_ ( .D(n10594), .CK(clk), .Q(ram[2826]) );
  DFF_X1 ram_reg_176__9_ ( .D(n10593), .CK(clk), .Q(ram[2825]) );
  DFF_X1 ram_reg_176__8_ ( .D(n10592), .CK(clk), .Q(ram[2824]) );
  DFF_X1 ram_reg_176__7_ ( .D(n10591), .CK(clk), .Q(ram[2823]) );
  DFF_X1 ram_reg_176__6_ ( .D(n10590), .CK(clk), .Q(ram[2822]) );
  DFF_X1 ram_reg_176__5_ ( .D(n10589), .CK(clk), .Q(ram[2821]) );
  DFF_X1 ram_reg_176__4_ ( .D(n10588), .CK(clk), .Q(ram[2820]) );
  DFF_X1 ram_reg_176__3_ ( .D(n10587), .CK(clk), .Q(ram[2819]) );
  DFF_X1 ram_reg_176__2_ ( .D(n10586), .CK(clk), .Q(ram[2818]) );
  DFF_X1 ram_reg_176__1_ ( .D(n10585), .CK(clk), .Q(ram[2817]) );
  DFF_X1 ram_reg_176__0_ ( .D(n10584), .CK(clk), .Q(ram[2816]) );
  DFF_X1 ram_reg_175__15_ ( .D(n10616), .CK(clk), .Q(ram[2815]) );
  DFF_X1 ram_reg_175__14_ ( .D(n10615), .CK(clk), .Q(ram[2814]) );
  DFF_X1 ram_reg_175__13_ ( .D(n10614), .CK(clk), .Q(ram[2813]) );
  DFF_X1 ram_reg_175__12_ ( .D(n10613), .CK(clk), .Q(ram[2812]) );
  DFF_X1 ram_reg_175__11_ ( .D(n10612), .CK(clk), .Q(ram[2811]) );
  DFF_X1 ram_reg_175__10_ ( .D(n10611), .CK(clk), .Q(ram[2810]) );
  DFF_X1 ram_reg_175__9_ ( .D(n10610), .CK(clk), .Q(ram[2809]) );
  DFF_X1 ram_reg_175__8_ ( .D(n10609), .CK(clk), .Q(ram[2808]) );
  DFF_X1 ram_reg_175__7_ ( .D(n10608), .CK(clk), .Q(ram[2807]) );
  DFF_X1 ram_reg_175__6_ ( .D(n10607), .CK(clk), .Q(ram[2806]) );
  DFF_X1 ram_reg_175__5_ ( .D(n10606), .CK(clk), .Q(ram[2805]) );
  DFF_X1 ram_reg_175__4_ ( .D(n10605), .CK(clk), .Q(ram[2804]) );
  DFF_X1 ram_reg_175__3_ ( .D(n10604), .CK(clk), .Q(ram[2803]) );
  DFF_X1 ram_reg_175__2_ ( .D(n10603), .CK(clk), .Q(ram[2802]) );
  DFF_X1 ram_reg_175__1_ ( .D(n10602), .CK(clk), .Q(ram[2801]) );
  DFF_X1 ram_reg_175__0_ ( .D(n10601), .CK(clk), .Q(ram[2800]) );
  DFF_X1 ram_reg_174__15_ ( .D(n10633), .CK(clk), .Q(ram[2799]) );
  DFF_X1 ram_reg_174__14_ ( .D(n10632), .CK(clk), .Q(ram[2798]) );
  DFF_X1 ram_reg_174__13_ ( .D(n10631), .CK(clk), .Q(ram[2797]) );
  DFF_X1 ram_reg_174__12_ ( .D(n10630), .CK(clk), .Q(ram[2796]) );
  DFF_X1 ram_reg_174__11_ ( .D(n10629), .CK(clk), .Q(ram[2795]) );
  DFF_X1 ram_reg_174__10_ ( .D(n10628), .CK(clk), .Q(ram[2794]) );
  DFF_X1 ram_reg_174__9_ ( .D(n10627), .CK(clk), .Q(ram[2793]) );
  DFF_X1 ram_reg_174__8_ ( .D(n10626), .CK(clk), .Q(ram[2792]) );
  DFF_X1 ram_reg_174__7_ ( .D(n10625), .CK(clk), .Q(ram[2791]) );
  DFF_X1 ram_reg_174__6_ ( .D(n10624), .CK(clk), .Q(ram[2790]) );
  DFF_X1 ram_reg_174__5_ ( .D(n10623), .CK(clk), .Q(ram[2789]) );
  DFF_X1 ram_reg_174__4_ ( .D(n10622), .CK(clk), .Q(ram[2788]) );
  DFF_X1 ram_reg_174__3_ ( .D(n10621), .CK(clk), .Q(ram[2787]) );
  DFF_X1 ram_reg_174__2_ ( .D(n10620), .CK(clk), .Q(ram[2786]) );
  DFF_X1 ram_reg_174__1_ ( .D(n10619), .CK(clk), .Q(ram[2785]) );
  DFF_X1 ram_reg_174__0_ ( .D(n10618), .CK(clk), .Q(ram[2784]) );
  DFF_X1 ram_reg_173__15_ ( .D(n10650), .CK(clk), .Q(ram[2783]) );
  DFF_X1 ram_reg_173__14_ ( .D(n10649), .CK(clk), .Q(ram[2782]) );
  DFF_X1 ram_reg_173__13_ ( .D(n10648), .CK(clk), .Q(ram[2781]) );
  DFF_X1 ram_reg_173__12_ ( .D(n10647), .CK(clk), .Q(ram[2780]) );
  DFF_X1 ram_reg_173__11_ ( .D(n10646), .CK(clk), .Q(ram[2779]) );
  DFF_X1 ram_reg_173__10_ ( .D(n10645), .CK(clk), .Q(ram[2778]) );
  DFF_X1 ram_reg_173__9_ ( .D(n10644), .CK(clk), .Q(ram[2777]) );
  DFF_X1 ram_reg_173__8_ ( .D(n10643), .CK(clk), .Q(ram[2776]) );
  DFF_X1 ram_reg_173__7_ ( .D(n10642), .CK(clk), .Q(ram[2775]) );
  DFF_X1 ram_reg_173__6_ ( .D(n10641), .CK(clk), .Q(ram[2774]) );
  DFF_X1 ram_reg_173__5_ ( .D(n10640), .CK(clk), .Q(ram[2773]) );
  DFF_X1 ram_reg_173__4_ ( .D(n10639), .CK(clk), .Q(ram[2772]) );
  DFF_X1 ram_reg_173__3_ ( .D(n10638), .CK(clk), .Q(ram[2771]) );
  DFF_X1 ram_reg_173__2_ ( .D(n10637), .CK(clk), .Q(ram[2770]) );
  DFF_X1 ram_reg_173__1_ ( .D(n10636), .CK(clk), .Q(ram[2769]) );
  DFF_X1 ram_reg_173__0_ ( .D(n10635), .CK(clk), .Q(ram[2768]) );
  DFF_X1 ram_reg_172__15_ ( .D(n10667), .CK(clk), .Q(ram[2767]) );
  DFF_X1 ram_reg_172__14_ ( .D(n10666), .CK(clk), .Q(ram[2766]) );
  DFF_X1 ram_reg_172__13_ ( .D(n10665), .CK(clk), .Q(ram[2765]) );
  DFF_X1 ram_reg_172__12_ ( .D(n10664), .CK(clk), .Q(ram[2764]) );
  DFF_X1 ram_reg_172__11_ ( .D(n10663), .CK(clk), .Q(ram[2763]) );
  DFF_X1 ram_reg_172__10_ ( .D(n10662), .CK(clk), .Q(ram[2762]) );
  DFF_X1 ram_reg_172__9_ ( .D(n10661), .CK(clk), .Q(ram[2761]) );
  DFF_X1 ram_reg_172__8_ ( .D(n10660), .CK(clk), .Q(ram[2760]) );
  DFF_X1 ram_reg_172__7_ ( .D(n10659), .CK(clk), .Q(ram[2759]) );
  DFF_X1 ram_reg_172__6_ ( .D(n10658), .CK(clk), .Q(ram[2758]) );
  DFF_X1 ram_reg_172__5_ ( .D(n10657), .CK(clk), .Q(ram[2757]) );
  DFF_X1 ram_reg_172__4_ ( .D(n10656), .CK(clk), .Q(ram[2756]) );
  DFF_X1 ram_reg_172__3_ ( .D(n10655), .CK(clk), .Q(ram[2755]) );
  DFF_X1 ram_reg_172__2_ ( .D(n10654), .CK(clk), .Q(ram[2754]) );
  DFF_X1 ram_reg_172__1_ ( .D(n10653), .CK(clk), .Q(ram[2753]) );
  DFF_X1 ram_reg_172__0_ ( .D(n10652), .CK(clk), .Q(ram[2752]) );
  DFF_X1 ram_reg_171__15_ ( .D(n10684), .CK(clk), .Q(ram[2751]) );
  DFF_X1 ram_reg_171__14_ ( .D(n10683), .CK(clk), .Q(ram[2750]) );
  DFF_X1 ram_reg_171__13_ ( .D(n10682), .CK(clk), .Q(ram[2749]) );
  DFF_X1 ram_reg_171__12_ ( .D(n10681), .CK(clk), .Q(ram[2748]) );
  DFF_X1 ram_reg_171__11_ ( .D(n10680), .CK(clk), .Q(ram[2747]) );
  DFF_X1 ram_reg_171__10_ ( .D(n10679), .CK(clk), .Q(ram[2746]) );
  DFF_X1 ram_reg_171__9_ ( .D(n10678), .CK(clk), .Q(ram[2745]) );
  DFF_X1 ram_reg_171__8_ ( .D(n10677), .CK(clk), .Q(ram[2744]) );
  DFF_X1 ram_reg_171__7_ ( .D(n10676), .CK(clk), .Q(ram[2743]) );
  DFF_X1 ram_reg_171__6_ ( .D(n10675), .CK(clk), .Q(ram[2742]) );
  DFF_X1 ram_reg_171__5_ ( .D(n10674), .CK(clk), .Q(ram[2741]) );
  DFF_X1 ram_reg_171__4_ ( .D(n10673), .CK(clk), .Q(ram[2740]) );
  DFF_X1 ram_reg_171__3_ ( .D(n10672), .CK(clk), .Q(ram[2739]) );
  DFF_X1 ram_reg_171__2_ ( .D(n10671), .CK(clk), .Q(ram[2738]) );
  DFF_X1 ram_reg_171__1_ ( .D(n10670), .CK(clk), .Q(ram[2737]) );
  DFF_X1 ram_reg_171__0_ ( .D(n10669), .CK(clk), .Q(ram[2736]) );
  DFF_X1 ram_reg_170__15_ ( .D(n10701), .CK(clk), .Q(ram[2735]) );
  DFF_X1 ram_reg_170__14_ ( .D(n10700), .CK(clk), .Q(ram[2734]) );
  DFF_X1 ram_reg_170__13_ ( .D(n10699), .CK(clk), .Q(ram[2733]) );
  DFF_X1 ram_reg_170__12_ ( .D(n10698), .CK(clk), .Q(ram[2732]) );
  DFF_X1 ram_reg_170__11_ ( .D(n10697), .CK(clk), .Q(ram[2731]) );
  DFF_X1 ram_reg_170__10_ ( .D(n10696), .CK(clk), .Q(ram[2730]) );
  DFF_X1 ram_reg_170__9_ ( .D(n10695), .CK(clk), .Q(ram[2729]) );
  DFF_X1 ram_reg_170__8_ ( .D(n10694), .CK(clk), .Q(ram[2728]) );
  DFF_X1 ram_reg_170__7_ ( .D(n10693), .CK(clk), .Q(ram[2727]) );
  DFF_X1 ram_reg_170__6_ ( .D(n10692), .CK(clk), .Q(ram[2726]) );
  DFF_X1 ram_reg_170__5_ ( .D(n10691), .CK(clk), .Q(ram[2725]) );
  DFF_X1 ram_reg_170__4_ ( .D(n10690), .CK(clk), .Q(ram[2724]) );
  DFF_X1 ram_reg_170__3_ ( .D(n10689), .CK(clk), .Q(ram[2723]) );
  DFF_X1 ram_reg_170__2_ ( .D(n10688), .CK(clk), .Q(ram[2722]) );
  DFF_X1 ram_reg_170__1_ ( .D(n10687), .CK(clk), .Q(ram[2721]) );
  DFF_X1 ram_reg_170__0_ ( .D(n10686), .CK(clk), .Q(ram[2720]) );
  DFF_X1 ram_reg_169__15_ ( .D(n10718), .CK(clk), .Q(ram[2719]) );
  DFF_X1 ram_reg_169__14_ ( .D(n10717), .CK(clk), .Q(ram[2718]) );
  DFF_X1 ram_reg_169__13_ ( .D(n10716), .CK(clk), .Q(ram[2717]) );
  DFF_X1 ram_reg_169__12_ ( .D(n10715), .CK(clk), .Q(ram[2716]) );
  DFF_X1 ram_reg_169__11_ ( .D(n10714), .CK(clk), .Q(ram[2715]) );
  DFF_X1 ram_reg_169__10_ ( .D(n10713), .CK(clk), .Q(ram[2714]) );
  DFF_X1 ram_reg_169__9_ ( .D(n10712), .CK(clk), .Q(ram[2713]) );
  DFF_X1 ram_reg_169__8_ ( .D(n10711), .CK(clk), .Q(ram[2712]) );
  DFF_X1 ram_reg_169__7_ ( .D(n10710), .CK(clk), .Q(ram[2711]) );
  DFF_X1 ram_reg_169__6_ ( .D(n10709), .CK(clk), .Q(ram[2710]) );
  DFF_X1 ram_reg_169__5_ ( .D(n10708), .CK(clk), .Q(ram[2709]) );
  DFF_X1 ram_reg_169__4_ ( .D(n10707), .CK(clk), .Q(ram[2708]) );
  DFF_X1 ram_reg_169__3_ ( .D(n10706), .CK(clk), .Q(ram[2707]) );
  DFF_X1 ram_reg_169__2_ ( .D(n10705), .CK(clk), .Q(ram[2706]) );
  DFF_X1 ram_reg_169__1_ ( .D(n10704), .CK(clk), .Q(ram[2705]) );
  DFF_X1 ram_reg_169__0_ ( .D(n10703), .CK(clk), .Q(ram[2704]) );
  DFF_X1 ram_reg_168__15_ ( .D(n10735), .CK(clk), .Q(ram[2703]) );
  DFF_X1 ram_reg_168__14_ ( .D(n10734), .CK(clk), .Q(ram[2702]) );
  DFF_X1 ram_reg_168__13_ ( .D(n10733), .CK(clk), .Q(ram[2701]) );
  DFF_X1 ram_reg_168__12_ ( .D(n10732), .CK(clk), .Q(ram[2700]) );
  DFF_X1 ram_reg_168__11_ ( .D(n10731), .CK(clk), .Q(ram[2699]) );
  DFF_X1 ram_reg_168__10_ ( .D(n10730), .CK(clk), .Q(ram[2698]) );
  DFF_X1 ram_reg_168__9_ ( .D(n10729), .CK(clk), .Q(ram[2697]) );
  DFF_X1 ram_reg_168__8_ ( .D(n10728), .CK(clk), .Q(ram[2696]) );
  DFF_X1 ram_reg_168__7_ ( .D(n10727), .CK(clk), .Q(ram[2695]) );
  DFF_X1 ram_reg_168__6_ ( .D(n10726), .CK(clk), .Q(ram[2694]) );
  DFF_X1 ram_reg_168__5_ ( .D(n10725), .CK(clk), .Q(ram[2693]) );
  DFF_X1 ram_reg_168__4_ ( .D(n10724), .CK(clk), .Q(ram[2692]) );
  DFF_X1 ram_reg_168__3_ ( .D(n10723), .CK(clk), .Q(ram[2691]) );
  DFF_X1 ram_reg_168__2_ ( .D(n10722), .CK(clk), .Q(ram[2690]) );
  DFF_X1 ram_reg_168__1_ ( .D(n10721), .CK(clk), .Q(ram[2689]) );
  DFF_X1 ram_reg_168__0_ ( .D(n10720), .CK(clk), .Q(ram[2688]) );
  DFF_X1 ram_reg_167__15_ ( .D(n10752), .CK(clk), .Q(ram[2687]) );
  DFF_X1 ram_reg_167__14_ ( .D(n10751), .CK(clk), .Q(ram[2686]) );
  DFF_X1 ram_reg_167__13_ ( .D(n10750), .CK(clk), .Q(ram[2685]) );
  DFF_X1 ram_reg_167__12_ ( .D(n10749), .CK(clk), .Q(ram[2684]) );
  DFF_X1 ram_reg_167__11_ ( .D(n10748), .CK(clk), .Q(ram[2683]) );
  DFF_X1 ram_reg_167__10_ ( .D(n10747), .CK(clk), .Q(ram[2682]) );
  DFF_X1 ram_reg_167__9_ ( .D(n10746), .CK(clk), .Q(ram[2681]) );
  DFF_X1 ram_reg_167__8_ ( .D(n10745), .CK(clk), .Q(ram[2680]) );
  DFF_X1 ram_reg_167__7_ ( .D(n10744), .CK(clk), .Q(ram[2679]) );
  DFF_X1 ram_reg_167__6_ ( .D(n10743), .CK(clk), .Q(ram[2678]) );
  DFF_X1 ram_reg_167__5_ ( .D(n10742), .CK(clk), .Q(ram[2677]) );
  DFF_X1 ram_reg_167__4_ ( .D(n10741), .CK(clk), .Q(ram[2676]) );
  DFF_X1 ram_reg_167__3_ ( .D(n10740), .CK(clk), .Q(ram[2675]) );
  DFF_X1 ram_reg_167__2_ ( .D(n10739), .CK(clk), .Q(ram[2674]) );
  DFF_X1 ram_reg_167__1_ ( .D(n10738), .CK(clk), .Q(ram[2673]) );
  DFF_X1 ram_reg_167__0_ ( .D(n10737), .CK(clk), .Q(ram[2672]) );
  DFF_X1 ram_reg_166__15_ ( .D(n10769), .CK(clk), .Q(ram[2671]) );
  DFF_X1 ram_reg_166__14_ ( .D(n10768), .CK(clk), .Q(ram[2670]) );
  DFF_X1 ram_reg_166__13_ ( .D(n10767), .CK(clk), .Q(ram[2669]) );
  DFF_X1 ram_reg_166__12_ ( .D(n10766), .CK(clk), .Q(ram[2668]) );
  DFF_X1 ram_reg_166__11_ ( .D(n10765), .CK(clk), .Q(ram[2667]) );
  DFF_X1 ram_reg_166__10_ ( .D(n10764), .CK(clk), .Q(ram[2666]) );
  DFF_X1 ram_reg_166__9_ ( .D(n10763), .CK(clk), .Q(ram[2665]) );
  DFF_X1 ram_reg_166__8_ ( .D(n10762), .CK(clk), .Q(ram[2664]) );
  DFF_X1 ram_reg_166__7_ ( .D(n10761), .CK(clk), .Q(ram[2663]) );
  DFF_X1 ram_reg_166__6_ ( .D(n10760), .CK(clk), .Q(ram[2662]) );
  DFF_X1 ram_reg_166__5_ ( .D(n10759), .CK(clk), .Q(ram[2661]) );
  DFF_X1 ram_reg_166__4_ ( .D(n10758), .CK(clk), .Q(ram[2660]) );
  DFF_X1 ram_reg_166__3_ ( .D(n10757), .CK(clk), .Q(ram[2659]) );
  DFF_X1 ram_reg_166__2_ ( .D(n10756), .CK(clk), .Q(ram[2658]) );
  DFF_X1 ram_reg_166__1_ ( .D(n10755), .CK(clk), .Q(ram[2657]) );
  DFF_X1 ram_reg_166__0_ ( .D(n10754), .CK(clk), .Q(ram[2656]) );
  DFF_X1 ram_reg_165__15_ ( .D(n10786), .CK(clk), .Q(ram[2655]) );
  DFF_X1 ram_reg_165__14_ ( .D(n10785), .CK(clk), .Q(ram[2654]) );
  DFF_X1 ram_reg_165__13_ ( .D(n10784), .CK(clk), .Q(ram[2653]) );
  DFF_X1 ram_reg_165__12_ ( .D(n10783), .CK(clk), .Q(ram[2652]) );
  DFF_X1 ram_reg_165__11_ ( .D(n10782), .CK(clk), .Q(ram[2651]) );
  DFF_X1 ram_reg_165__10_ ( .D(n10781), .CK(clk), .Q(ram[2650]) );
  DFF_X1 ram_reg_165__9_ ( .D(n10780), .CK(clk), .Q(ram[2649]) );
  DFF_X1 ram_reg_165__8_ ( .D(n10779), .CK(clk), .Q(ram[2648]) );
  DFF_X1 ram_reg_165__7_ ( .D(n10778), .CK(clk), .Q(ram[2647]) );
  DFF_X1 ram_reg_165__6_ ( .D(n10777), .CK(clk), .Q(ram[2646]) );
  DFF_X1 ram_reg_165__5_ ( .D(n10776), .CK(clk), .Q(ram[2645]) );
  DFF_X1 ram_reg_165__4_ ( .D(n10775), .CK(clk), .Q(ram[2644]) );
  DFF_X1 ram_reg_165__3_ ( .D(n10774), .CK(clk), .Q(ram[2643]) );
  DFF_X1 ram_reg_165__2_ ( .D(n10773), .CK(clk), .Q(ram[2642]) );
  DFF_X1 ram_reg_165__1_ ( .D(n10772), .CK(clk), .Q(ram[2641]) );
  DFF_X1 ram_reg_165__0_ ( .D(n10771), .CK(clk), .Q(ram[2640]) );
  DFF_X1 ram_reg_164__15_ ( .D(n10803), .CK(clk), .Q(ram[2639]) );
  DFF_X1 ram_reg_164__14_ ( .D(n10802), .CK(clk), .Q(ram[2638]) );
  DFF_X1 ram_reg_164__13_ ( .D(n10801), .CK(clk), .Q(ram[2637]) );
  DFF_X1 ram_reg_164__12_ ( .D(n10800), .CK(clk), .Q(ram[2636]) );
  DFF_X1 ram_reg_164__11_ ( .D(n10799), .CK(clk), .Q(ram[2635]) );
  DFF_X1 ram_reg_164__10_ ( .D(n10798), .CK(clk), .Q(ram[2634]) );
  DFF_X1 ram_reg_164__9_ ( .D(n10797), .CK(clk), .Q(ram[2633]) );
  DFF_X1 ram_reg_164__8_ ( .D(n10796), .CK(clk), .Q(ram[2632]) );
  DFF_X1 ram_reg_164__7_ ( .D(n10795), .CK(clk), .Q(ram[2631]) );
  DFF_X1 ram_reg_164__6_ ( .D(n10794), .CK(clk), .Q(ram[2630]) );
  DFF_X1 ram_reg_164__5_ ( .D(n10793), .CK(clk), .Q(ram[2629]) );
  DFF_X1 ram_reg_164__4_ ( .D(n10792), .CK(clk), .Q(ram[2628]) );
  DFF_X1 ram_reg_164__3_ ( .D(n10791), .CK(clk), .Q(ram[2627]) );
  DFF_X1 ram_reg_164__2_ ( .D(n10790), .CK(clk), .Q(ram[2626]) );
  DFF_X1 ram_reg_164__1_ ( .D(n10789), .CK(clk), .Q(ram[2625]) );
  DFF_X1 ram_reg_164__0_ ( .D(n10788), .CK(clk), .Q(ram[2624]) );
  DFF_X1 ram_reg_163__15_ ( .D(n10820), .CK(clk), .Q(ram[2623]) );
  DFF_X1 ram_reg_163__14_ ( .D(n10819), .CK(clk), .Q(ram[2622]) );
  DFF_X1 ram_reg_163__13_ ( .D(n10818), .CK(clk), .Q(ram[2621]) );
  DFF_X1 ram_reg_163__12_ ( .D(n10817), .CK(clk), .Q(ram[2620]) );
  DFF_X1 ram_reg_163__11_ ( .D(n10816), .CK(clk), .Q(ram[2619]) );
  DFF_X1 ram_reg_163__10_ ( .D(n10815), .CK(clk), .Q(ram[2618]) );
  DFF_X1 ram_reg_163__9_ ( .D(n10814), .CK(clk), .Q(ram[2617]) );
  DFF_X1 ram_reg_163__8_ ( .D(n10813), .CK(clk), .Q(ram[2616]) );
  DFF_X1 ram_reg_163__7_ ( .D(n10812), .CK(clk), .Q(ram[2615]) );
  DFF_X1 ram_reg_163__6_ ( .D(n10811), .CK(clk), .Q(ram[2614]) );
  DFF_X1 ram_reg_163__5_ ( .D(n10810), .CK(clk), .Q(ram[2613]) );
  DFF_X1 ram_reg_163__4_ ( .D(n10809), .CK(clk), .Q(ram[2612]) );
  DFF_X1 ram_reg_163__3_ ( .D(n10808), .CK(clk), .Q(ram[2611]) );
  DFF_X1 ram_reg_163__2_ ( .D(n10807), .CK(clk), .Q(ram[2610]) );
  DFF_X1 ram_reg_163__1_ ( .D(n10806), .CK(clk), .Q(ram[2609]) );
  DFF_X1 ram_reg_163__0_ ( .D(n10805), .CK(clk), .Q(ram[2608]) );
  DFF_X1 ram_reg_162__15_ ( .D(n10837), .CK(clk), .Q(ram[2607]) );
  DFF_X1 ram_reg_162__14_ ( .D(n10836), .CK(clk), .Q(ram[2606]) );
  DFF_X1 ram_reg_162__13_ ( .D(n10835), .CK(clk), .Q(ram[2605]) );
  DFF_X1 ram_reg_162__12_ ( .D(n10834), .CK(clk), .Q(ram[2604]) );
  DFF_X1 ram_reg_162__11_ ( .D(n10833), .CK(clk), .Q(ram[2603]) );
  DFF_X1 ram_reg_162__10_ ( .D(n10832), .CK(clk), .Q(ram[2602]) );
  DFF_X1 ram_reg_162__9_ ( .D(n10831), .CK(clk), .Q(ram[2601]) );
  DFF_X1 ram_reg_162__8_ ( .D(n10830), .CK(clk), .Q(ram[2600]) );
  DFF_X1 ram_reg_162__7_ ( .D(n10829), .CK(clk), .Q(ram[2599]) );
  DFF_X1 ram_reg_162__6_ ( .D(n10828), .CK(clk), .Q(ram[2598]) );
  DFF_X1 ram_reg_162__5_ ( .D(n10827), .CK(clk), .Q(ram[2597]) );
  DFF_X1 ram_reg_162__4_ ( .D(n10826), .CK(clk), .Q(ram[2596]) );
  DFF_X1 ram_reg_162__3_ ( .D(n10825), .CK(clk), .Q(ram[2595]) );
  DFF_X1 ram_reg_162__2_ ( .D(n10824), .CK(clk), .Q(ram[2594]) );
  DFF_X1 ram_reg_162__1_ ( .D(n10823), .CK(clk), .Q(ram[2593]) );
  DFF_X1 ram_reg_162__0_ ( .D(n10822), .CK(clk), .Q(ram[2592]) );
  DFF_X1 ram_reg_161__15_ ( .D(n10854), .CK(clk), .Q(ram[2591]) );
  DFF_X1 ram_reg_161__14_ ( .D(n10853), .CK(clk), .Q(ram[2590]) );
  DFF_X1 ram_reg_161__13_ ( .D(n10852), .CK(clk), .Q(ram[2589]) );
  DFF_X1 ram_reg_161__12_ ( .D(n10851), .CK(clk), .Q(ram[2588]) );
  DFF_X1 ram_reg_161__11_ ( .D(n10850), .CK(clk), .Q(ram[2587]) );
  DFF_X1 ram_reg_161__10_ ( .D(n10849), .CK(clk), .Q(ram[2586]) );
  DFF_X1 ram_reg_161__9_ ( .D(n10848), .CK(clk), .Q(ram[2585]) );
  DFF_X1 ram_reg_161__8_ ( .D(n10847), .CK(clk), .Q(ram[2584]) );
  DFF_X1 ram_reg_161__7_ ( .D(n10846), .CK(clk), .Q(ram[2583]) );
  DFF_X1 ram_reg_161__6_ ( .D(n10845), .CK(clk), .Q(ram[2582]) );
  DFF_X1 ram_reg_161__5_ ( .D(n10844), .CK(clk), .Q(ram[2581]) );
  DFF_X1 ram_reg_161__4_ ( .D(n10843), .CK(clk), .Q(ram[2580]) );
  DFF_X1 ram_reg_161__3_ ( .D(n10842), .CK(clk), .Q(ram[2579]) );
  DFF_X1 ram_reg_161__2_ ( .D(n10841), .CK(clk), .Q(ram[2578]) );
  DFF_X1 ram_reg_161__1_ ( .D(n10840), .CK(clk), .Q(ram[2577]) );
  DFF_X1 ram_reg_161__0_ ( .D(n10839), .CK(clk), .Q(ram[2576]) );
  DFF_X1 ram_reg_160__15_ ( .D(n10871), .CK(clk), .Q(ram[2575]) );
  DFF_X1 ram_reg_160__14_ ( .D(n10870), .CK(clk), .Q(ram[2574]) );
  DFF_X1 ram_reg_160__13_ ( .D(n10869), .CK(clk), .Q(ram[2573]) );
  DFF_X1 ram_reg_160__12_ ( .D(n10868), .CK(clk), .Q(ram[2572]) );
  DFF_X1 ram_reg_160__11_ ( .D(n10867), .CK(clk), .Q(ram[2571]) );
  DFF_X1 ram_reg_160__10_ ( .D(n10866), .CK(clk), .Q(ram[2570]) );
  DFF_X1 ram_reg_160__9_ ( .D(n10865), .CK(clk), .Q(ram[2569]) );
  DFF_X1 ram_reg_160__8_ ( .D(n10864), .CK(clk), .Q(ram[2568]) );
  DFF_X1 ram_reg_160__7_ ( .D(n10863), .CK(clk), .Q(ram[2567]) );
  DFF_X1 ram_reg_160__6_ ( .D(n10862), .CK(clk), .Q(ram[2566]) );
  DFF_X1 ram_reg_160__5_ ( .D(n10861), .CK(clk), .Q(ram[2565]) );
  DFF_X1 ram_reg_160__4_ ( .D(n10860), .CK(clk), .Q(ram[2564]) );
  DFF_X1 ram_reg_160__3_ ( .D(n10859), .CK(clk), .Q(ram[2563]) );
  DFF_X1 ram_reg_160__2_ ( .D(n10858), .CK(clk), .Q(ram[2562]) );
  DFF_X1 ram_reg_160__1_ ( .D(n10857), .CK(clk), .Q(ram[2561]) );
  DFF_X1 ram_reg_160__0_ ( .D(n10856), .CK(clk), .Q(ram[2560]) );
  DFF_X1 ram_reg_159__15_ ( .D(n10888), .CK(clk), .Q(ram[2559]) );
  DFF_X1 ram_reg_159__14_ ( .D(n10887), .CK(clk), .Q(ram[2558]) );
  DFF_X1 ram_reg_159__13_ ( .D(n10886), .CK(clk), .Q(ram[2557]) );
  DFF_X1 ram_reg_159__12_ ( .D(n10885), .CK(clk), .Q(ram[2556]) );
  DFF_X1 ram_reg_159__11_ ( .D(n10884), .CK(clk), .Q(ram[2555]) );
  DFF_X1 ram_reg_159__10_ ( .D(n10883), .CK(clk), .Q(ram[2554]) );
  DFF_X1 ram_reg_159__9_ ( .D(n10882), .CK(clk), .Q(ram[2553]) );
  DFF_X1 ram_reg_159__8_ ( .D(n10881), .CK(clk), .Q(ram[2552]) );
  DFF_X1 ram_reg_159__7_ ( .D(n10880), .CK(clk), .Q(ram[2551]) );
  DFF_X1 ram_reg_159__6_ ( .D(n10879), .CK(clk), .Q(ram[2550]) );
  DFF_X1 ram_reg_159__5_ ( .D(n10878), .CK(clk), .Q(ram[2549]) );
  DFF_X1 ram_reg_159__4_ ( .D(n10877), .CK(clk), .Q(ram[2548]) );
  DFF_X1 ram_reg_159__3_ ( .D(n10876), .CK(clk), .Q(ram[2547]) );
  DFF_X1 ram_reg_159__2_ ( .D(n10875), .CK(clk), .Q(ram[2546]) );
  DFF_X1 ram_reg_159__1_ ( .D(n10874), .CK(clk), .Q(ram[2545]) );
  DFF_X1 ram_reg_159__0_ ( .D(n10873), .CK(clk), .Q(ram[2544]) );
  DFF_X1 ram_reg_158__15_ ( .D(n10905), .CK(clk), .Q(ram[2543]) );
  DFF_X1 ram_reg_158__14_ ( .D(n10904), .CK(clk), .Q(ram[2542]) );
  DFF_X1 ram_reg_158__13_ ( .D(n10903), .CK(clk), .Q(ram[2541]) );
  DFF_X1 ram_reg_158__12_ ( .D(n10902), .CK(clk), .Q(ram[2540]) );
  DFF_X1 ram_reg_158__11_ ( .D(n10901), .CK(clk), .Q(ram[2539]) );
  DFF_X1 ram_reg_158__10_ ( .D(n10900), .CK(clk), .Q(ram[2538]) );
  DFF_X1 ram_reg_158__9_ ( .D(n10899), .CK(clk), .Q(ram[2537]) );
  DFF_X1 ram_reg_158__8_ ( .D(n10898), .CK(clk), .Q(ram[2536]) );
  DFF_X1 ram_reg_158__7_ ( .D(n10897), .CK(clk), .Q(ram[2535]) );
  DFF_X1 ram_reg_158__6_ ( .D(n10896), .CK(clk), .Q(ram[2534]) );
  DFF_X1 ram_reg_158__5_ ( .D(n10895), .CK(clk), .Q(ram[2533]) );
  DFF_X1 ram_reg_158__4_ ( .D(n10894), .CK(clk), .Q(ram[2532]) );
  DFF_X1 ram_reg_158__3_ ( .D(n10893), .CK(clk), .Q(ram[2531]) );
  DFF_X1 ram_reg_158__2_ ( .D(n10892), .CK(clk), .Q(ram[2530]) );
  DFF_X1 ram_reg_158__1_ ( .D(n10891), .CK(clk), .Q(ram[2529]) );
  DFF_X1 ram_reg_158__0_ ( .D(n10890), .CK(clk), .Q(ram[2528]) );
  DFF_X1 ram_reg_157__15_ ( .D(n10922), .CK(clk), .Q(ram[2527]) );
  DFF_X1 ram_reg_157__14_ ( .D(n10921), .CK(clk), .Q(ram[2526]) );
  DFF_X1 ram_reg_157__13_ ( .D(n10920), .CK(clk), .Q(ram[2525]) );
  DFF_X1 ram_reg_157__12_ ( .D(n10919), .CK(clk), .Q(ram[2524]) );
  DFF_X1 ram_reg_157__11_ ( .D(n10918), .CK(clk), .Q(ram[2523]) );
  DFF_X1 ram_reg_157__10_ ( .D(n10917), .CK(clk), .Q(ram[2522]) );
  DFF_X1 ram_reg_157__9_ ( .D(n10916), .CK(clk), .Q(ram[2521]) );
  DFF_X1 ram_reg_157__8_ ( .D(n10915), .CK(clk), .Q(ram[2520]) );
  DFF_X1 ram_reg_157__7_ ( .D(n10914), .CK(clk), .Q(ram[2519]) );
  DFF_X1 ram_reg_157__6_ ( .D(n10913), .CK(clk), .Q(ram[2518]) );
  DFF_X1 ram_reg_157__5_ ( .D(n10912), .CK(clk), .Q(ram[2517]) );
  DFF_X1 ram_reg_157__4_ ( .D(n10911), .CK(clk), .Q(ram[2516]) );
  DFF_X1 ram_reg_157__3_ ( .D(n10910), .CK(clk), .Q(ram[2515]) );
  DFF_X1 ram_reg_157__2_ ( .D(n10909), .CK(clk), .Q(ram[2514]) );
  DFF_X1 ram_reg_157__1_ ( .D(n10908), .CK(clk), .Q(ram[2513]) );
  DFF_X1 ram_reg_157__0_ ( .D(n10907), .CK(clk), .Q(ram[2512]) );
  DFF_X1 ram_reg_156__15_ ( .D(n10939), .CK(clk), .Q(ram[2511]) );
  DFF_X1 ram_reg_156__14_ ( .D(n10938), .CK(clk), .Q(ram[2510]) );
  DFF_X1 ram_reg_156__13_ ( .D(n10937), .CK(clk), .Q(ram[2509]) );
  DFF_X1 ram_reg_156__12_ ( .D(n10936), .CK(clk), .Q(ram[2508]) );
  DFF_X1 ram_reg_156__11_ ( .D(n10935), .CK(clk), .Q(ram[2507]) );
  DFF_X1 ram_reg_156__10_ ( .D(n10934), .CK(clk), .Q(ram[2506]) );
  DFF_X1 ram_reg_156__9_ ( .D(n10933), .CK(clk), .Q(ram[2505]) );
  DFF_X1 ram_reg_156__8_ ( .D(n10932), .CK(clk), .Q(ram[2504]) );
  DFF_X1 ram_reg_156__7_ ( .D(n10931), .CK(clk), .Q(ram[2503]) );
  DFF_X1 ram_reg_156__6_ ( .D(n10930), .CK(clk), .Q(ram[2502]) );
  DFF_X1 ram_reg_156__5_ ( .D(n10929), .CK(clk), .Q(ram[2501]) );
  DFF_X1 ram_reg_156__4_ ( .D(n10928), .CK(clk), .Q(ram[2500]) );
  DFF_X1 ram_reg_156__3_ ( .D(n10927), .CK(clk), .Q(ram[2499]) );
  DFF_X1 ram_reg_156__2_ ( .D(n10926), .CK(clk), .Q(ram[2498]) );
  DFF_X1 ram_reg_156__1_ ( .D(n10925), .CK(clk), .Q(ram[2497]) );
  DFF_X1 ram_reg_156__0_ ( .D(n10924), .CK(clk), .Q(ram[2496]) );
  DFF_X1 ram_reg_155__15_ ( .D(n10956), .CK(clk), .Q(ram[2495]) );
  DFF_X1 ram_reg_155__14_ ( .D(n10955), .CK(clk), .Q(ram[2494]) );
  DFF_X1 ram_reg_155__13_ ( .D(n10954), .CK(clk), .Q(ram[2493]) );
  DFF_X1 ram_reg_155__12_ ( .D(n10953), .CK(clk), .Q(ram[2492]) );
  DFF_X1 ram_reg_155__11_ ( .D(n10952), .CK(clk), .Q(ram[2491]) );
  DFF_X1 ram_reg_155__10_ ( .D(n10951), .CK(clk), .Q(ram[2490]) );
  DFF_X1 ram_reg_155__9_ ( .D(n10950), .CK(clk), .Q(ram[2489]) );
  DFF_X1 ram_reg_155__8_ ( .D(n10949), .CK(clk), .Q(ram[2488]) );
  DFF_X1 ram_reg_155__7_ ( .D(n10948), .CK(clk), .Q(ram[2487]) );
  DFF_X1 ram_reg_155__6_ ( .D(n10947), .CK(clk), .Q(ram[2486]) );
  DFF_X1 ram_reg_155__5_ ( .D(n10946), .CK(clk), .Q(ram[2485]) );
  DFF_X1 ram_reg_155__4_ ( .D(n10945), .CK(clk), .Q(ram[2484]) );
  DFF_X1 ram_reg_155__3_ ( .D(n10944), .CK(clk), .Q(ram[2483]) );
  DFF_X1 ram_reg_155__2_ ( .D(n10943), .CK(clk), .Q(ram[2482]) );
  DFF_X1 ram_reg_155__1_ ( .D(n10942), .CK(clk), .Q(ram[2481]) );
  DFF_X1 ram_reg_155__0_ ( .D(n10941), .CK(clk), .Q(ram[2480]) );
  DFF_X1 ram_reg_154__15_ ( .D(n10973), .CK(clk), .Q(ram[2479]) );
  DFF_X1 ram_reg_154__14_ ( .D(n10972), .CK(clk), .Q(ram[2478]) );
  DFF_X1 ram_reg_154__13_ ( .D(n10971), .CK(clk), .Q(ram[2477]) );
  DFF_X1 ram_reg_154__12_ ( .D(n10970), .CK(clk), .Q(ram[2476]) );
  DFF_X1 ram_reg_154__11_ ( .D(n10969), .CK(clk), .Q(ram[2475]) );
  DFF_X1 ram_reg_154__10_ ( .D(n10968), .CK(clk), .Q(ram[2474]) );
  DFF_X1 ram_reg_154__9_ ( .D(n10967), .CK(clk), .Q(ram[2473]) );
  DFF_X1 ram_reg_154__8_ ( .D(n10966), .CK(clk), .Q(ram[2472]) );
  DFF_X1 ram_reg_154__7_ ( .D(n10965), .CK(clk), .Q(ram[2471]) );
  DFF_X1 ram_reg_154__6_ ( .D(n10964), .CK(clk), .Q(ram[2470]) );
  DFF_X1 ram_reg_154__5_ ( .D(n10963), .CK(clk), .Q(ram[2469]) );
  DFF_X1 ram_reg_154__4_ ( .D(n10962), .CK(clk), .Q(ram[2468]) );
  DFF_X1 ram_reg_154__3_ ( .D(n10961), .CK(clk), .Q(ram[2467]) );
  DFF_X1 ram_reg_154__2_ ( .D(n10960), .CK(clk), .Q(ram[2466]) );
  DFF_X1 ram_reg_154__1_ ( .D(n10959), .CK(clk), .Q(ram[2465]) );
  DFF_X1 ram_reg_154__0_ ( .D(n10958), .CK(clk), .Q(ram[2464]) );
  DFF_X1 ram_reg_153__15_ ( .D(n10990), .CK(clk), .Q(ram[2463]) );
  DFF_X1 ram_reg_153__14_ ( .D(n10989), .CK(clk), .Q(ram[2462]) );
  DFF_X1 ram_reg_153__13_ ( .D(n10988), .CK(clk), .Q(ram[2461]) );
  DFF_X1 ram_reg_153__12_ ( .D(n10987), .CK(clk), .Q(ram[2460]) );
  DFF_X1 ram_reg_153__11_ ( .D(n10986), .CK(clk), .Q(ram[2459]) );
  DFF_X1 ram_reg_153__10_ ( .D(n10985), .CK(clk), .Q(ram[2458]) );
  DFF_X1 ram_reg_153__9_ ( .D(n10984), .CK(clk), .Q(ram[2457]) );
  DFF_X1 ram_reg_153__8_ ( .D(n10983), .CK(clk), .Q(ram[2456]) );
  DFF_X1 ram_reg_153__7_ ( .D(n10982), .CK(clk), .Q(ram[2455]) );
  DFF_X1 ram_reg_153__6_ ( .D(n10981), .CK(clk), .Q(ram[2454]) );
  DFF_X1 ram_reg_153__5_ ( .D(n10980), .CK(clk), .Q(ram[2453]) );
  DFF_X1 ram_reg_153__4_ ( .D(n10979), .CK(clk), .Q(ram[2452]) );
  DFF_X1 ram_reg_153__3_ ( .D(n10978), .CK(clk), .Q(ram[2451]) );
  DFF_X1 ram_reg_153__2_ ( .D(n10977), .CK(clk), .Q(ram[2450]) );
  DFF_X1 ram_reg_153__1_ ( .D(n10976), .CK(clk), .Q(ram[2449]) );
  DFF_X1 ram_reg_153__0_ ( .D(n10975), .CK(clk), .Q(ram[2448]) );
  DFF_X1 ram_reg_152__15_ ( .D(n11007), .CK(clk), .Q(ram[2447]) );
  DFF_X1 ram_reg_152__14_ ( .D(n11006), .CK(clk), .Q(ram[2446]) );
  DFF_X1 ram_reg_152__13_ ( .D(n11005), .CK(clk), .Q(ram[2445]) );
  DFF_X1 ram_reg_152__12_ ( .D(n11004), .CK(clk), .Q(ram[2444]) );
  DFF_X1 ram_reg_152__11_ ( .D(n11003), .CK(clk), .Q(ram[2443]) );
  DFF_X1 ram_reg_152__10_ ( .D(n11002), .CK(clk), .Q(ram[2442]) );
  DFF_X1 ram_reg_152__9_ ( .D(n11001), .CK(clk), .Q(ram[2441]) );
  DFF_X1 ram_reg_152__8_ ( .D(n11000), .CK(clk), .Q(ram[2440]) );
  DFF_X1 ram_reg_152__7_ ( .D(n10999), .CK(clk), .Q(ram[2439]) );
  DFF_X1 ram_reg_152__6_ ( .D(n10998), .CK(clk), .Q(ram[2438]) );
  DFF_X1 ram_reg_152__5_ ( .D(n10997), .CK(clk), .Q(ram[2437]) );
  DFF_X1 ram_reg_152__4_ ( .D(n10996), .CK(clk), .Q(ram[2436]) );
  DFF_X1 ram_reg_152__3_ ( .D(n10995), .CK(clk), .Q(ram[2435]) );
  DFF_X1 ram_reg_152__2_ ( .D(n10994), .CK(clk), .Q(ram[2434]) );
  DFF_X1 ram_reg_152__1_ ( .D(n10993), .CK(clk), .Q(ram[2433]) );
  DFF_X1 ram_reg_152__0_ ( .D(n10992), .CK(clk), .Q(ram[2432]) );
  DFF_X1 ram_reg_151__15_ ( .D(n11024), .CK(clk), .Q(ram[2431]) );
  DFF_X1 ram_reg_151__14_ ( .D(n11023), .CK(clk), .Q(ram[2430]) );
  DFF_X1 ram_reg_151__13_ ( .D(n11022), .CK(clk), .Q(ram[2429]) );
  DFF_X1 ram_reg_151__12_ ( .D(n11021), .CK(clk), .Q(ram[2428]) );
  DFF_X1 ram_reg_151__11_ ( .D(n11020), .CK(clk), .Q(ram[2427]) );
  DFF_X1 ram_reg_151__10_ ( .D(n11019), .CK(clk), .Q(ram[2426]) );
  DFF_X1 ram_reg_151__9_ ( .D(n11018), .CK(clk), .Q(ram[2425]) );
  DFF_X1 ram_reg_151__8_ ( .D(n11017), .CK(clk), .Q(ram[2424]) );
  DFF_X1 ram_reg_151__7_ ( .D(n11016), .CK(clk), .Q(ram[2423]) );
  DFF_X1 ram_reg_151__6_ ( .D(n11015), .CK(clk), .Q(ram[2422]) );
  DFF_X1 ram_reg_151__5_ ( .D(n11014), .CK(clk), .Q(ram[2421]) );
  DFF_X1 ram_reg_151__4_ ( .D(n11013), .CK(clk), .Q(ram[2420]) );
  DFF_X1 ram_reg_151__3_ ( .D(n11012), .CK(clk), .Q(ram[2419]) );
  DFF_X1 ram_reg_151__2_ ( .D(n11011), .CK(clk), .Q(ram[2418]) );
  DFF_X1 ram_reg_151__1_ ( .D(n11010), .CK(clk), .Q(ram[2417]) );
  DFF_X1 ram_reg_151__0_ ( .D(n11009), .CK(clk), .Q(ram[2416]) );
  DFF_X1 ram_reg_150__15_ ( .D(n11041), .CK(clk), .Q(ram[2415]) );
  DFF_X1 ram_reg_150__14_ ( .D(n11040), .CK(clk), .Q(ram[2414]) );
  DFF_X1 ram_reg_150__13_ ( .D(n11039), .CK(clk), .Q(ram[2413]) );
  DFF_X1 ram_reg_150__12_ ( .D(n11038), .CK(clk), .Q(ram[2412]) );
  DFF_X1 ram_reg_150__11_ ( .D(n11037), .CK(clk), .Q(ram[2411]) );
  DFF_X1 ram_reg_150__10_ ( .D(n11036), .CK(clk), .Q(ram[2410]) );
  DFF_X1 ram_reg_150__9_ ( .D(n11035), .CK(clk), .Q(ram[2409]) );
  DFF_X1 ram_reg_150__8_ ( .D(n11034), .CK(clk), .Q(ram[2408]) );
  DFF_X1 ram_reg_150__7_ ( .D(n11033), .CK(clk), .Q(ram[2407]) );
  DFF_X1 ram_reg_150__6_ ( .D(n11032), .CK(clk), .Q(ram[2406]) );
  DFF_X1 ram_reg_150__5_ ( .D(n11031), .CK(clk), .Q(ram[2405]) );
  DFF_X1 ram_reg_150__4_ ( .D(n11030), .CK(clk), .Q(ram[2404]) );
  DFF_X1 ram_reg_150__3_ ( .D(n11029), .CK(clk), .Q(ram[2403]) );
  DFF_X1 ram_reg_150__2_ ( .D(n11028), .CK(clk), .Q(ram[2402]) );
  DFF_X1 ram_reg_150__1_ ( .D(n11027), .CK(clk), .Q(ram[2401]) );
  DFF_X1 ram_reg_150__0_ ( .D(n11026), .CK(clk), .Q(ram[2400]) );
  DFF_X1 ram_reg_149__15_ ( .D(n11058), .CK(clk), .Q(ram[2399]) );
  DFF_X1 ram_reg_149__14_ ( .D(n11057), .CK(clk), .Q(ram[2398]) );
  DFF_X1 ram_reg_149__13_ ( .D(n11056), .CK(clk), .Q(ram[2397]) );
  DFF_X1 ram_reg_149__12_ ( .D(n11055), .CK(clk), .Q(ram[2396]) );
  DFF_X1 ram_reg_149__11_ ( .D(n11054), .CK(clk), .Q(ram[2395]) );
  DFF_X1 ram_reg_149__10_ ( .D(n11053), .CK(clk), .Q(ram[2394]) );
  DFF_X1 ram_reg_149__9_ ( .D(n11052), .CK(clk), .Q(ram[2393]) );
  DFF_X1 ram_reg_149__8_ ( .D(n11051), .CK(clk), .Q(ram[2392]) );
  DFF_X1 ram_reg_149__7_ ( .D(n11050), .CK(clk), .Q(ram[2391]) );
  DFF_X1 ram_reg_149__6_ ( .D(n11049), .CK(clk), .Q(ram[2390]) );
  DFF_X1 ram_reg_149__5_ ( .D(n11048), .CK(clk), .Q(ram[2389]) );
  DFF_X1 ram_reg_149__4_ ( .D(n11047), .CK(clk), .Q(ram[2388]) );
  DFF_X1 ram_reg_149__3_ ( .D(n11046), .CK(clk), .Q(ram[2387]) );
  DFF_X1 ram_reg_149__2_ ( .D(n11045), .CK(clk), .Q(ram[2386]) );
  DFF_X1 ram_reg_149__1_ ( .D(n11044), .CK(clk), .Q(ram[2385]) );
  DFF_X1 ram_reg_149__0_ ( .D(n11043), .CK(clk), .Q(ram[2384]) );
  DFF_X1 ram_reg_148__15_ ( .D(n11075), .CK(clk), .Q(ram[2383]) );
  DFF_X1 ram_reg_148__14_ ( .D(n11074), .CK(clk), .Q(ram[2382]) );
  DFF_X1 ram_reg_148__13_ ( .D(n11073), .CK(clk), .Q(ram[2381]) );
  DFF_X1 ram_reg_148__12_ ( .D(n11072), .CK(clk), .Q(ram[2380]) );
  DFF_X1 ram_reg_148__11_ ( .D(n11071), .CK(clk), .Q(ram[2379]) );
  DFF_X1 ram_reg_148__10_ ( .D(n11070), .CK(clk), .Q(ram[2378]) );
  DFF_X1 ram_reg_148__9_ ( .D(n11069), .CK(clk), .Q(ram[2377]) );
  DFF_X1 ram_reg_148__8_ ( .D(n11068), .CK(clk), .Q(ram[2376]) );
  DFF_X1 ram_reg_148__7_ ( .D(n11067), .CK(clk), .Q(ram[2375]) );
  DFF_X1 ram_reg_148__6_ ( .D(n11066), .CK(clk), .Q(ram[2374]) );
  DFF_X1 ram_reg_148__5_ ( .D(n11065), .CK(clk), .Q(ram[2373]) );
  DFF_X1 ram_reg_148__4_ ( .D(n11064), .CK(clk), .Q(ram[2372]) );
  DFF_X1 ram_reg_148__3_ ( .D(n11063), .CK(clk), .Q(ram[2371]) );
  DFF_X1 ram_reg_148__2_ ( .D(n11062), .CK(clk), .Q(ram[2370]) );
  DFF_X1 ram_reg_148__1_ ( .D(n11061), .CK(clk), .Q(ram[2369]) );
  DFF_X1 ram_reg_148__0_ ( .D(n11060), .CK(clk), .Q(ram[2368]) );
  DFF_X1 ram_reg_147__15_ ( .D(n11092), .CK(clk), .Q(ram[2367]) );
  DFF_X1 ram_reg_147__14_ ( .D(n11091), .CK(clk), .Q(ram[2366]) );
  DFF_X1 ram_reg_147__13_ ( .D(n11090), .CK(clk), .Q(ram[2365]) );
  DFF_X1 ram_reg_147__12_ ( .D(n11089), .CK(clk), .Q(ram[2364]) );
  DFF_X1 ram_reg_147__11_ ( .D(n11088), .CK(clk), .Q(ram[2363]) );
  DFF_X1 ram_reg_147__10_ ( .D(n11087), .CK(clk), .Q(ram[2362]) );
  DFF_X1 ram_reg_147__9_ ( .D(n11086), .CK(clk), .Q(ram[2361]) );
  DFF_X1 ram_reg_147__8_ ( .D(n11085), .CK(clk), .Q(ram[2360]) );
  DFF_X1 ram_reg_147__7_ ( .D(n11084), .CK(clk), .Q(ram[2359]) );
  DFF_X1 ram_reg_147__6_ ( .D(n11083), .CK(clk), .Q(ram[2358]) );
  DFF_X1 ram_reg_147__5_ ( .D(n11082), .CK(clk), .Q(ram[2357]) );
  DFF_X1 ram_reg_147__4_ ( .D(n11081), .CK(clk), .Q(ram[2356]) );
  DFF_X1 ram_reg_147__3_ ( .D(n11080), .CK(clk), .Q(ram[2355]) );
  DFF_X1 ram_reg_147__2_ ( .D(n11079), .CK(clk), .Q(ram[2354]) );
  DFF_X1 ram_reg_147__1_ ( .D(n11078), .CK(clk), .Q(ram[2353]) );
  DFF_X1 ram_reg_147__0_ ( .D(n11077), .CK(clk), .Q(ram[2352]) );
  DFF_X1 ram_reg_146__15_ ( .D(n11109), .CK(clk), .Q(ram[2351]) );
  DFF_X1 ram_reg_146__14_ ( .D(n11108), .CK(clk), .Q(ram[2350]) );
  DFF_X1 ram_reg_146__13_ ( .D(n11107), .CK(clk), .Q(ram[2349]) );
  DFF_X1 ram_reg_146__12_ ( .D(n11106), .CK(clk), .Q(ram[2348]) );
  DFF_X1 ram_reg_146__11_ ( .D(n11105), .CK(clk), .Q(ram[2347]) );
  DFF_X1 ram_reg_146__10_ ( .D(n11104), .CK(clk), .Q(ram[2346]) );
  DFF_X1 ram_reg_146__9_ ( .D(n11103), .CK(clk), .Q(ram[2345]) );
  DFF_X1 ram_reg_146__8_ ( .D(n11102), .CK(clk), .Q(ram[2344]) );
  DFF_X1 ram_reg_146__7_ ( .D(n11101), .CK(clk), .Q(ram[2343]) );
  DFF_X1 ram_reg_146__6_ ( .D(n11100), .CK(clk), .Q(ram[2342]) );
  DFF_X1 ram_reg_146__5_ ( .D(n11099), .CK(clk), .Q(ram[2341]) );
  DFF_X1 ram_reg_146__4_ ( .D(n11098), .CK(clk), .Q(ram[2340]) );
  DFF_X1 ram_reg_146__3_ ( .D(n11097), .CK(clk), .Q(ram[2339]) );
  DFF_X1 ram_reg_146__2_ ( .D(n11096), .CK(clk), .Q(ram[2338]) );
  DFF_X1 ram_reg_146__1_ ( .D(n11095), .CK(clk), .Q(ram[2337]) );
  DFF_X1 ram_reg_146__0_ ( .D(n11094), .CK(clk), .Q(ram[2336]) );
  DFF_X1 ram_reg_145__15_ ( .D(n11126), .CK(clk), .Q(ram[2335]) );
  DFF_X1 ram_reg_145__14_ ( .D(n11125), .CK(clk), .Q(ram[2334]) );
  DFF_X1 ram_reg_145__13_ ( .D(n11124), .CK(clk), .Q(ram[2333]) );
  DFF_X1 ram_reg_145__12_ ( .D(n11123), .CK(clk), .Q(ram[2332]) );
  DFF_X1 ram_reg_145__11_ ( .D(n11122), .CK(clk), .Q(ram[2331]) );
  DFF_X1 ram_reg_145__10_ ( .D(n11121), .CK(clk), .Q(ram[2330]) );
  DFF_X1 ram_reg_145__9_ ( .D(n11120), .CK(clk), .Q(ram[2329]) );
  DFF_X1 ram_reg_145__8_ ( .D(n11119), .CK(clk), .Q(ram[2328]) );
  DFF_X1 ram_reg_145__7_ ( .D(n11118), .CK(clk), .Q(ram[2327]) );
  DFF_X1 ram_reg_145__6_ ( .D(n11117), .CK(clk), .Q(ram[2326]) );
  DFF_X1 ram_reg_145__5_ ( .D(n11116), .CK(clk), .Q(ram[2325]) );
  DFF_X1 ram_reg_145__4_ ( .D(n11115), .CK(clk), .Q(ram[2324]) );
  DFF_X1 ram_reg_145__3_ ( .D(n11114), .CK(clk), .Q(ram[2323]) );
  DFF_X1 ram_reg_145__2_ ( .D(n11113), .CK(clk), .Q(ram[2322]) );
  DFF_X1 ram_reg_145__1_ ( .D(n11112), .CK(clk), .Q(ram[2321]) );
  DFF_X1 ram_reg_145__0_ ( .D(n11111), .CK(clk), .Q(ram[2320]) );
  DFF_X1 ram_reg_144__15_ ( .D(n11143), .CK(clk), .Q(ram[2319]) );
  DFF_X1 ram_reg_144__14_ ( .D(n11142), .CK(clk), .Q(ram[2318]) );
  DFF_X1 ram_reg_144__13_ ( .D(n11141), .CK(clk), .Q(ram[2317]) );
  DFF_X1 ram_reg_144__12_ ( .D(n11140), .CK(clk), .Q(ram[2316]) );
  DFF_X1 ram_reg_144__11_ ( .D(n11139), .CK(clk), .Q(ram[2315]) );
  DFF_X1 ram_reg_144__10_ ( .D(n11138), .CK(clk), .Q(ram[2314]) );
  DFF_X1 ram_reg_144__9_ ( .D(n11137), .CK(clk), .Q(ram[2313]) );
  DFF_X1 ram_reg_144__8_ ( .D(n11136), .CK(clk), .Q(ram[2312]) );
  DFF_X1 ram_reg_144__7_ ( .D(n11135), .CK(clk), .Q(ram[2311]) );
  DFF_X1 ram_reg_144__6_ ( .D(n11134), .CK(clk), .Q(ram[2310]) );
  DFF_X1 ram_reg_144__5_ ( .D(n11133), .CK(clk), .Q(ram[2309]) );
  DFF_X1 ram_reg_144__4_ ( .D(n11132), .CK(clk), .Q(ram[2308]) );
  DFF_X1 ram_reg_144__3_ ( .D(n11131), .CK(clk), .Q(ram[2307]) );
  DFF_X1 ram_reg_144__2_ ( .D(n11130), .CK(clk), .Q(ram[2306]) );
  DFF_X1 ram_reg_144__1_ ( .D(n11129), .CK(clk), .Q(ram[2305]) );
  DFF_X1 ram_reg_144__0_ ( .D(n11128), .CK(clk), .Q(ram[2304]) );
  DFF_X1 ram_reg_143__15_ ( .D(n11160), .CK(clk), .Q(ram[2303]) );
  DFF_X1 ram_reg_143__14_ ( .D(n11159), .CK(clk), .Q(ram[2302]) );
  DFF_X1 ram_reg_143__13_ ( .D(n11158), .CK(clk), .Q(ram[2301]) );
  DFF_X1 ram_reg_143__12_ ( .D(n11157), .CK(clk), .Q(ram[2300]) );
  DFF_X1 ram_reg_143__11_ ( .D(n11156), .CK(clk), .Q(ram[2299]) );
  DFF_X1 ram_reg_143__10_ ( .D(n11155), .CK(clk), .Q(ram[2298]) );
  DFF_X1 ram_reg_143__9_ ( .D(n11154), .CK(clk), .Q(ram[2297]) );
  DFF_X1 ram_reg_143__8_ ( .D(n11153), .CK(clk), .Q(ram[2296]) );
  DFF_X1 ram_reg_143__7_ ( .D(n11152), .CK(clk), .Q(ram[2295]) );
  DFF_X1 ram_reg_143__6_ ( .D(n11151), .CK(clk), .Q(ram[2294]) );
  DFF_X1 ram_reg_143__5_ ( .D(n11150), .CK(clk), .Q(ram[2293]) );
  DFF_X1 ram_reg_143__4_ ( .D(n11149), .CK(clk), .Q(ram[2292]) );
  DFF_X1 ram_reg_143__3_ ( .D(n11148), .CK(clk), .Q(ram[2291]) );
  DFF_X1 ram_reg_143__2_ ( .D(n11147), .CK(clk), .Q(ram[2290]) );
  DFF_X1 ram_reg_143__1_ ( .D(n11146), .CK(clk), .Q(ram[2289]) );
  DFF_X1 ram_reg_143__0_ ( .D(n11145), .CK(clk), .Q(ram[2288]) );
  DFF_X1 ram_reg_142__15_ ( .D(n11177), .CK(clk), .Q(ram[2287]) );
  DFF_X1 ram_reg_142__14_ ( .D(n11176), .CK(clk), .Q(ram[2286]) );
  DFF_X1 ram_reg_142__13_ ( .D(n11175), .CK(clk), .Q(ram[2285]) );
  DFF_X1 ram_reg_142__12_ ( .D(n11174), .CK(clk), .Q(ram[2284]) );
  DFF_X1 ram_reg_142__11_ ( .D(n11173), .CK(clk), .Q(ram[2283]) );
  DFF_X1 ram_reg_142__10_ ( .D(n11172), .CK(clk), .Q(ram[2282]) );
  DFF_X1 ram_reg_142__9_ ( .D(n11171), .CK(clk), .Q(ram[2281]) );
  DFF_X1 ram_reg_142__8_ ( .D(n11170), .CK(clk), .Q(ram[2280]) );
  DFF_X1 ram_reg_142__7_ ( .D(n11169), .CK(clk), .Q(ram[2279]) );
  DFF_X1 ram_reg_142__6_ ( .D(n11168), .CK(clk), .Q(ram[2278]) );
  DFF_X1 ram_reg_142__5_ ( .D(n11167), .CK(clk), .Q(ram[2277]) );
  DFF_X1 ram_reg_142__4_ ( .D(n11166), .CK(clk), .Q(ram[2276]) );
  DFF_X1 ram_reg_142__3_ ( .D(n11165), .CK(clk), .Q(ram[2275]) );
  DFF_X1 ram_reg_142__2_ ( .D(n11164), .CK(clk), .Q(ram[2274]) );
  DFF_X1 ram_reg_142__1_ ( .D(n11163), .CK(clk), .Q(ram[2273]) );
  DFF_X1 ram_reg_142__0_ ( .D(n11162), .CK(clk), .Q(ram[2272]) );
  DFF_X1 ram_reg_141__15_ ( .D(n11194), .CK(clk), .Q(ram[2271]) );
  DFF_X1 ram_reg_141__14_ ( .D(n11193), .CK(clk), .Q(ram[2270]) );
  DFF_X1 ram_reg_141__13_ ( .D(n11192), .CK(clk), .Q(ram[2269]) );
  DFF_X1 ram_reg_141__12_ ( .D(n11191), .CK(clk), .Q(ram[2268]) );
  DFF_X1 ram_reg_141__11_ ( .D(n11190), .CK(clk), .Q(ram[2267]) );
  DFF_X1 ram_reg_141__10_ ( .D(n11189), .CK(clk), .Q(ram[2266]) );
  DFF_X1 ram_reg_141__9_ ( .D(n11188), .CK(clk), .Q(ram[2265]) );
  DFF_X1 ram_reg_141__8_ ( .D(n11187), .CK(clk), .Q(ram[2264]) );
  DFF_X1 ram_reg_141__7_ ( .D(n11186), .CK(clk), .Q(ram[2263]) );
  DFF_X1 ram_reg_141__6_ ( .D(n11185), .CK(clk), .Q(ram[2262]) );
  DFF_X1 ram_reg_141__5_ ( .D(n11184), .CK(clk), .Q(ram[2261]) );
  DFF_X1 ram_reg_141__4_ ( .D(n11183), .CK(clk), .Q(ram[2260]) );
  DFF_X1 ram_reg_141__3_ ( .D(n11182), .CK(clk), .Q(ram[2259]) );
  DFF_X1 ram_reg_141__2_ ( .D(n11181), .CK(clk), .Q(ram[2258]) );
  DFF_X1 ram_reg_141__1_ ( .D(n11180), .CK(clk), .Q(ram[2257]) );
  DFF_X1 ram_reg_141__0_ ( .D(n11179), .CK(clk), .Q(ram[2256]) );
  DFF_X1 ram_reg_140__15_ ( .D(n11211), .CK(clk), .Q(ram[2255]) );
  DFF_X1 ram_reg_140__14_ ( .D(n11210), .CK(clk), .Q(ram[2254]) );
  DFF_X1 ram_reg_140__13_ ( .D(n11209), .CK(clk), .Q(ram[2253]) );
  DFF_X1 ram_reg_140__12_ ( .D(n11208), .CK(clk), .Q(ram[2252]) );
  DFF_X1 ram_reg_140__11_ ( .D(n11207), .CK(clk), .Q(ram[2251]) );
  DFF_X1 ram_reg_140__10_ ( .D(n11206), .CK(clk), .Q(ram[2250]) );
  DFF_X1 ram_reg_140__9_ ( .D(n11205), .CK(clk), .Q(ram[2249]) );
  DFF_X1 ram_reg_140__8_ ( .D(n11204), .CK(clk), .Q(ram[2248]) );
  DFF_X1 ram_reg_140__7_ ( .D(n11203), .CK(clk), .Q(ram[2247]) );
  DFF_X1 ram_reg_140__6_ ( .D(n11202), .CK(clk), .Q(ram[2246]) );
  DFF_X1 ram_reg_140__5_ ( .D(n11201), .CK(clk), .Q(ram[2245]) );
  DFF_X1 ram_reg_140__4_ ( .D(n11200), .CK(clk), .Q(ram[2244]) );
  DFF_X1 ram_reg_140__3_ ( .D(n11199), .CK(clk), .Q(ram[2243]) );
  DFF_X1 ram_reg_140__2_ ( .D(n11198), .CK(clk), .Q(ram[2242]) );
  DFF_X1 ram_reg_140__1_ ( .D(n11197), .CK(clk), .Q(ram[2241]) );
  DFF_X1 ram_reg_140__0_ ( .D(n11196), .CK(clk), .Q(ram[2240]) );
  DFF_X1 ram_reg_139__15_ ( .D(n11228), .CK(clk), .Q(ram[2239]) );
  DFF_X1 ram_reg_139__14_ ( .D(n11227), .CK(clk), .Q(ram[2238]) );
  DFF_X1 ram_reg_139__13_ ( .D(n11226), .CK(clk), .Q(ram[2237]) );
  DFF_X1 ram_reg_139__12_ ( .D(n11225), .CK(clk), .Q(ram[2236]) );
  DFF_X1 ram_reg_139__11_ ( .D(n11224), .CK(clk), .Q(ram[2235]) );
  DFF_X1 ram_reg_139__10_ ( .D(n11223), .CK(clk), .Q(ram[2234]) );
  DFF_X1 ram_reg_139__9_ ( .D(n11222), .CK(clk), .Q(ram[2233]) );
  DFF_X1 ram_reg_139__8_ ( .D(n11221), .CK(clk), .Q(ram[2232]) );
  DFF_X1 ram_reg_139__7_ ( .D(n11220), .CK(clk), .Q(ram[2231]) );
  DFF_X1 ram_reg_139__6_ ( .D(n11219), .CK(clk), .Q(ram[2230]) );
  DFF_X1 ram_reg_139__5_ ( .D(n11218), .CK(clk), .Q(ram[2229]) );
  DFF_X1 ram_reg_139__4_ ( .D(n11217), .CK(clk), .Q(ram[2228]) );
  DFF_X1 ram_reg_139__3_ ( .D(n11216), .CK(clk), .Q(ram[2227]) );
  DFF_X1 ram_reg_139__2_ ( .D(n11215), .CK(clk), .Q(ram[2226]) );
  DFF_X1 ram_reg_139__1_ ( .D(n11214), .CK(clk), .Q(ram[2225]) );
  DFF_X1 ram_reg_139__0_ ( .D(n11213), .CK(clk), .Q(ram[2224]) );
  DFF_X1 ram_reg_138__15_ ( .D(n11245), .CK(clk), .Q(ram[2223]) );
  DFF_X1 ram_reg_138__14_ ( .D(n11244), .CK(clk), .Q(ram[2222]) );
  DFF_X1 ram_reg_138__13_ ( .D(n11243), .CK(clk), .Q(ram[2221]) );
  DFF_X1 ram_reg_138__12_ ( .D(n11242), .CK(clk), .Q(ram[2220]) );
  DFF_X1 ram_reg_138__11_ ( .D(n11241), .CK(clk), .Q(ram[2219]) );
  DFF_X1 ram_reg_138__10_ ( .D(n11240), .CK(clk), .Q(ram[2218]) );
  DFF_X1 ram_reg_138__9_ ( .D(n11239), .CK(clk), .Q(ram[2217]) );
  DFF_X1 ram_reg_138__8_ ( .D(n11238), .CK(clk), .Q(ram[2216]) );
  DFF_X1 ram_reg_138__7_ ( .D(n11237), .CK(clk), .Q(ram[2215]) );
  DFF_X1 ram_reg_138__6_ ( .D(n11236), .CK(clk), .Q(ram[2214]) );
  DFF_X1 ram_reg_138__5_ ( .D(n11235), .CK(clk), .Q(ram[2213]) );
  DFF_X1 ram_reg_138__4_ ( .D(n11234), .CK(clk), .Q(ram[2212]) );
  DFF_X1 ram_reg_138__3_ ( .D(n11233), .CK(clk), .Q(ram[2211]) );
  DFF_X1 ram_reg_138__2_ ( .D(n11232), .CK(clk), .Q(ram[2210]) );
  DFF_X1 ram_reg_138__1_ ( .D(n11231), .CK(clk), .Q(ram[2209]) );
  DFF_X1 ram_reg_138__0_ ( .D(n11230), .CK(clk), .Q(ram[2208]) );
  DFF_X1 ram_reg_137__15_ ( .D(n11262), .CK(clk), .Q(ram[2207]) );
  DFF_X1 ram_reg_137__14_ ( .D(n11261), .CK(clk), .Q(ram[2206]) );
  DFF_X1 ram_reg_137__13_ ( .D(n11260), .CK(clk), .Q(ram[2205]) );
  DFF_X1 ram_reg_137__12_ ( .D(n11259), .CK(clk), .Q(ram[2204]) );
  DFF_X1 ram_reg_137__11_ ( .D(n11258), .CK(clk), .Q(ram[2203]) );
  DFF_X1 ram_reg_137__10_ ( .D(n11257), .CK(clk), .Q(ram[2202]) );
  DFF_X1 ram_reg_137__9_ ( .D(n11256), .CK(clk), .Q(ram[2201]) );
  DFF_X1 ram_reg_137__8_ ( .D(n11255), .CK(clk), .Q(ram[2200]) );
  DFF_X1 ram_reg_137__7_ ( .D(n11254), .CK(clk), .Q(ram[2199]) );
  DFF_X1 ram_reg_137__6_ ( .D(n11253), .CK(clk), .Q(ram[2198]) );
  DFF_X1 ram_reg_137__5_ ( .D(n11252), .CK(clk), .Q(ram[2197]) );
  DFF_X1 ram_reg_137__4_ ( .D(n11251), .CK(clk), .Q(ram[2196]) );
  DFF_X1 ram_reg_137__3_ ( .D(n11250), .CK(clk), .Q(ram[2195]) );
  DFF_X1 ram_reg_137__2_ ( .D(n11249), .CK(clk), .Q(ram[2194]) );
  DFF_X1 ram_reg_137__1_ ( .D(n11248), .CK(clk), .Q(ram[2193]) );
  DFF_X1 ram_reg_137__0_ ( .D(n11247), .CK(clk), .Q(ram[2192]) );
  DFF_X1 ram_reg_136__15_ ( .D(n11279), .CK(clk), .Q(ram[2191]) );
  DFF_X1 ram_reg_136__14_ ( .D(n11278), .CK(clk), .Q(ram[2190]) );
  DFF_X1 ram_reg_136__13_ ( .D(n11277), .CK(clk), .Q(ram[2189]) );
  DFF_X1 ram_reg_136__12_ ( .D(n11276), .CK(clk), .Q(ram[2188]) );
  DFF_X1 ram_reg_136__11_ ( .D(n11275), .CK(clk), .Q(ram[2187]) );
  DFF_X1 ram_reg_136__10_ ( .D(n11274), .CK(clk), .Q(ram[2186]) );
  DFF_X1 ram_reg_136__9_ ( .D(n11273), .CK(clk), .Q(ram[2185]) );
  DFF_X1 ram_reg_136__8_ ( .D(n11272), .CK(clk), .Q(ram[2184]) );
  DFF_X1 ram_reg_136__7_ ( .D(n11271), .CK(clk), .Q(ram[2183]) );
  DFF_X1 ram_reg_136__6_ ( .D(n11270), .CK(clk), .Q(ram[2182]) );
  DFF_X1 ram_reg_136__5_ ( .D(n11269), .CK(clk), .Q(ram[2181]) );
  DFF_X1 ram_reg_136__4_ ( .D(n11268), .CK(clk), .Q(ram[2180]) );
  DFF_X1 ram_reg_136__3_ ( .D(n11267), .CK(clk), .Q(ram[2179]) );
  DFF_X1 ram_reg_136__2_ ( .D(n11266), .CK(clk), .Q(ram[2178]) );
  DFF_X1 ram_reg_136__1_ ( .D(n11265), .CK(clk), .Q(ram[2177]) );
  DFF_X1 ram_reg_136__0_ ( .D(n11264), .CK(clk), .Q(ram[2176]) );
  DFF_X1 ram_reg_135__15_ ( .D(n11296), .CK(clk), .Q(ram[2175]) );
  DFF_X1 ram_reg_135__14_ ( .D(n11295), .CK(clk), .Q(ram[2174]) );
  DFF_X1 ram_reg_135__13_ ( .D(n11294), .CK(clk), .Q(ram[2173]) );
  DFF_X1 ram_reg_135__12_ ( .D(n11293), .CK(clk), .Q(ram[2172]) );
  DFF_X1 ram_reg_135__11_ ( .D(n11292), .CK(clk), .Q(ram[2171]) );
  DFF_X1 ram_reg_135__10_ ( .D(n11291), .CK(clk), .Q(ram[2170]) );
  DFF_X1 ram_reg_135__9_ ( .D(n11290), .CK(clk), .Q(ram[2169]) );
  DFF_X1 ram_reg_135__8_ ( .D(n11289), .CK(clk), .Q(ram[2168]) );
  DFF_X1 ram_reg_135__7_ ( .D(n11288), .CK(clk), .Q(ram[2167]) );
  DFF_X1 ram_reg_135__6_ ( .D(n11287), .CK(clk), .Q(ram[2166]) );
  DFF_X1 ram_reg_135__5_ ( .D(n11286), .CK(clk), .Q(ram[2165]) );
  DFF_X1 ram_reg_135__4_ ( .D(n11285), .CK(clk), .Q(ram[2164]) );
  DFF_X1 ram_reg_135__3_ ( .D(n11284), .CK(clk), .Q(ram[2163]) );
  DFF_X1 ram_reg_135__2_ ( .D(n11283), .CK(clk), .Q(ram[2162]) );
  DFF_X1 ram_reg_135__1_ ( .D(n11282), .CK(clk), .Q(ram[2161]) );
  DFF_X1 ram_reg_135__0_ ( .D(n11281), .CK(clk), .Q(ram[2160]) );
  DFF_X1 ram_reg_134__15_ ( .D(n11313), .CK(clk), .Q(ram[2159]) );
  DFF_X1 ram_reg_134__14_ ( .D(n11312), .CK(clk), .Q(ram[2158]) );
  DFF_X1 ram_reg_134__13_ ( .D(n11311), .CK(clk), .Q(ram[2157]) );
  DFF_X1 ram_reg_134__12_ ( .D(n11310), .CK(clk), .Q(ram[2156]) );
  DFF_X1 ram_reg_134__11_ ( .D(n11309), .CK(clk), .Q(ram[2155]) );
  DFF_X1 ram_reg_134__10_ ( .D(n11308), .CK(clk), .Q(ram[2154]) );
  DFF_X1 ram_reg_134__9_ ( .D(n11307), .CK(clk), .Q(ram[2153]) );
  DFF_X1 ram_reg_134__8_ ( .D(n11306), .CK(clk), .Q(ram[2152]) );
  DFF_X1 ram_reg_134__7_ ( .D(n11305), .CK(clk), .Q(ram[2151]) );
  DFF_X1 ram_reg_134__6_ ( .D(n11304), .CK(clk), .Q(ram[2150]) );
  DFF_X1 ram_reg_134__5_ ( .D(n11303), .CK(clk), .Q(ram[2149]) );
  DFF_X1 ram_reg_134__4_ ( .D(n11302), .CK(clk), .Q(ram[2148]) );
  DFF_X1 ram_reg_134__3_ ( .D(n11301), .CK(clk), .Q(ram[2147]) );
  DFF_X1 ram_reg_134__2_ ( .D(n11300), .CK(clk), .Q(ram[2146]) );
  DFF_X1 ram_reg_134__1_ ( .D(n11299), .CK(clk), .Q(ram[2145]) );
  DFF_X1 ram_reg_134__0_ ( .D(n11298), .CK(clk), .Q(ram[2144]) );
  DFF_X1 ram_reg_133__15_ ( .D(n11330), .CK(clk), .Q(ram[2143]) );
  DFF_X1 ram_reg_133__14_ ( .D(n11329), .CK(clk), .Q(ram[2142]) );
  DFF_X1 ram_reg_133__13_ ( .D(n11328), .CK(clk), .Q(ram[2141]) );
  DFF_X1 ram_reg_133__12_ ( .D(n11327), .CK(clk), .Q(ram[2140]) );
  DFF_X1 ram_reg_133__11_ ( .D(n11326), .CK(clk), .Q(ram[2139]) );
  DFF_X1 ram_reg_133__10_ ( .D(n11325), .CK(clk), .Q(ram[2138]) );
  DFF_X1 ram_reg_133__9_ ( .D(n11324), .CK(clk), .Q(ram[2137]) );
  DFF_X1 ram_reg_133__8_ ( .D(n11323), .CK(clk), .Q(ram[2136]) );
  DFF_X1 ram_reg_133__7_ ( .D(n11322), .CK(clk), .Q(ram[2135]) );
  DFF_X1 ram_reg_133__6_ ( .D(n11321), .CK(clk), .Q(ram[2134]) );
  DFF_X1 ram_reg_133__5_ ( .D(n11320), .CK(clk), .Q(ram[2133]) );
  DFF_X1 ram_reg_133__4_ ( .D(n11319), .CK(clk), .Q(ram[2132]) );
  DFF_X1 ram_reg_133__3_ ( .D(n11318), .CK(clk), .Q(ram[2131]) );
  DFF_X1 ram_reg_133__2_ ( .D(n11317), .CK(clk), .Q(ram[2130]) );
  DFF_X1 ram_reg_133__1_ ( .D(n11316), .CK(clk), .Q(ram[2129]) );
  DFF_X1 ram_reg_133__0_ ( .D(n11315), .CK(clk), .Q(ram[2128]) );
  DFF_X1 ram_reg_132__15_ ( .D(n11347), .CK(clk), .Q(ram[2127]) );
  DFF_X1 ram_reg_132__14_ ( .D(n11346), .CK(clk), .Q(ram[2126]) );
  DFF_X1 ram_reg_132__13_ ( .D(n11345), .CK(clk), .Q(ram[2125]) );
  DFF_X1 ram_reg_132__12_ ( .D(n11344), .CK(clk), .Q(ram[2124]) );
  DFF_X1 ram_reg_132__11_ ( .D(n11343), .CK(clk), .Q(ram[2123]) );
  DFF_X1 ram_reg_132__10_ ( .D(n11342), .CK(clk), .Q(ram[2122]) );
  DFF_X1 ram_reg_132__9_ ( .D(n11341), .CK(clk), .Q(ram[2121]) );
  DFF_X1 ram_reg_132__8_ ( .D(n11340), .CK(clk), .Q(ram[2120]) );
  DFF_X1 ram_reg_132__7_ ( .D(n11339), .CK(clk), .Q(ram[2119]) );
  DFF_X1 ram_reg_132__6_ ( .D(n11338), .CK(clk), .Q(ram[2118]) );
  DFF_X1 ram_reg_132__5_ ( .D(n11337), .CK(clk), .Q(ram[2117]) );
  DFF_X1 ram_reg_132__4_ ( .D(n11336), .CK(clk), .Q(ram[2116]) );
  DFF_X1 ram_reg_132__3_ ( .D(n11335), .CK(clk), .Q(ram[2115]) );
  DFF_X1 ram_reg_132__2_ ( .D(n11334), .CK(clk), .Q(ram[2114]) );
  DFF_X1 ram_reg_132__1_ ( .D(n11333), .CK(clk), .Q(ram[2113]) );
  DFF_X1 ram_reg_132__0_ ( .D(n11332), .CK(clk), .Q(ram[2112]) );
  DFF_X1 ram_reg_131__15_ ( .D(n11364), .CK(clk), .Q(ram[2111]) );
  DFF_X1 ram_reg_131__14_ ( .D(n11363), .CK(clk), .Q(ram[2110]) );
  DFF_X1 ram_reg_131__13_ ( .D(n11362), .CK(clk), .Q(ram[2109]) );
  DFF_X1 ram_reg_131__12_ ( .D(n11361), .CK(clk), .Q(ram[2108]) );
  DFF_X1 ram_reg_131__11_ ( .D(n11360), .CK(clk), .Q(ram[2107]) );
  DFF_X1 ram_reg_131__10_ ( .D(n11359), .CK(clk), .Q(ram[2106]) );
  DFF_X1 ram_reg_131__9_ ( .D(n11358), .CK(clk), .Q(ram[2105]) );
  DFF_X1 ram_reg_131__8_ ( .D(n11357), .CK(clk), .Q(ram[2104]) );
  DFF_X1 ram_reg_131__7_ ( .D(n11356), .CK(clk), .Q(ram[2103]) );
  DFF_X1 ram_reg_131__6_ ( .D(n11355), .CK(clk), .Q(ram[2102]) );
  DFF_X1 ram_reg_131__5_ ( .D(n11354), .CK(clk), .Q(ram[2101]) );
  DFF_X1 ram_reg_131__4_ ( .D(n11353), .CK(clk), .Q(ram[2100]) );
  DFF_X1 ram_reg_131__3_ ( .D(n11352), .CK(clk), .Q(ram[2099]) );
  DFF_X1 ram_reg_131__2_ ( .D(n11351), .CK(clk), .Q(ram[2098]) );
  DFF_X1 ram_reg_131__1_ ( .D(n11350), .CK(clk), .Q(ram[2097]) );
  DFF_X1 ram_reg_131__0_ ( .D(n11349), .CK(clk), .Q(ram[2096]) );
  DFF_X1 ram_reg_130__15_ ( .D(n11381), .CK(clk), .Q(ram[2095]) );
  DFF_X1 ram_reg_130__14_ ( .D(n11380), .CK(clk), .Q(ram[2094]) );
  DFF_X1 ram_reg_130__13_ ( .D(n11379), .CK(clk), .Q(ram[2093]) );
  DFF_X1 ram_reg_130__12_ ( .D(n11378), .CK(clk), .Q(ram[2092]) );
  DFF_X1 ram_reg_130__11_ ( .D(n11377), .CK(clk), .Q(ram[2091]) );
  DFF_X1 ram_reg_130__10_ ( .D(n11376), .CK(clk), .Q(ram[2090]) );
  DFF_X1 ram_reg_130__9_ ( .D(n11375), .CK(clk), .Q(ram[2089]) );
  DFF_X1 ram_reg_130__8_ ( .D(n11374), .CK(clk), .Q(ram[2088]) );
  DFF_X1 ram_reg_130__7_ ( .D(n11373), .CK(clk), .Q(ram[2087]) );
  DFF_X1 ram_reg_130__6_ ( .D(n11372), .CK(clk), .Q(ram[2086]) );
  DFF_X1 ram_reg_130__5_ ( .D(n11371), .CK(clk), .Q(ram[2085]) );
  DFF_X1 ram_reg_130__4_ ( .D(n11370), .CK(clk), .Q(ram[2084]) );
  DFF_X1 ram_reg_130__3_ ( .D(n11369), .CK(clk), .Q(ram[2083]) );
  DFF_X1 ram_reg_130__2_ ( .D(n11368), .CK(clk), .Q(ram[2082]) );
  DFF_X1 ram_reg_130__1_ ( .D(n11367), .CK(clk), .Q(ram[2081]) );
  DFF_X1 ram_reg_130__0_ ( .D(n11366), .CK(clk), .Q(ram[2080]) );
  DFF_X1 ram_reg_129__15_ ( .D(n11398), .CK(clk), .Q(ram[2079]) );
  DFF_X1 ram_reg_129__14_ ( .D(n11397), .CK(clk), .Q(ram[2078]) );
  DFF_X1 ram_reg_129__13_ ( .D(n11396), .CK(clk), .Q(ram[2077]) );
  DFF_X1 ram_reg_129__12_ ( .D(n11395), .CK(clk), .Q(ram[2076]) );
  DFF_X1 ram_reg_129__11_ ( .D(n11394), .CK(clk), .Q(ram[2075]) );
  DFF_X1 ram_reg_129__10_ ( .D(n11393), .CK(clk), .Q(ram[2074]) );
  DFF_X1 ram_reg_129__9_ ( .D(n11392), .CK(clk), .Q(ram[2073]) );
  DFF_X1 ram_reg_129__8_ ( .D(n11391), .CK(clk), .Q(ram[2072]) );
  DFF_X1 ram_reg_129__7_ ( .D(n11390), .CK(clk), .Q(ram[2071]) );
  DFF_X1 ram_reg_129__6_ ( .D(n11389), .CK(clk), .Q(ram[2070]) );
  DFF_X1 ram_reg_129__5_ ( .D(n11388), .CK(clk), .Q(ram[2069]) );
  DFF_X1 ram_reg_129__4_ ( .D(n11387), .CK(clk), .Q(ram[2068]) );
  DFF_X1 ram_reg_129__3_ ( .D(n11386), .CK(clk), .Q(ram[2067]) );
  DFF_X1 ram_reg_129__2_ ( .D(n11385), .CK(clk), .Q(ram[2066]) );
  DFF_X1 ram_reg_129__1_ ( .D(n11384), .CK(clk), .Q(ram[2065]) );
  DFF_X1 ram_reg_129__0_ ( .D(n11383), .CK(clk), .Q(ram[2064]) );
  DFF_X1 ram_reg_128__15_ ( .D(n11415), .CK(clk), .Q(ram[2063]) );
  DFF_X1 ram_reg_128__14_ ( .D(n11414), .CK(clk), .Q(ram[2062]) );
  DFF_X1 ram_reg_128__13_ ( .D(n11413), .CK(clk), .Q(ram[2061]) );
  DFF_X1 ram_reg_128__12_ ( .D(n11412), .CK(clk), .Q(ram[2060]) );
  DFF_X1 ram_reg_128__11_ ( .D(n11411), .CK(clk), .Q(ram[2059]) );
  DFF_X1 ram_reg_128__10_ ( .D(n11410), .CK(clk), .Q(ram[2058]) );
  DFF_X1 ram_reg_128__9_ ( .D(n11409), .CK(clk), .Q(ram[2057]) );
  DFF_X1 ram_reg_128__8_ ( .D(n11408), .CK(clk), .Q(ram[2056]) );
  DFF_X1 ram_reg_128__7_ ( .D(n11407), .CK(clk), .Q(ram[2055]) );
  DFF_X1 ram_reg_128__6_ ( .D(n11406), .CK(clk), .Q(ram[2054]) );
  DFF_X1 ram_reg_128__5_ ( .D(n11405), .CK(clk), .Q(ram[2053]) );
  DFF_X1 ram_reg_128__4_ ( .D(n11404), .CK(clk), .Q(ram[2052]) );
  DFF_X1 ram_reg_128__3_ ( .D(n11403), .CK(clk), .Q(ram[2051]) );
  DFF_X1 ram_reg_128__2_ ( .D(n11402), .CK(clk), .Q(ram[2050]) );
  DFF_X1 ram_reg_128__1_ ( .D(n11401), .CK(clk), .Q(ram[2049]) );
  DFF_X1 ram_reg_128__0_ ( .D(n11400), .CK(clk), .Q(ram[2048]) );
  DFF_X1 ram_reg_127__15_ ( .D(n11432), .CK(clk), .Q(ram[2047]) );
  DFF_X1 ram_reg_127__14_ ( .D(n11431), .CK(clk), .Q(ram[2046]) );
  DFF_X1 ram_reg_127__13_ ( .D(n11430), .CK(clk), .Q(ram[2045]) );
  DFF_X1 ram_reg_127__12_ ( .D(n11429), .CK(clk), .Q(ram[2044]) );
  DFF_X1 ram_reg_127__11_ ( .D(n11428), .CK(clk), .Q(ram[2043]) );
  DFF_X1 ram_reg_127__10_ ( .D(n11427), .CK(clk), .Q(ram[2042]) );
  DFF_X1 ram_reg_127__9_ ( .D(n11426), .CK(clk), .Q(ram[2041]) );
  DFF_X1 ram_reg_127__8_ ( .D(n11425), .CK(clk), .Q(ram[2040]) );
  DFF_X1 ram_reg_127__7_ ( .D(n11424), .CK(clk), .Q(ram[2039]) );
  DFF_X1 ram_reg_127__6_ ( .D(n11423), .CK(clk), .Q(ram[2038]) );
  DFF_X1 ram_reg_127__5_ ( .D(n11422), .CK(clk), .Q(ram[2037]) );
  DFF_X1 ram_reg_127__4_ ( .D(n11421), .CK(clk), .Q(ram[2036]) );
  DFF_X1 ram_reg_127__3_ ( .D(n11420), .CK(clk), .Q(ram[2035]) );
  DFF_X1 ram_reg_127__2_ ( .D(n11419), .CK(clk), .Q(ram[2034]) );
  DFF_X1 ram_reg_127__1_ ( .D(n11418), .CK(clk), .Q(ram[2033]) );
  DFF_X1 ram_reg_127__0_ ( .D(n11417), .CK(clk), .Q(ram[2032]) );
  DFF_X1 ram_reg_126__15_ ( .D(n11449), .CK(clk), .Q(ram[2031]) );
  DFF_X1 ram_reg_126__14_ ( .D(n11448), .CK(clk), .Q(ram[2030]) );
  DFF_X1 ram_reg_126__13_ ( .D(n11447), .CK(clk), .Q(ram[2029]) );
  DFF_X1 ram_reg_126__12_ ( .D(n11446), .CK(clk), .Q(ram[2028]) );
  DFF_X1 ram_reg_126__11_ ( .D(n11445), .CK(clk), .Q(ram[2027]) );
  DFF_X1 ram_reg_126__10_ ( .D(n11444), .CK(clk), .Q(ram[2026]) );
  DFF_X1 ram_reg_126__9_ ( .D(n11443), .CK(clk), .Q(ram[2025]) );
  DFF_X1 ram_reg_126__8_ ( .D(n11442), .CK(clk), .Q(ram[2024]) );
  DFF_X1 ram_reg_126__7_ ( .D(n11441), .CK(clk), .Q(ram[2023]) );
  DFF_X1 ram_reg_126__6_ ( .D(n11440), .CK(clk), .Q(ram[2022]) );
  DFF_X1 ram_reg_126__5_ ( .D(n11439), .CK(clk), .Q(ram[2021]) );
  DFF_X1 ram_reg_126__4_ ( .D(n11438), .CK(clk), .Q(ram[2020]) );
  DFF_X1 ram_reg_126__3_ ( .D(n11437), .CK(clk), .Q(ram[2019]) );
  DFF_X1 ram_reg_126__2_ ( .D(n11436), .CK(clk), .Q(ram[2018]) );
  DFF_X1 ram_reg_126__1_ ( .D(n11435), .CK(clk), .Q(ram[2017]) );
  DFF_X1 ram_reg_126__0_ ( .D(n11434), .CK(clk), .Q(ram[2016]) );
  DFF_X1 ram_reg_125__15_ ( .D(n11466), .CK(clk), .Q(ram[2015]) );
  DFF_X1 ram_reg_125__14_ ( .D(n11465), .CK(clk), .Q(ram[2014]) );
  DFF_X1 ram_reg_125__13_ ( .D(n11464), .CK(clk), .Q(ram[2013]) );
  DFF_X1 ram_reg_125__12_ ( .D(n11463), .CK(clk), .Q(ram[2012]) );
  DFF_X1 ram_reg_125__11_ ( .D(n11462), .CK(clk), .Q(ram[2011]) );
  DFF_X1 ram_reg_125__10_ ( .D(n11461), .CK(clk), .Q(ram[2010]) );
  DFF_X1 ram_reg_125__9_ ( .D(n11460), .CK(clk), .Q(ram[2009]) );
  DFF_X1 ram_reg_125__8_ ( .D(n11459), .CK(clk), .Q(ram[2008]) );
  DFF_X1 ram_reg_125__7_ ( .D(n11458), .CK(clk), .Q(ram[2007]) );
  DFF_X1 ram_reg_125__6_ ( .D(n11457), .CK(clk), .Q(ram[2006]) );
  DFF_X1 ram_reg_125__5_ ( .D(n11456), .CK(clk), .Q(ram[2005]) );
  DFF_X1 ram_reg_125__4_ ( .D(n11455), .CK(clk), .Q(ram[2004]) );
  DFF_X1 ram_reg_125__3_ ( .D(n11454), .CK(clk), .Q(ram[2003]) );
  DFF_X1 ram_reg_125__2_ ( .D(n11453), .CK(clk), .Q(ram[2002]) );
  DFF_X1 ram_reg_125__1_ ( .D(n11452), .CK(clk), .Q(ram[2001]) );
  DFF_X1 ram_reg_125__0_ ( .D(n11451), .CK(clk), .Q(ram[2000]) );
  DFF_X1 ram_reg_124__15_ ( .D(n11483), .CK(clk), .Q(ram[1999]) );
  DFF_X1 ram_reg_124__14_ ( .D(n11482), .CK(clk), .Q(ram[1998]) );
  DFF_X1 ram_reg_124__13_ ( .D(n11481), .CK(clk), .Q(ram[1997]) );
  DFF_X1 ram_reg_124__12_ ( .D(n11480), .CK(clk), .Q(ram[1996]) );
  DFF_X1 ram_reg_124__11_ ( .D(n11479), .CK(clk), .Q(ram[1995]) );
  DFF_X1 ram_reg_124__10_ ( .D(n11478), .CK(clk), .Q(ram[1994]) );
  DFF_X1 ram_reg_124__9_ ( .D(n11477), .CK(clk), .Q(ram[1993]) );
  DFF_X1 ram_reg_124__8_ ( .D(n11476), .CK(clk), .Q(ram[1992]) );
  DFF_X1 ram_reg_124__7_ ( .D(n11475), .CK(clk), .Q(ram[1991]) );
  DFF_X1 ram_reg_124__6_ ( .D(n11474), .CK(clk), .Q(ram[1990]) );
  DFF_X1 ram_reg_124__5_ ( .D(n11473), .CK(clk), .Q(ram[1989]) );
  DFF_X1 ram_reg_124__4_ ( .D(n11472), .CK(clk), .Q(ram[1988]) );
  DFF_X1 ram_reg_124__3_ ( .D(n11471), .CK(clk), .Q(ram[1987]) );
  DFF_X1 ram_reg_124__2_ ( .D(n11470), .CK(clk), .Q(ram[1986]) );
  DFF_X1 ram_reg_124__1_ ( .D(n11469), .CK(clk), .Q(ram[1985]) );
  DFF_X1 ram_reg_124__0_ ( .D(n11468), .CK(clk), .Q(ram[1984]) );
  DFF_X1 ram_reg_123__15_ ( .D(n11500), .CK(clk), .Q(ram[1983]) );
  DFF_X1 ram_reg_123__14_ ( .D(n11499), .CK(clk), .Q(ram[1982]) );
  DFF_X1 ram_reg_123__13_ ( .D(n11498), .CK(clk), .Q(ram[1981]) );
  DFF_X1 ram_reg_123__12_ ( .D(n11497), .CK(clk), .Q(ram[1980]) );
  DFF_X1 ram_reg_123__11_ ( .D(n11496), .CK(clk), .Q(ram[1979]) );
  DFF_X1 ram_reg_123__10_ ( .D(n11495), .CK(clk), .Q(ram[1978]) );
  DFF_X1 ram_reg_123__9_ ( .D(n11494), .CK(clk), .Q(ram[1977]) );
  DFF_X1 ram_reg_123__8_ ( .D(n11493), .CK(clk), .Q(ram[1976]) );
  DFF_X1 ram_reg_123__7_ ( .D(n11492), .CK(clk), .Q(ram[1975]) );
  DFF_X1 ram_reg_123__6_ ( .D(n11491), .CK(clk), .Q(ram[1974]) );
  DFF_X1 ram_reg_123__5_ ( .D(n11490), .CK(clk), .Q(ram[1973]) );
  DFF_X1 ram_reg_123__4_ ( .D(n11489), .CK(clk), .Q(ram[1972]) );
  DFF_X1 ram_reg_123__3_ ( .D(n11488), .CK(clk), .Q(ram[1971]) );
  DFF_X1 ram_reg_123__2_ ( .D(n11487), .CK(clk), .Q(ram[1970]) );
  DFF_X1 ram_reg_123__1_ ( .D(n11486), .CK(clk), .Q(ram[1969]) );
  DFF_X1 ram_reg_123__0_ ( .D(n11485), .CK(clk), .Q(ram[1968]) );
  DFF_X1 ram_reg_122__15_ ( .D(n11517), .CK(clk), .Q(ram[1967]) );
  DFF_X1 ram_reg_122__14_ ( .D(n11516), .CK(clk), .Q(ram[1966]) );
  DFF_X1 ram_reg_122__13_ ( .D(n11515), .CK(clk), .Q(ram[1965]) );
  DFF_X1 ram_reg_122__12_ ( .D(n11514), .CK(clk), .Q(ram[1964]) );
  DFF_X1 ram_reg_122__11_ ( .D(n11513), .CK(clk), .Q(ram[1963]) );
  DFF_X1 ram_reg_122__10_ ( .D(n11512), .CK(clk), .Q(ram[1962]) );
  DFF_X1 ram_reg_122__9_ ( .D(n11511), .CK(clk), .Q(ram[1961]) );
  DFF_X1 ram_reg_122__8_ ( .D(n11510), .CK(clk), .Q(ram[1960]) );
  DFF_X1 ram_reg_122__7_ ( .D(n11509), .CK(clk), .Q(ram[1959]) );
  DFF_X1 ram_reg_122__6_ ( .D(n11508), .CK(clk), .Q(ram[1958]) );
  DFF_X1 ram_reg_122__5_ ( .D(n11507), .CK(clk), .Q(ram[1957]) );
  DFF_X1 ram_reg_122__4_ ( .D(n11506), .CK(clk), .Q(ram[1956]) );
  DFF_X1 ram_reg_122__3_ ( .D(n11505), .CK(clk), .Q(ram[1955]) );
  DFF_X1 ram_reg_122__2_ ( .D(n11504), .CK(clk), .Q(ram[1954]) );
  DFF_X1 ram_reg_122__1_ ( .D(n11503), .CK(clk), .Q(ram[1953]) );
  DFF_X1 ram_reg_122__0_ ( .D(n11502), .CK(clk), .Q(ram[1952]) );
  DFF_X1 ram_reg_121__15_ ( .D(n11534), .CK(clk), .Q(ram[1951]) );
  DFF_X1 ram_reg_121__14_ ( .D(n11533), .CK(clk), .Q(ram[1950]) );
  DFF_X1 ram_reg_121__13_ ( .D(n11532), .CK(clk), .Q(ram[1949]) );
  DFF_X1 ram_reg_121__12_ ( .D(n11531), .CK(clk), .Q(ram[1948]) );
  DFF_X1 ram_reg_121__11_ ( .D(n11530), .CK(clk), .Q(ram[1947]) );
  DFF_X1 ram_reg_121__10_ ( .D(n11529), .CK(clk), .Q(ram[1946]) );
  DFF_X1 ram_reg_121__9_ ( .D(n11528), .CK(clk), .Q(ram[1945]) );
  DFF_X1 ram_reg_121__8_ ( .D(n11527), .CK(clk), .Q(ram[1944]) );
  DFF_X1 ram_reg_121__7_ ( .D(n11526), .CK(clk), .Q(ram[1943]) );
  DFF_X1 ram_reg_121__6_ ( .D(n11525), .CK(clk), .Q(ram[1942]) );
  DFF_X1 ram_reg_121__5_ ( .D(n11524), .CK(clk), .Q(ram[1941]) );
  DFF_X1 ram_reg_121__4_ ( .D(n11523), .CK(clk), .Q(ram[1940]) );
  DFF_X1 ram_reg_121__3_ ( .D(n11522), .CK(clk), .Q(ram[1939]) );
  DFF_X1 ram_reg_121__2_ ( .D(n11521), .CK(clk), .Q(ram[1938]) );
  DFF_X1 ram_reg_121__1_ ( .D(n11520), .CK(clk), .Q(ram[1937]) );
  DFF_X1 ram_reg_121__0_ ( .D(n11519), .CK(clk), .Q(ram[1936]) );
  DFF_X1 ram_reg_120__15_ ( .D(n11551), .CK(clk), .Q(ram[1935]) );
  DFF_X1 ram_reg_120__14_ ( .D(n11550), .CK(clk), .Q(ram[1934]) );
  DFF_X1 ram_reg_120__13_ ( .D(n11549), .CK(clk), .Q(ram[1933]) );
  DFF_X1 ram_reg_120__12_ ( .D(n11548), .CK(clk), .Q(ram[1932]) );
  DFF_X1 ram_reg_120__11_ ( .D(n11547), .CK(clk), .Q(ram[1931]) );
  DFF_X1 ram_reg_120__10_ ( .D(n11546), .CK(clk), .Q(ram[1930]) );
  DFF_X1 ram_reg_120__9_ ( .D(n11545), .CK(clk), .Q(ram[1929]) );
  DFF_X1 ram_reg_120__8_ ( .D(n11544), .CK(clk), .Q(ram[1928]) );
  DFF_X1 ram_reg_120__7_ ( .D(n11543), .CK(clk), .Q(ram[1927]) );
  DFF_X1 ram_reg_120__6_ ( .D(n11542), .CK(clk), .Q(ram[1926]) );
  DFF_X1 ram_reg_120__5_ ( .D(n11541), .CK(clk), .Q(ram[1925]) );
  DFF_X1 ram_reg_120__4_ ( .D(n11540), .CK(clk), .Q(ram[1924]) );
  DFF_X1 ram_reg_120__3_ ( .D(n11539), .CK(clk), .Q(ram[1923]) );
  DFF_X1 ram_reg_120__2_ ( .D(n11538), .CK(clk), .Q(ram[1922]) );
  DFF_X1 ram_reg_120__1_ ( .D(n11537), .CK(clk), .Q(ram[1921]) );
  DFF_X1 ram_reg_120__0_ ( .D(n11536), .CK(clk), .Q(ram[1920]) );
  DFF_X1 ram_reg_119__15_ ( .D(n11568), .CK(clk), .Q(ram[1919]) );
  DFF_X1 ram_reg_119__14_ ( .D(n11567), .CK(clk), .Q(ram[1918]) );
  DFF_X1 ram_reg_119__13_ ( .D(n11566), .CK(clk), .Q(ram[1917]) );
  DFF_X1 ram_reg_119__12_ ( .D(n11565), .CK(clk), .Q(ram[1916]) );
  DFF_X1 ram_reg_119__11_ ( .D(n11564), .CK(clk), .Q(ram[1915]) );
  DFF_X1 ram_reg_119__10_ ( .D(n11563), .CK(clk), .Q(ram[1914]) );
  DFF_X1 ram_reg_119__9_ ( .D(n11562), .CK(clk), .Q(ram[1913]) );
  DFF_X1 ram_reg_119__8_ ( .D(n11561), .CK(clk), .Q(ram[1912]) );
  DFF_X1 ram_reg_119__7_ ( .D(n11560), .CK(clk), .Q(ram[1911]) );
  DFF_X1 ram_reg_119__6_ ( .D(n11559), .CK(clk), .Q(ram[1910]) );
  DFF_X1 ram_reg_119__5_ ( .D(n11558), .CK(clk), .Q(ram[1909]) );
  DFF_X1 ram_reg_119__4_ ( .D(n11557), .CK(clk), .Q(ram[1908]) );
  DFF_X1 ram_reg_119__3_ ( .D(n11556), .CK(clk), .Q(ram[1907]) );
  DFF_X1 ram_reg_119__2_ ( .D(n11555), .CK(clk), .Q(ram[1906]) );
  DFF_X1 ram_reg_119__1_ ( .D(n11554), .CK(clk), .Q(ram[1905]) );
  DFF_X1 ram_reg_119__0_ ( .D(n11553), .CK(clk), .Q(ram[1904]) );
  DFF_X1 ram_reg_118__15_ ( .D(n11585), .CK(clk), .Q(ram[1903]) );
  DFF_X1 ram_reg_118__14_ ( .D(n11584), .CK(clk), .Q(ram[1902]) );
  DFF_X1 ram_reg_118__13_ ( .D(n11583), .CK(clk), .Q(ram[1901]) );
  DFF_X1 ram_reg_118__12_ ( .D(n11582), .CK(clk), .Q(ram[1900]) );
  DFF_X1 ram_reg_118__11_ ( .D(n11581), .CK(clk), .Q(ram[1899]) );
  DFF_X1 ram_reg_118__10_ ( .D(n11580), .CK(clk), .Q(ram[1898]) );
  DFF_X1 ram_reg_118__9_ ( .D(n11579), .CK(clk), .Q(ram[1897]) );
  DFF_X1 ram_reg_118__8_ ( .D(n11578), .CK(clk), .Q(ram[1896]) );
  DFF_X1 ram_reg_118__7_ ( .D(n11577), .CK(clk), .Q(ram[1895]) );
  DFF_X1 ram_reg_118__6_ ( .D(n11576), .CK(clk), .Q(ram[1894]) );
  DFF_X1 ram_reg_118__5_ ( .D(n11575), .CK(clk), .Q(ram[1893]) );
  DFF_X1 ram_reg_118__4_ ( .D(n11574), .CK(clk), .Q(ram[1892]) );
  DFF_X1 ram_reg_118__3_ ( .D(n11573), .CK(clk), .Q(ram[1891]) );
  DFF_X1 ram_reg_118__2_ ( .D(n11572), .CK(clk), .Q(ram[1890]) );
  DFF_X1 ram_reg_118__1_ ( .D(n11571), .CK(clk), .Q(ram[1889]) );
  DFF_X1 ram_reg_118__0_ ( .D(n11570), .CK(clk), .Q(ram[1888]) );
  DFF_X1 ram_reg_117__15_ ( .D(n11602), .CK(clk), .Q(ram[1887]) );
  DFF_X1 ram_reg_117__14_ ( .D(n11601), .CK(clk), .Q(ram[1886]) );
  DFF_X1 ram_reg_117__13_ ( .D(n11600), .CK(clk), .Q(ram[1885]) );
  DFF_X1 ram_reg_117__12_ ( .D(n11599), .CK(clk), .Q(ram[1884]) );
  DFF_X1 ram_reg_117__11_ ( .D(n11598), .CK(clk), .Q(ram[1883]) );
  DFF_X1 ram_reg_117__10_ ( .D(n11597), .CK(clk), .Q(ram[1882]) );
  DFF_X1 ram_reg_117__9_ ( .D(n11596), .CK(clk), .Q(ram[1881]) );
  DFF_X1 ram_reg_117__8_ ( .D(n11595), .CK(clk), .Q(ram[1880]) );
  DFF_X1 ram_reg_117__7_ ( .D(n11594), .CK(clk), .Q(ram[1879]) );
  DFF_X1 ram_reg_117__6_ ( .D(n11593), .CK(clk), .Q(ram[1878]) );
  DFF_X1 ram_reg_117__5_ ( .D(n11592), .CK(clk), .Q(ram[1877]) );
  DFF_X1 ram_reg_117__4_ ( .D(n11591), .CK(clk), .Q(ram[1876]) );
  DFF_X1 ram_reg_117__3_ ( .D(n11590), .CK(clk), .Q(ram[1875]) );
  DFF_X1 ram_reg_117__2_ ( .D(n11589), .CK(clk), .Q(ram[1874]) );
  DFF_X1 ram_reg_117__1_ ( .D(n11588), .CK(clk), .Q(ram[1873]) );
  DFF_X1 ram_reg_117__0_ ( .D(n11587), .CK(clk), .Q(ram[1872]) );
  DFF_X1 ram_reg_116__15_ ( .D(n11619), .CK(clk), .Q(ram[1871]) );
  DFF_X1 ram_reg_116__14_ ( .D(n11618), .CK(clk), .Q(ram[1870]) );
  DFF_X1 ram_reg_116__13_ ( .D(n11617), .CK(clk), .Q(ram[1869]) );
  DFF_X1 ram_reg_116__12_ ( .D(n11616), .CK(clk), .Q(ram[1868]) );
  DFF_X1 ram_reg_116__11_ ( .D(n11615), .CK(clk), .Q(ram[1867]) );
  DFF_X1 ram_reg_116__10_ ( .D(n11614), .CK(clk), .Q(ram[1866]) );
  DFF_X1 ram_reg_116__9_ ( .D(n11613), .CK(clk), .Q(ram[1865]) );
  DFF_X1 ram_reg_116__8_ ( .D(n11612), .CK(clk), .Q(ram[1864]) );
  DFF_X1 ram_reg_116__7_ ( .D(n11611), .CK(clk), .Q(ram[1863]) );
  DFF_X1 ram_reg_116__6_ ( .D(n11610), .CK(clk), .Q(ram[1862]) );
  DFF_X1 ram_reg_116__5_ ( .D(n11609), .CK(clk), .Q(ram[1861]) );
  DFF_X1 ram_reg_116__4_ ( .D(n11608), .CK(clk), .Q(ram[1860]) );
  DFF_X1 ram_reg_116__3_ ( .D(n11607), .CK(clk), .Q(ram[1859]) );
  DFF_X1 ram_reg_116__2_ ( .D(n11606), .CK(clk), .Q(ram[1858]) );
  DFF_X1 ram_reg_116__1_ ( .D(n11605), .CK(clk), .Q(ram[1857]) );
  DFF_X1 ram_reg_116__0_ ( .D(n11604), .CK(clk), .Q(ram[1856]) );
  DFF_X1 ram_reg_115__15_ ( .D(n11636), .CK(clk), .Q(ram[1855]) );
  DFF_X1 ram_reg_115__14_ ( .D(n11635), .CK(clk), .Q(ram[1854]) );
  DFF_X1 ram_reg_115__13_ ( .D(n11634), .CK(clk), .Q(ram[1853]) );
  DFF_X1 ram_reg_115__12_ ( .D(n11633), .CK(clk), .Q(ram[1852]) );
  DFF_X1 ram_reg_115__11_ ( .D(n11632), .CK(clk), .Q(ram[1851]) );
  DFF_X1 ram_reg_115__10_ ( .D(n11631), .CK(clk), .Q(ram[1850]) );
  DFF_X1 ram_reg_115__9_ ( .D(n11630), .CK(clk), .Q(ram[1849]) );
  DFF_X1 ram_reg_115__8_ ( .D(n11629), .CK(clk), .Q(ram[1848]) );
  DFF_X1 ram_reg_115__7_ ( .D(n11628), .CK(clk), .Q(ram[1847]) );
  DFF_X1 ram_reg_115__6_ ( .D(n11627), .CK(clk), .Q(ram[1846]) );
  DFF_X1 ram_reg_115__5_ ( .D(n11626), .CK(clk), .Q(ram[1845]) );
  DFF_X1 ram_reg_115__4_ ( .D(n11625), .CK(clk), .Q(ram[1844]) );
  DFF_X1 ram_reg_115__3_ ( .D(n11624), .CK(clk), .Q(ram[1843]) );
  DFF_X1 ram_reg_115__2_ ( .D(n11623), .CK(clk), .Q(ram[1842]) );
  DFF_X1 ram_reg_115__1_ ( .D(n11622), .CK(clk), .Q(ram[1841]) );
  DFF_X1 ram_reg_115__0_ ( .D(n11621), .CK(clk), .Q(ram[1840]) );
  DFF_X1 ram_reg_114__15_ ( .D(n11653), .CK(clk), .Q(ram[1839]) );
  DFF_X1 ram_reg_114__14_ ( .D(n11652), .CK(clk), .Q(ram[1838]) );
  DFF_X1 ram_reg_114__13_ ( .D(n11651), .CK(clk), .Q(ram[1837]) );
  DFF_X1 ram_reg_114__12_ ( .D(n11650), .CK(clk), .Q(ram[1836]) );
  DFF_X1 ram_reg_114__11_ ( .D(n11649), .CK(clk), .Q(ram[1835]) );
  DFF_X1 ram_reg_114__10_ ( .D(n11648), .CK(clk), .Q(ram[1834]) );
  DFF_X1 ram_reg_114__9_ ( .D(n11647), .CK(clk), .Q(ram[1833]) );
  DFF_X1 ram_reg_114__8_ ( .D(n11646), .CK(clk), .Q(ram[1832]) );
  DFF_X1 ram_reg_114__7_ ( .D(n11645), .CK(clk), .Q(ram[1831]) );
  DFF_X1 ram_reg_114__6_ ( .D(n11644), .CK(clk), .Q(ram[1830]) );
  DFF_X1 ram_reg_114__5_ ( .D(n11643), .CK(clk), .Q(ram[1829]) );
  DFF_X1 ram_reg_114__4_ ( .D(n11642), .CK(clk), .Q(ram[1828]) );
  DFF_X1 ram_reg_114__3_ ( .D(n11641), .CK(clk), .Q(ram[1827]) );
  DFF_X1 ram_reg_114__2_ ( .D(n11640), .CK(clk), .Q(ram[1826]) );
  DFF_X1 ram_reg_114__1_ ( .D(n11639), .CK(clk), .Q(ram[1825]) );
  DFF_X1 ram_reg_114__0_ ( .D(n11638), .CK(clk), .Q(ram[1824]) );
  DFF_X1 ram_reg_113__15_ ( .D(n11670), .CK(clk), .Q(ram[1823]) );
  DFF_X1 ram_reg_113__14_ ( .D(n11669), .CK(clk), .Q(ram[1822]) );
  DFF_X1 ram_reg_113__13_ ( .D(n11668), .CK(clk), .Q(ram[1821]) );
  DFF_X1 ram_reg_113__12_ ( .D(n11667), .CK(clk), .Q(ram[1820]) );
  DFF_X1 ram_reg_113__11_ ( .D(n11666), .CK(clk), .Q(ram[1819]) );
  DFF_X1 ram_reg_113__10_ ( .D(n11665), .CK(clk), .Q(ram[1818]) );
  DFF_X1 ram_reg_113__9_ ( .D(n11664), .CK(clk), .Q(ram[1817]) );
  DFF_X1 ram_reg_113__8_ ( .D(n11663), .CK(clk), .Q(ram[1816]) );
  DFF_X1 ram_reg_113__7_ ( .D(n11662), .CK(clk), .Q(ram[1815]) );
  DFF_X1 ram_reg_113__6_ ( .D(n11661), .CK(clk), .Q(ram[1814]) );
  DFF_X1 ram_reg_113__5_ ( .D(n11660), .CK(clk), .Q(ram[1813]) );
  DFF_X1 ram_reg_113__4_ ( .D(n11659), .CK(clk), .Q(ram[1812]) );
  DFF_X1 ram_reg_113__3_ ( .D(n11658), .CK(clk), .Q(ram[1811]) );
  DFF_X1 ram_reg_113__2_ ( .D(n11657), .CK(clk), .Q(ram[1810]) );
  DFF_X1 ram_reg_113__1_ ( .D(n11656), .CK(clk), .Q(ram[1809]) );
  DFF_X1 ram_reg_113__0_ ( .D(n11655), .CK(clk), .Q(ram[1808]) );
  DFF_X1 ram_reg_112__15_ ( .D(n11687), .CK(clk), .Q(ram[1807]) );
  DFF_X1 ram_reg_112__14_ ( .D(n11686), .CK(clk), .Q(ram[1806]) );
  DFF_X1 ram_reg_112__13_ ( .D(n11685), .CK(clk), .Q(ram[1805]) );
  DFF_X1 ram_reg_112__12_ ( .D(n11684), .CK(clk), .Q(ram[1804]) );
  DFF_X1 ram_reg_112__11_ ( .D(n11683), .CK(clk), .Q(ram[1803]) );
  DFF_X1 ram_reg_112__10_ ( .D(n11682), .CK(clk), .Q(ram[1802]) );
  DFF_X1 ram_reg_112__9_ ( .D(n11681), .CK(clk), .Q(ram[1801]) );
  DFF_X1 ram_reg_112__8_ ( .D(n11680), .CK(clk), .Q(ram[1800]) );
  DFF_X1 ram_reg_112__7_ ( .D(n11679), .CK(clk), .Q(ram[1799]) );
  DFF_X1 ram_reg_112__6_ ( .D(n11678), .CK(clk), .Q(ram[1798]) );
  DFF_X1 ram_reg_112__5_ ( .D(n11677), .CK(clk), .Q(ram[1797]) );
  DFF_X1 ram_reg_112__4_ ( .D(n11676), .CK(clk), .Q(ram[1796]) );
  DFF_X1 ram_reg_112__3_ ( .D(n11675), .CK(clk), .Q(ram[1795]) );
  DFF_X1 ram_reg_112__2_ ( .D(n11674), .CK(clk), .Q(ram[1794]) );
  DFF_X1 ram_reg_112__1_ ( .D(n11673), .CK(clk), .Q(ram[1793]) );
  DFF_X1 ram_reg_112__0_ ( .D(n11672), .CK(clk), .Q(ram[1792]) );
  DFF_X1 ram_reg_111__15_ ( .D(n11704), .CK(clk), .Q(ram[1791]) );
  DFF_X1 ram_reg_111__14_ ( .D(n11703), .CK(clk), .Q(ram[1790]) );
  DFF_X1 ram_reg_111__13_ ( .D(n11702), .CK(clk), .Q(ram[1789]) );
  DFF_X1 ram_reg_111__12_ ( .D(n11701), .CK(clk), .Q(ram[1788]) );
  DFF_X1 ram_reg_111__11_ ( .D(n11700), .CK(clk), .Q(ram[1787]) );
  DFF_X1 ram_reg_111__10_ ( .D(n11699), .CK(clk), .Q(ram[1786]) );
  DFF_X1 ram_reg_111__9_ ( .D(n11698), .CK(clk), .Q(ram[1785]) );
  DFF_X1 ram_reg_111__8_ ( .D(n11697), .CK(clk), .Q(ram[1784]) );
  DFF_X1 ram_reg_111__7_ ( .D(n11696), .CK(clk), .Q(ram[1783]) );
  DFF_X1 ram_reg_111__6_ ( .D(n11695), .CK(clk), .Q(ram[1782]) );
  DFF_X1 ram_reg_111__5_ ( .D(n11694), .CK(clk), .Q(ram[1781]) );
  DFF_X1 ram_reg_111__4_ ( .D(n11693), .CK(clk), .Q(ram[1780]) );
  DFF_X1 ram_reg_111__3_ ( .D(n11692), .CK(clk), .Q(ram[1779]) );
  DFF_X1 ram_reg_111__2_ ( .D(n11691), .CK(clk), .Q(ram[1778]) );
  DFF_X1 ram_reg_111__1_ ( .D(n11690), .CK(clk), .Q(ram[1777]) );
  DFF_X1 ram_reg_111__0_ ( .D(n11689), .CK(clk), .Q(ram[1776]) );
  DFF_X1 ram_reg_110__15_ ( .D(n11721), .CK(clk), .Q(ram[1775]) );
  DFF_X1 ram_reg_110__14_ ( .D(n11720), .CK(clk), .Q(ram[1774]) );
  DFF_X1 ram_reg_110__13_ ( .D(n11719), .CK(clk), .Q(ram[1773]) );
  DFF_X1 ram_reg_110__12_ ( .D(n11718), .CK(clk), .Q(ram[1772]) );
  DFF_X1 ram_reg_110__11_ ( .D(n11717), .CK(clk), .Q(ram[1771]) );
  DFF_X1 ram_reg_110__10_ ( .D(n11716), .CK(clk), .Q(ram[1770]) );
  DFF_X1 ram_reg_110__9_ ( .D(n11715), .CK(clk), .Q(ram[1769]) );
  DFF_X1 ram_reg_110__8_ ( .D(n11714), .CK(clk), .Q(ram[1768]) );
  DFF_X1 ram_reg_110__7_ ( .D(n11713), .CK(clk), .Q(ram[1767]) );
  DFF_X1 ram_reg_110__6_ ( .D(n11712), .CK(clk), .Q(ram[1766]) );
  DFF_X1 ram_reg_110__5_ ( .D(n11711), .CK(clk), .Q(ram[1765]) );
  DFF_X1 ram_reg_110__4_ ( .D(n11710), .CK(clk), .Q(ram[1764]) );
  DFF_X1 ram_reg_110__3_ ( .D(n11709), .CK(clk), .Q(ram[1763]) );
  DFF_X1 ram_reg_110__2_ ( .D(n11708), .CK(clk), .Q(ram[1762]) );
  DFF_X1 ram_reg_110__1_ ( .D(n11707), .CK(clk), .Q(ram[1761]) );
  DFF_X1 ram_reg_110__0_ ( .D(n11706), .CK(clk), .Q(ram[1760]) );
  DFF_X1 ram_reg_109__15_ ( .D(n11738), .CK(clk), .Q(ram[1759]) );
  DFF_X1 ram_reg_109__14_ ( .D(n11737), .CK(clk), .Q(ram[1758]) );
  DFF_X1 ram_reg_109__13_ ( .D(n11736), .CK(clk), .Q(ram[1757]) );
  DFF_X1 ram_reg_109__12_ ( .D(n11735), .CK(clk), .Q(ram[1756]) );
  DFF_X1 ram_reg_109__11_ ( .D(n11734), .CK(clk), .Q(ram[1755]) );
  DFF_X1 ram_reg_109__10_ ( .D(n11733), .CK(clk), .Q(ram[1754]) );
  DFF_X1 ram_reg_109__9_ ( .D(n11732), .CK(clk), .Q(ram[1753]) );
  DFF_X1 ram_reg_109__8_ ( .D(n11731), .CK(clk), .Q(ram[1752]) );
  DFF_X1 ram_reg_109__7_ ( .D(n11730), .CK(clk), .Q(ram[1751]) );
  DFF_X1 ram_reg_109__6_ ( .D(n11729), .CK(clk), .Q(ram[1750]) );
  DFF_X1 ram_reg_109__5_ ( .D(n11728), .CK(clk), .Q(ram[1749]) );
  DFF_X1 ram_reg_109__4_ ( .D(n11727), .CK(clk), .Q(ram[1748]) );
  DFF_X1 ram_reg_109__3_ ( .D(n11726), .CK(clk), .Q(ram[1747]) );
  DFF_X1 ram_reg_109__2_ ( .D(n11725), .CK(clk), .Q(ram[1746]) );
  DFF_X1 ram_reg_109__1_ ( .D(n11724), .CK(clk), .Q(ram[1745]) );
  DFF_X1 ram_reg_109__0_ ( .D(n11723), .CK(clk), .Q(ram[1744]) );
  DFF_X1 ram_reg_108__15_ ( .D(n11755), .CK(clk), .Q(ram[1743]) );
  DFF_X1 ram_reg_108__14_ ( .D(n11754), .CK(clk), .Q(ram[1742]) );
  DFF_X1 ram_reg_108__13_ ( .D(n11753), .CK(clk), .Q(ram[1741]) );
  DFF_X1 ram_reg_108__12_ ( .D(n11752), .CK(clk), .Q(ram[1740]) );
  DFF_X1 ram_reg_108__11_ ( .D(n11751), .CK(clk), .Q(ram[1739]) );
  DFF_X1 ram_reg_108__10_ ( .D(n11750), .CK(clk), .Q(ram[1738]) );
  DFF_X1 ram_reg_108__9_ ( .D(n11749), .CK(clk), .Q(ram[1737]) );
  DFF_X1 ram_reg_108__8_ ( .D(n11748), .CK(clk), .Q(ram[1736]) );
  DFF_X1 ram_reg_108__7_ ( .D(n11747), .CK(clk), .Q(ram[1735]) );
  DFF_X1 ram_reg_108__6_ ( .D(n11746), .CK(clk), .Q(ram[1734]) );
  DFF_X1 ram_reg_108__5_ ( .D(n11745), .CK(clk), .Q(ram[1733]) );
  DFF_X1 ram_reg_108__4_ ( .D(n11744), .CK(clk), .Q(ram[1732]) );
  DFF_X1 ram_reg_108__3_ ( .D(n11743), .CK(clk), .Q(ram[1731]) );
  DFF_X1 ram_reg_108__2_ ( .D(n11742), .CK(clk), .Q(ram[1730]) );
  DFF_X1 ram_reg_108__1_ ( .D(n11741), .CK(clk), .Q(ram[1729]) );
  DFF_X1 ram_reg_108__0_ ( .D(n11740), .CK(clk), .Q(ram[1728]) );
  DFF_X1 ram_reg_107__15_ ( .D(n11772), .CK(clk), .Q(ram[1727]) );
  DFF_X1 ram_reg_107__14_ ( .D(n11771), .CK(clk), .Q(ram[1726]) );
  DFF_X1 ram_reg_107__13_ ( .D(n11770), .CK(clk), .Q(ram[1725]) );
  DFF_X1 ram_reg_107__12_ ( .D(n11769), .CK(clk), .Q(ram[1724]) );
  DFF_X1 ram_reg_107__11_ ( .D(n11768), .CK(clk), .Q(ram[1723]) );
  DFF_X1 ram_reg_107__10_ ( .D(n11767), .CK(clk), .Q(ram[1722]) );
  DFF_X1 ram_reg_107__9_ ( .D(n11766), .CK(clk), .Q(ram[1721]) );
  DFF_X1 ram_reg_107__8_ ( .D(n11765), .CK(clk), .Q(ram[1720]) );
  DFF_X1 ram_reg_107__7_ ( .D(n11764), .CK(clk), .Q(ram[1719]) );
  DFF_X1 ram_reg_107__6_ ( .D(n11763), .CK(clk), .Q(ram[1718]) );
  DFF_X1 ram_reg_107__5_ ( .D(n11762), .CK(clk), .Q(ram[1717]) );
  DFF_X1 ram_reg_107__4_ ( .D(n11761), .CK(clk), .Q(ram[1716]) );
  DFF_X1 ram_reg_107__3_ ( .D(n11760), .CK(clk), .Q(ram[1715]) );
  DFF_X1 ram_reg_107__2_ ( .D(n11759), .CK(clk), .Q(ram[1714]) );
  DFF_X1 ram_reg_107__1_ ( .D(n11758), .CK(clk), .Q(ram[1713]) );
  DFF_X1 ram_reg_107__0_ ( .D(n11757), .CK(clk), .Q(ram[1712]) );
  DFF_X1 ram_reg_106__15_ ( .D(n11789), .CK(clk), .Q(ram[1711]) );
  DFF_X1 ram_reg_106__14_ ( .D(n11788), .CK(clk), .Q(ram[1710]) );
  DFF_X1 ram_reg_106__13_ ( .D(n11787), .CK(clk), .Q(ram[1709]) );
  DFF_X1 ram_reg_106__12_ ( .D(n11786), .CK(clk), .Q(ram[1708]) );
  DFF_X1 ram_reg_106__11_ ( .D(n11785), .CK(clk), .Q(ram[1707]) );
  DFF_X1 ram_reg_106__10_ ( .D(n11784), .CK(clk), .Q(ram[1706]) );
  DFF_X1 ram_reg_106__9_ ( .D(n11783), .CK(clk), .Q(ram[1705]) );
  DFF_X1 ram_reg_106__8_ ( .D(n11782), .CK(clk), .Q(ram[1704]) );
  DFF_X1 ram_reg_106__7_ ( .D(n11781), .CK(clk), .Q(ram[1703]) );
  DFF_X1 ram_reg_106__6_ ( .D(n11780), .CK(clk), .Q(ram[1702]) );
  DFF_X1 ram_reg_106__5_ ( .D(n11779), .CK(clk), .Q(ram[1701]) );
  DFF_X1 ram_reg_106__4_ ( .D(n11778), .CK(clk), .Q(ram[1700]) );
  DFF_X1 ram_reg_106__3_ ( .D(n11777), .CK(clk), .Q(ram[1699]) );
  DFF_X1 ram_reg_106__2_ ( .D(n11776), .CK(clk), .Q(ram[1698]) );
  DFF_X1 ram_reg_106__1_ ( .D(n11775), .CK(clk), .Q(ram[1697]) );
  DFF_X1 ram_reg_106__0_ ( .D(n11774), .CK(clk), .Q(ram[1696]) );
  DFF_X1 ram_reg_105__15_ ( .D(n11806), .CK(clk), .Q(ram[1695]) );
  DFF_X1 ram_reg_105__14_ ( .D(n11805), .CK(clk), .Q(ram[1694]) );
  DFF_X1 ram_reg_105__13_ ( .D(n11804), .CK(clk), .Q(ram[1693]) );
  DFF_X1 ram_reg_105__12_ ( .D(n11803), .CK(clk), .Q(ram[1692]) );
  DFF_X1 ram_reg_105__11_ ( .D(n11802), .CK(clk), .Q(ram[1691]) );
  DFF_X1 ram_reg_105__10_ ( .D(n11801), .CK(clk), .Q(ram[1690]) );
  DFF_X1 ram_reg_105__9_ ( .D(n11800), .CK(clk), .Q(ram[1689]) );
  DFF_X1 ram_reg_105__8_ ( .D(n11799), .CK(clk), .Q(ram[1688]) );
  DFF_X1 ram_reg_105__7_ ( .D(n11798), .CK(clk), .Q(ram[1687]) );
  DFF_X1 ram_reg_105__6_ ( .D(n11797), .CK(clk), .Q(ram[1686]) );
  DFF_X1 ram_reg_105__5_ ( .D(n11796), .CK(clk), .Q(ram[1685]) );
  DFF_X1 ram_reg_105__4_ ( .D(n11795), .CK(clk), .Q(ram[1684]) );
  DFF_X1 ram_reg_105__3_ ( .D(n11794), .CK(clk), .Q(ram[1683]) );
  DFF_X1 ram_reg_105__2_ ( .D(n11793), .CK(clk), .Q(ram[1682]) );
  DFF_X1 ram_reg_105__1_ ( .D(n11792), .CK(clk), .Q(ram[1681]) );
  DFF_X1 ram_reg_105__0_ ( .D(n11791), .CK(clk), .Q(ram[1680]) );
  DFF_X1 ram_reg_104__15_ ( .D(n11823), .CK(clk), .Q(ram[1679]) );
  DFF_X1 ram_reg_104__14_ ( .D(n11822), .CK(clk), .Q(ram[1678]) );
  DFF_X1 ram_reg_104__13_ ( .D(n11821), .CK(clk), .Q(ram[1677]) );
  DFF_X1 ram_reg_104__12_ ( .D(n11820), .CK(clk), .Q(ram[1676]) );
  DFF_X1 ram_reg_104__11_ ( .D(n11819), .CK(clk), .Q(ram[1675]) );
  DFF_X1 ram_reg_104__10_ ( .D(n11818), .CK(clk), .Q(ram[1674]) );
  DFF_X1 ram_reg_104__9_ ( .D(n11817), .CK(clk), .Q(ram[1673]) );
  DFF_X1 ram_reg_104__8_ ( .D(n11816), .CK(clk), .Q(ram[1672]) );
  DFF_X1 ram_reg_104__7_ ( .D(n11815), .CK(clk), .Q(ram[1671]) );
  DFF_X1 ram_reg_104__6_ ( .D(n11814), .CK(clk), .Q(ram[1670]) );
  DFF_X1 ram_reg_104__5_ ( .D(n11813), .CK(clk), .Q(ram[1669]) );
  DFF_X1 ram_reg_104__4_ ( .D(n11812), .CK(clk), .Q(ram[1668]) );
  DFF_X1 ram_reg_104__3_ ( .D(n11811), .CK(clk), .Q(ram[1667]) );
  DFF_X1 ram_reg_104__2_ ( .D(n11810), .CK(clk), .Q(ram[1666]) );
  DFF_X1 ram_reg_104__1_ ( .D(n11809), .CK(clk), .Q(ram[1665]) );
  DFF_X1 ram_reg_104__0_ ( .D(n11808), .CK(clk), .Q(ram[1664]) );
  DFF_X1 ram_reg_103__15_ ( .D(n11840), .CK(clk), .Q(ram[1663]) );
  DFF_X1 ram_reg_103__14_ ( .D(n11839), .CK(clk), .Q(ram[1662]) );
  DFF_X1 ram_reg_103__13_ ( .D(n11838), .CK(clk), .Q(ram[1661]) );
  DFF_X1 ram_reg_103__12_ ( .D(n11837), .CK(clk), .Q(ram[1660]) );
  DFF_X1 ram_reg_103__11_ ( .D(n11836), .CK(clk), .Q(ram[1659]) );
  DFF_X1 ram_reg_103__10_ ( .D(n11835), .CK(clk), .Q(ram[1658]) );
  DFF_X1 ram_reg_103__9_ ( .D(n11834), .CK(clk), .Q(ram[1657]) );
  DFF_X1 ram_reg_103__8_ ( .D(n11833), .CK(clk), .Q(ram[1656]) );
  DFF_X1 ram_reg_103__7_ ( .D(n11832), .CK(clk), .Q(ram[1655]) );
  DFF_X1 ram_reg_103__6_ ( .D(n11831), .CK(clk), .Q(ram[1654]) );
  DFF_X1 ram_reg_103__5_ ( .D(n11830), .CK(clk), .Q(ram[1653]) );
  DFF_X1 ram_reg_103__4_ ( .D(n11829), .CK(clk), .Q(ram[1652]) );
  DFF_X1 ram_reg_103__3_ ( .D(n11828), .CK(clk), .Q(ram[1651]) );
  DFF_X1 ram_reg_103__2_ ( .D(n11827), .CK(clk), .Q(ram[1650]) );
  DFF_X1 ram_reg_103__1_ ( .D(n11826), .CK(clk), .Q(ram[1649]) );
  DFF_X1 ram_reg_103__0_ ( .D(n11825), .CK(clk), .Q(ram[1648]) );
  DFF_X1 ram_reg_102__15_ ( .D(n11857), .CK(clk), .Q(ram[1647]) );
  DFF_X1 ram_reg_102__14_ ( .D(n11856), .CK(clk), .Q(ram[1646]) );
  DFF_X1 ram_reg_102__13_ ( .D(n11855), .CK(clk), .Q(ram[1645]) );
  DFF_X1 ram_reg_102__12_ ( .D(n11854), .CK(clk), .Q(ram[1644]) );
  DFF_X1 ram_reg_102__11_ ( .D(n11853), .CK(clk), .Q(ram[1643]) );
  DFF_X1 ram_reg_102__10_ ( .D(n11852), .CK(clk), .Q(ram[1642]) );
  DFF_X1 ram_reg_102__9_ ( .D(n11851), .CK(clk), .Q(ram[1641]) );
  DFF_X1 ram_reg_102__8_ ( .D(n11850), .CK(clk), .Q(ram[1640]) );
  DFF_X1 ram_reg_102__7_ ( .D(n11849), .CK(clk), .Q(ram[1639]) );
  DFF_X1 ram_reg_102__6_ ( .D(n11848), .CK(clk), .Q(ram[1638]) );
  DFF_X1 ram_reg_102__5_ ( .D(n11847), .CK(clk), .Q(ram[1637]) );
  DFF_X1 ram_reg_102__4_ ( .D(n11846), .CK(clk), .Q(ram[1636]) );
  DFF_X1 ram_reg_102__3_ ( .D(n11845), .CK(clk), .Q(ram[1635]) );
  DFF_X1 ram_reg_102__2_ ( .D(n11844), .CK(clk), .Q(ram[1634]) );
  DFF_X1 ram_reg_102__1_ ( .D(n11843), .CK(clk), .Q(ram[1633]) );
  DFF_X1 ram_reg_102__0_ ( .D(n11842), .CK(clk), .Q(ram[1632]) );
  DFF_X1 ram_reg_101__15_ ( .D(n11874), .CK(clk), .Q(ram[1631]) );
  DFF_X1 ram_reg_101__14_ ( .D(n11873), .CK(clk), .Q(ram[1630]) );
  DFF_X1 ram_reg_101__13_ ( .D(n11872), .CK(clk), .Q(ram[1629]) );
  DFF_X1 ram_reg_101__12_ ( .D(n11871), .CK(clk), .Q(ram[1628]) );
  DFF_X1 ram_reg_101__11_ ( .D(n11870), .CK(clk), .Q(ram[1627]) );
  DFF_X1 ram_reg_101__10_ ( .D(n11869), .CK(clk), .Q(ram[1626]) );
  DFF_X1 ram_reg_101__9_ ( .D(n11868), .CK(clk), .Q(ram[1625]) );
  DFF_X1 ram_reg_101__8_ ( .D(n11867), .CK(clk), .Q(ram[1624]) );
  DFF_X1 ram_reg_101__7_ ( .D(n11866), .CK(clk), .Q(ram[1623]) );
  DFF_X1 ram_reg_101__6_ ( .D(n11865), .CK(clk), .Q(ram[1622]) );
  DFF_X1 ram_reg_101__5_ ( .D(n11864), .CK(clk), .Q(ram[1621]) );
  DFF_X1 ram_reg_101__4_ ( .D(n11863), .CK(clk), .Q(ram[1620]) );
  DFF_X1 ram_reg_101__3_ ( .D(n11862), .CK(clk), .Q(ram[1619]) );
  DFF_X1 ram_reg_101__2_ ( .D(n11861), .CK(clk), .Q(ram[1618]) );
  DFF_X1 ram_reg_101__1_ ( .D(n11860), .CK(clk), .Q(ram[1617]) );
  DFF_X1 ram_reg_101__0_ ( .D(n11859), .CK(clk), .Q(ram[1616]) );
  DFF_X1 ram_reg_100__15_ ( .D(n11891), .CK(clk), .Q(ram[1615]) );
  DFF_X1 ram_reg_100__14_ ( .D(n11890), .CK(clk), .Q(ram[1614]) );
  DFF_X1 ram_reg_100__13_ ( .D(n11889), .CK(clk), .Q(ram[1613]) );
  DFF_X1 ram_reg_100__12_ ( .D(n11888), .CK(clk), .Q(ram[1612]) );
  DFF_X1 ram_reg_100__11_ ( .D(n11887), .CK(clk), .Q(ram[1611]) );
  DFF_X1 ram_reg_100__10_ ( .D(n11886), .CK(clk), .Q(ram[1610]) );
  DFF_X1 ram_reg_100__9_ ( .D(n11885), .CK(clk), .Q(ram[1609]) );
  DFF_X1 ram_reg_100__8_ ( .D(n11884), .CK(clk), .Q(ram[1608]) );
  DFF_X1 ram_reg_100__7_ ( .D(n11883), .CK(clk), .Q(ram[1607]) );
  DFF_X1 ram_reg_100__6_ ( .D(n11882), .CK(clk), .Q(ram[1606]) );
  DFF_X1 ram_reg_100__5_ ( .D(n11881), .CK(clk), .Q(ram[1605]) );
  DFF_X1 ram_reg_100__4_ ( .D(n11880), .CK(clk), .Q(ram[1604]) );
  DFF_X1 ram_reg_100__3_ ( .D(n11879), .CK(clk), .Q(ram[1603]) );
  DFF_X1 ram_reg_100__2_ ( .D(n11878), .CK(clk), .Q(ram[1602]) );
  DFF_X1 ram_reg_100__1_ ( .D(n11877), .CK(clk), .Q(ram[1601]) );
  DFF_X1 ram_reg_100__0_ ( .D(n11876), .CK(clk), .Q(ram[1600]) );
  DFF_X1 ram_reg_99__15_ ( .D(n11908), .CK(clk), .Q(ram[1599]) );
  DFF_X1 ram_reg_99__14_ ( .D(n11907), .CK(clk), .Q(ram[1598]) );
  DFF_X1 ram_reg_99__13_ ( .D(n11906), .CK(clk), .Q(ram[1597]) );
  DFF_X1 ram_reg_99__12_ ( .D(n11905), .CK(clk), .Q(ram[1596]) );
  DFF_X1 ram_reg_99__11_ ( .D(n11904), .CK(clk), .Q(ram[1595]) );
  DFF_X1 ram_reg_99__10_ ( .D(n11903), .CK(clk), .Q(ram[1594]) );
  DFF_X1 ram_reg_99__9_ ( .D(n11902), .CK(clk), .Q(ram[1593]) );
  DFF_X1 ram_reg_99__8_ ( .D(n11901), .CK(clk), .Q(ram[1592]) );
  DFF_X1 ram_reg_99__7_ ( .D(n11900), .CK(clk), .Q(ram[1591]) );
  DFF_X1 ram_reg_99__6_ ( .D(n11899), .CK(clk), .Q(ram[1590]) );
  DFF_X1 ram_reg_99__5_ ( .D(n11898), .CK(clk), .Q(ram[1589]) );
  DFF_X1 ram_reg_99__4_ ( .D(n11897), .CK(clk), .Q(ram[1588]) );
  DFF_X1 ram_reg_99__3_ ( .D(n11896), .CK(clk), .Q(ram[1587]) );
  DFF_X1 ram_reg_99__2_ ( .D(n11895), .CK(clk), .Q(ram[1586]) );
  DFF_X1 ram_reg_99__1_ ( .D(n11894), .CK(clk), .Q(ram[1585]) );
  DFF_X1 ram_reg_99__0_ ( .D(n11893), .CK(clk), .Q(ram[1584]) );
  DFF_X1 ram_reg_98__15_ ( .D(n11925), .CK(clk), .Q(ram[1583]) );
  DFF_X1 ram_reg_98__14_ ( .D(n11924), .CK(clk), .Q(ram[1582]) );
  DFF_X1 ram_reg_98__13_ ( .D(n11923), .CK(clk), .Q(ram[1581]) );
  DFF_X1 ram_reg_98__12_ ( .D(n11922), .CK(clk), .Q(ram[1580]) );
  DFF_X1 ram_reg_98__11_ ( .D(n11921), .CK(clk), .Q(ram[1579]) );
  DFF_X1 ram_reg_98__10_ ( .D(n11920), .CK(clk), .Q(ram[1578]) );
  DFF_X1 ram_reg_98__9_ ( .D(n11919), .CK(clk), .Q(ram[1577]) );
  DFF_X1 ram_reg_98__8_ ( .D(n11918), .CK(clk), .Q(ram[1576]) );
  DFF_X1 ram_reg_98__7_ ( .D(n11917), .CK(clk), .Q(ram[1575]) );
  DFF_X1 ram_reg_98__6_ ( .D(n11916), .CK(clk), .Q(ram[1574]) );
  DFF_X1 ram_reg_98__5_ ( .D(n11915), .CK(clk), .Q(ram[1573]) );
  DFF_X1 ram_reg_98__4_ ( .D(n11914), .CK(clk), .Q(ram[1572]) );
  DFF_X1 ram_reg_98__3_ ( .D(n11913), .CK(clk), .Q(ram[1571]) );
  DFF_X1 ram_reg_98__2_ ( .D(n11912), .CK(clk), .Q(ram[1570]) );
  DFF_X1 ram_reg_98__1_ ( .D(n11911), .CK(clk), .Q(ram[1569]) );
  DFF_X1 ram_reg_98__0_ ( .D(n11910), .CK(clk), .Q(ram[1568]) );
  DFF_X1 ram_reg_97__15_ ( .D(n11942), .CK(clk), .Q(ram[1567]) );
  DFF_X1 ram_reg_97__14_ ( .D(n11941), .CK(clk), .Q(ram[1566]) );
  DFF_X1 ram_reg_97__13_ ( .D(n11940), .CK(clk), .Q(ram[1565]) );
  DFF_X1 ram_reg_97__12_ ( .D(n11939), .CK(clk), .Q(ram[1564]) );
  DFF_X1 ram_reg_97__11_ ( .D(n11938), .CK(clk), .Q(ram[1563]) );
  DFF_X1 ram_reg_97__10_ ( .D(n11937), .CK(clk), .Q(ram[1562]) );
  DFF_X1 ram_reg_97__9_ ( .D(n11936), .CK(clk), .Q(ram[1561]) );
  DFF_X1 ram_reg_97__8_ ( .D(n11935), .CK(clk), .Q(ram[1560]) );
  DFF_X1 ram_reg_97__7_ ( .D(n11934), .CK(clk), .Q(ram[1559]) );
  DFF_X1 ram_reg_97__6_ ( .D(n11933), .CK(clk), .Q(ram[1558]) );
  DFF_X1 ram_reg_97__5_ ( .D(n11932), .CK(clk), .Q(ram[1557]) );
  DFF_X1 ram_reg_97__4_ ( .D(n11931), .CK(clk), .Q(ram[1556]) );
  DFF_X1 ram_reg_97__3_ ( .D(n11930), .CK(clk), .Q(ram[1555]) );
  DFF_X1 ram_reg_97__2_ ( .D(n11929), .CK(clk), .Q(ram[1554]) );
  DFF_X1 ram_reg_97__1_ ( .D(n11928), .CK(clk), .Q(ram[1553]) );
  DFF_X1 ram_reg_97__0_ ( .D(n11927), .CK(clk), .Q(ram[1552]) );
  DFF_X1 ram_reg_96__15_ ( .D(n11959), .CK(clk), .Q(ram[1551]) );
  DFF_X1 ram_reg_96__14_ ( .D(n11958), .CK(clk), .Q(ram[1550]) );
  DFF_X1 ram_reg_96__13_ ( .D(n11957), .CK(clk), .Q(ram[1549]) );
  DFF_X1 ram_reg_96__12_ ( .D(n11956), .CK(clk), .Q(ram[1548]) );
  DFF_X1 ram_reg_96__11_ ( .D(n11955), .CK(clk), .Q(ram[1547]) );
  DFF_X1 ram_reg_96__10_ ( .D(n11954), .CK(clk), .Q(ram[1546]) );
  DFF_X1 ram_reg_96__9_ ( .D(n11953), .CK(clk), .Q(ram[1545]) );
  DFF_X1 ram_reg_96__8_ ( .D(n11952), .CK(clk), .Q(ram[1544]) );
  DFF_X1 ram_reg_96__7_ ( .D(n11951), .CK(clk), .Q(ram[1543]) );
  DFF_X1 ram_reg_96__6_ ( .D(n11950), .CK(clk), .Q(ram[1542]) );
  DFF_X1 ram_reg_96__5_ ( .D(n11949), .CK(clk), .Q(ram[1541]) );
  DFF_X1 ram_reg_96__4_ ( .D(n11948), .CK(clk), .Q(ram[1540]) );
  DFF_X1 ram_reg_96__3_ ( .D(n11947), .CK(clk), .Q(ram[1539]) );
  DFF_X1 ram_reg_96__2_ ( .D(n11946), .CK(clk), .Q(ram[1538]) );
  DFF_X1 ram_reg_96__1_ ( .D(n11945), .CK(clk), .Q(ram[1537]) );
  DFF_X1 ram_reg_96__0_ ( .D(n11944), .CK(clk), .Q(ram[1536]) );
  DFF_X1 ram_reg_95__15_ ( .D(n11976), .CK(clk), .Q(ram[1535]) );
  DFF_X1 ram_reg_95__14_ ( .D(n11975), .CK(clk), .Q(ram[1534]) );
  DFF_X1 ram_reg_95__13_ ( .D(n11974), .CK(clk), .Q(ram[1533]) );
  DFF_X1 ram_reg_95__12_ ( .D(n11973), .CK(clk), .Q(ram[1532]) );
  DFF_X1 ram_reg_95__11_ ( .D(n11972), .CK(clk), .Q(ram[1531]) );
  DFF_X1 ram_reg_95__10_ ( .D(n11971), .CK(clk), .Q(ram[1530]) );
  DFF_X1 ram_reg_95__9_ ( .D(n11970), .CK(clk), .Q(ram[1529]) );
  DFF_X1 ram_reg_95__8_ ( .D(n11969), .CK(clk), .Q(ram[1528]) );
  DFF_X1 ram_reg_95__7_ ( .D(n11968), .CK(clk), .Q(ram[1527]) );
  DFF_X1 ram_reg_95__6_ ( .D(n11967), .CK(clk), .Q(ram[1526]) );
  DFF_X1 ram_reg_95__5_ ( .D(n11966), .CK(clk), .Q(ram[1525]) );
  DFF_X1 ram_reg_95__4_ ( .D(n11965), .CK(clk), .Q(ram[1524]) );
  DFF_X1 ram_reg_95__3_ ( .D(n11964), .CK(clk), .Q(ram[1523]) );
  DFF_X1 ram_reg_95__2_ ( .D(n11963), .CK(clk), .Q(ram[1522]) );
  DFF_X1 ram_reg_95__1_ ( .D(n11962), .CK(clk), .Q(ram[1521]) );
  DFF_X1 ram_reg_95__0_ ( .D(n11961), .CK(clk), .Q(ram[1520]) );
  DFF_X1 ram_reg_94__15_ ( .D(n11993), .CK(clk), .Q(ram[1519]) );
  DFF_X1 ram_reg_94__14_ ( .D(n11992), .CK(clk), .Q(ram[1518]) );
  DFF_X1 ram_reg_94__13_ ( .D(n11991), .CK(clk), .Q(ram[1517]) );
  DFF_X1 ram_reg_94__12_ ( .D(n11990), .CK(clk), .Q(ram[1516]) );
  DFF_X1 ram_reg_94__11_ ( .D(n11989), .CK(clk), .Q(ram[1515]) );
  DFF_X1 ram_reg_94__10_ ( .D(n11988), .CK(clk), .Q(ram[1514]) );
  DFF_X1 ram_reg_94__9_ ( .D(n11987), .CK(clk), .Q(ram[1513]) );
  DFF_X1 ram_reg_94__8_ ( .D(n11986), .CK(clk), .Q(ram[1512]) );
  DFF_X1 ram_reg_94__7_ ( .D(n11985), .CK(clk), .Q(ram[1511]) );
  DFF_X1 ram_reg_94__6_ ( .D(n11984), .CK(clk), .Q(ram[1510]) );
  DFF_X1 ram_reg_94__5_ ( .D(n11983), .CK(clk), .Q(ram[1509]) );
  DFF_X1 ram_reg_94__4_ ( .D(n11982), .CK(clk), .Q(ram[1508]) );
  DFF_X1 ram_reg_94__3_ ( .D(n11981), .CK(clk), .Q(ram[1507]) );
  DFF_X1 ram_reg_94__2_ ( .D(n11980), .CK(clk), .Q(ram[1506]) );
  DFF_X1 ram_reg_94__1_ ( .D(n11979), .CK(clk), .Q(ram[1505]) );
  DFF_X1 ram_reg_94__0_ ( .D(n11978), .CK(clk), .Q(ram[1504]) );
  DFF_X1 ram_reg_93__15_ ( .D(n12010), .CK(clk), .Q(ram[1503]) );
  DFF_X1 ram_reg_93__14_ ( .D(n12009), .CK(clk), .Q(ram[1502]) );
  DFF_X1 ram_reg_93__13_ ( .D(n12008), .CK(clk), .Q(ram[1501]) );
  DFF_X1 ram_reg_93__12_ ( .D(n12007), .CK(clk), .Q(ram[1500]) );
  DFF_X1 ram_reg_93__11_ ( .D(n12006), .CK(clk), .Q(ram[1499]) );
  DFF_X1 ram_reg_93__10_ ( .D(n12005), .CK(clk), .Q(ram[1498]) );
  DFF_X1 ram_reg_93__9_ ( .D(n12004), .CK(clk), .Q(ram[1497]) );
  DFF_X1 ram_reg_93__8_ ( .D(n12003), .CK(clk), .Q(ram[1496]) );
  DFF_X1 ram_reg_93__7_ ( .D(n12002), .CK(clk), .Q(ram[1495]) );
  DFF_X1 ram_reg_93__6_ ( .D(n12001), .CK(clk), .Q(ram[1494]) );
  DFF_X1 ram_reg_93__5_ ( .D(n12000), .CK(clk), .Q(ram[1493]) );
  DFF_X1 ram_reg_93__4_ ( .D(n11999), .CK(clk), .Q(ram[1492]) );
  DFF_X1 ram_reg_93__3_ ( .D(n11998), .CK(clk), .Q(ram[1491]) );
  DFF_X1 ram_reg_93__2_ ( .D(n11997), .CK(clk), .Q(ram[1490]) );
  DFF_X1 ram_reg_93__1_ ( .D(n11996), .CK(clk), .Q(ram[1489]) );
  DFF_X1 ram_reg_93__0_ ( .D(n11995), .CK(clk), .Q(ram[1488]) );
  DFF_X1 ram_reg_92__15_ ( .D(n12027), .CK(clk), .Q(ram[1487]) );
  DFF_X1 ram_reg_92__14_ ( .D(n12026), .CK(clk), .Q(ram[1486]) );
  DFF_X1 ram_reg_92__13_ ( .D(n12025), .CK(clk), .Q(ram[1485]) );
  DFF_X1 ram_reg_92__12_ ( .D(n12024), .CK(clk), .Q(ram[1484]) );
  DFF_X1 ram_reg_92__11_ ( .D(n12023), .CK(clk), .Q(ram[1483]) );
  DFF_X1 ram_reg_92__10_ ( .D(n12022), .CK(clk), .Q(ram[1482]) );
  DFF_X1 ram_reg_92__9_ ( .D(n12021), .CK(clk), .Q(ram[1481]) );
  DFF_X1 ram_reg_92__8_ ( .D(n12020), .CK(clk), .Q(ram[1480]) );
  DFF_X1 ram_reg_92__7_ ( .D(n12019), .CK(clk), .Q(ram[1479]) );
  DFF_X1 ram_reg_92__6_ ( .D(n12018), .CK(clk), .Q(ram[1478]) );
  DFF_X1 ram_reg_92__5_ ( .D(n12017), .CK(clk), .Q(ram[1477]) );
  DFF_X1 ram_reg_92__4_ ( .D(n12016), .CK(clk), .Q(ram[1476]) );
  DFF_X1 ram_reg_92__3_ ( .D(n12015), .CK(clk), .Q(ram[1475]) );
  DFF_X1 ram_reg_92__2_ ( .D(n12014), .CK(clk), .Q(ram[1474]) );
  DFF_X1 ram_reg_92__1_ ( .D(n12013), .CK(clk), .Q(ram[1473]) );
  DFF_X1 ram_reg_92__0_ ( .D(n12012), .CK(clk), .Q(ram[1472]) );
  DFF_X1 ram_reg_91__15_ ( .D(n12044), .CK(clk), .Q(ram[1471]) );
  DFF_X1 ram_reg_91__14_ ( .D(n12043), .CK(clk), .Q(ram[1470]) );
  DFF_X1 ram_reg_91__13_ ( .D(n12042), .CK(clk), .Q(ram[1469]) );
  DFF_X1 ram_reg_91__12_ ( .D(n12041), .CK(clk), .Q(ram[1468]) );
  DFF_X1 ram_reg_91__11_ ( .D(n12040), .CK(clk), .Q(ram[1467]) );
  DFF_X1 ram_reg_91__10_ ( .D(n12039), .CK(clk), .Q(ram[1466]) );
  DFF_X1 ram_reg_91__9_ ( .D(n12038), .CK(clk), .Q(ram[1465]) );
  DFF_X1 ram_reg_91__8_ ( .D(n12037), .CK(clk), .Q(ram[1464]) );
  DFF_X1 ram_reg_91__7_ ( .D(n12036), .CK(clk), .Q(ram[1463]) );
  DFF_X1 ram_reg_91__6_ ( .D(n12035), .CK(clk), .Q(ram[1462]) );
  DFF_X1 ram_reg_91__5_ ( .D(n12034), .CK(clk), .Q(ram[1461]) );
  DFF_X1 ram_reg_91__4_ ( .D(n12033), .CK(clk), .Q(ram[1460]) );
  DFF_X1 ram_reg_91__3_ ( .D(n12032), .CK(clk), .Q(ram[1459]) );
  DFF_X1 ram_reg_91__2_ ( .D(n12031), .CK(clk), .Q(ram[1458]) );
  DFF_X1 ram_reg_91__1_ ( .D(n12030), .CK(clk), .Q(ram[1457]) );
  DFF_X1 ram_reg_91__0_ ( .D(n12029), .CK(clk), .Q(ram[1456]) );
  DFF_X1 ram_reg_90__15_ ( .D(n12061), .CK(clk), .Q(ram[1455]) );
  DFF_X1 ram_reg_90__14_ ( .D(n12060), .CK(clk), .Q(ram[1454]) );
  DFF_X1 ram_reg_90__13_ ( .D(n12059), .CK(clk), .Q(ram[1453]) );
  DFF_X1 ram_reg_90__12_ ( .D(n12058), .CK(clk), .Q(ram[1452]) );
  DFF_X1 ram_reg_90__11_ ( .D(n12057), .CK(clk), .Q(ram[1451]) );
  DFF_X1 ram_reg_90__10_ ( .D(n12056), .CK(clk), .Q(ram[1450]) );
  DFF_X1 ram_reg_90__9_ ( .D(n12055), .CK(clk), .Q(ram[1449]) );
  DFF_X1 ram_reg_90__8_ ( .D(n12054), .CK(clk), .Q(ram[1448]) );
  DFF_X1 ram_reg_90__7_ ( .D(n12053), .CK(clk), .Q(ram[1447]) );
  DFF_X1 ram_reg_90__6_ ( .D(n12052), .CK(clk), .Q(ram[1446]) );
  DFF_X1 ram_reg_90__5_ ( .D(n12051), .CK(clk), .Q(ram[1445]) );
  DFF_X1 ram_reg_90__4_ ( .D(n12050), .CK(clk), .Q(ram[1444]) );
  DFF_X1 ram_reg_90__3_ ( .D(n12049), .CK(clk), .Q(ram[1443]) );
  DFF_X1 ram_reg_90__2_ ( .D(n12048), .CK(clk), .Q(ram[1442]) );
  DFF_X1 ram_reg_90__1_ ( .D(n12047), .CK(clk), .Q(ram[1441]) );
  DFF_X1 ram_reg_90__0_ ( .D(n12046), .CK(clk), .Q(ram[1440]) );
  DFF_X1 ram_reg_89__15_ ( .D(n12078), .CK(clk), .Q(ram[1439]) );
  DFF_X1 ram_reg_89__14_ ( .D(n12077), .CK(clk), .Q(ram[1438]) );
  DFF_X1 ram_reg_89__13_ ( .D(n12076), .CK(clk), .Q(ram[1437]) );
  DFF_X1 ram_reg_89__12_ ( .D(n12075), .CK(clk), .Q(ram[1436]) );
  DFF_X1 ram_reg_89__11_ ( .D(n12074), .CK(clk), .Q(ram[1435]) );
  DFF_X1 ram_reg_89__10_ ( .D(n12073), .CK(clk), .Q(ram[1434]) );
  DFF_X1 ram_reg_89__9_ ( .D(n12072), .CK(clk), .Q(ram[1433]) );
  DFF_X1 ram_reg_89__8_ ( .D(n12071), .CK(clk), .Q(ram[1432]) );
  DFF_X1 ram_reg_89__7_ ( .D(n12070), .CK(clk), .Q(ram[1431]) );
  DFF_X1 ram_reg_89__6_ ( .D(n12069), .CK(clk), .Q(ram[1430]) );
  DFF_X1 ram_reg_89__5_ ( .D(n12068), .CK(clk), .Q(ram[1429]) );
  DFF_X1 ram_reg_89__4_ ( .D(n12067), .CK(clk), .Q(ram[1428]) );
  DFF_X1 ram_reg_89__3_ ( .D(n12066), .CK(clk), .Q(ram[1427]) );
  DFF_X1 ram_reg_89__2_ ( .D(n12065), .CK(clk), .Q(ram[1426]) );
  DFF_X1 ram_reg_89__1_ ( .D(n12064), .CK(clk), .Q(ram[1425]) );
  DFF_X1 ram_reg_89__0_ ( .D(n12063), .CK(clk), .Q(ram[1424]) );
  DFF_X1 ram_reg_88__15_ ( .D(n12095), .CK(clk), .Q(ram[1423]) );
  DFF_X1 ram_reg_88__14_ ( .D(n12094), .CK(clk), .Q(ram[1422]) );
  DFF_X1 ram_reg_88__13_ ( .D(n12093), .CK(clk), .Q(ram[1421]) );
  DFF_X1 ram_reg_88__12_ ( .D(n12092), .CK(clk), .Q(ram[1420]) );
  DFF_X1 ram_reg_88__11_ ( .D(n12091), .CK(clk), .Q(ram[1419]) );
  DFF_X1 ram_reg_88__10_ ( .D(n12090), .CK(clk), .Q(ram[1418]) );
  DFF_X1 ram_reg_88__9_ ( .D(n12089), .CK(clk), .Q(ram[1417]) );
  DFF_X1 ram_reg_88__8_ ( .D(n12088), .CK(clk), .Q(ram[1416]) );
  DFF_X1 ram_reg_88__7_ ( .D(n12087), .CK(clk), .Q(ram[1415]) );
  DFF_X1 ram_reg_88__6_ ( .D(n12086), .CK(clk), .Q(ram[1414]) );
  DFF_X1 ram_reg_88__5_ ( .D(n12085), .CK(clk), .Q(ram[1413]) );
  DFF_X1 ram_reg_88__4_ ( .D(n12084), .CK(clk), .Q(ram[1412]) );
  DFF_X1 ram_reg_88__3_ ( .D(n12083), .CK(clk), .Q(ram[1411]) );
  DFF_X1 ram_reg_88__2_ ( .D(n12082), .CK(clk), .Q(ram[1410]) );
  DFF_X1 ram_reg_88__1_ ( .D(n12081), .CK(clk), .Q(ram[1409]) );
  DFF_X1 ram_reg_88__0_ ( .D(n12080), .CK(clk), .Q(ram[1408]) );
  DFF_X1 ram_reg_87__15_ ( .D(n12112), .CK(clk), .Q(ram[1407]) );
  DFF_X1 ram_reg_87__14_ ( .D(n12111), .CK(clk), .Q(ram[1406]) );
  DFF_X1 ram_reg_87__13_ ( .D(n12110), .CK(clk), .Q(ram[1405]) );
  DFF_X1 ram_reg_87__12_ ( .D(n12109), .CK(clk), .Q(ram[1404]) );
  DFF_X1 ram_reg_87__11_ ( .D(n12108), .CK(clk), .Q(ram[1403]) );
  DFF_X1 ram_reg_87__10_ ( .D(n12107), .CK(clk), .Q(ram[1402]) );
  DFF_X1 ram_reg_87__9_ ( .D(n12106), .CK(clk), .Q(ram[1401]) );
  DFF_X1 ram_reg_87__8_ ( .D(n12105), .CK(clk), .Q(ram[1400]) );
  DFF_X1 ram_reg_87__7_ ( .D(n12104), .CK(clk), .Q(ram[1399]) );
  DFF_X1 ram_reg_87__6_ ( .D(n12103), .CK(clk), .Q(ram[1398]) );
  DFF_X1 ram_reg_87__5_ ( .D(n12102), .CK(clk), .Q(ram[1397]) );
  DFF_X1 ram_reg_87__4_ ( .D(n12101), .CK(clk), .Q(ram[1396]) );
  DFF_X1 ram_reg_87__3_ ( .D(n12100), .CK(clk), .Q(ram[1395]) );
  DFF_X1 ram_reg_87__2_ ( .D(n12099), .CK(clk), .Q(ram[1394]) );
  DFF_X1 ram_reg_87__1_ ( .D(n12098), .CK(clk), .Q(ram[1393]) );
  DFF_X1 ram_reg_87__0_ ( .D(n12097), .CK(clk), .Q(ram[1392]) );
  DFF_X1 ram_reg_86__15_ ( .D(n12129), .CK(clk), .Q(ram[1391]) );
  DFF_X1 ram_reg_86__14_ ( .D(n12128), .CK(clk), .Q(ram[1390]) );
  DFF_X1 ram_reg_86__13_ ( .D(n12127), .CK(clk), .Q(ram[1389]) );
  DFF_X1 ram_reg_86__12_ ( .D(n12126), .CK(clk), .Q(ram[1388]) );
  DFF_X1 ram_reg_86__11_ ( .D(n12125), .CK(clk), .Q(ram[1387]) );
  DFF_X1 ram_reg_86__10_ ( .D(n12124), .CK(clk), .Q(ram[1386]) );
  DFF_X1 ram_reg_86__9_ ( .D(n12123), .CK(clk), .Q(ram[1385]) );
  DFF_X1 ram_reg_86__8_ ( .D(n12122), .CK(clk), .Q(ram[1384]) );
  DFF_X1 ram_reg_86__7_ ( .D(n12121), .CK(clk), .Q(ram[1383]) );
  DFF_X1 ram_reg_86__6_ ( .D(n12120), .CK(clk), .Q(ram[1382]) );
  DFF_X1 ram_reg_86__5_ ( .D(n12119), .CK(clk), .Q(ram[1381]) );
  DFF_X1 ram_reg_86__4_ ( .D(n12118), .CK(clk), .Q(ram[1380]) );
  DFF_X1 ram_reg_86__3_ ( .D(n12117), .CK(clk), .Q(ram[1379]) );
  DFF_X1 ram_reg_86__2_ ( .D(n12116), .CK(clk), .Q(ram[1378]) );
  DFF_X1 ram_reg_86__1_ ( .D(n12115), .CK(clk), .Q(ram[1377]) );
  DFF_X1 ram_reg_86__0_ ( .D(n12114), .CK(clk), .Q(ram[1376]) );
  DFF_X1 ram_reg_85__15_ ( .D(n12146), .CK(clk), .Q(ram[1375]) );
  DFF_X1 ram_reg_85__14_ ( .D(n12145), .CK(clk), .Q(ram[1374]) );
  DFF_X1 ram_reg_85__13_ ( .D(n12144), .CK(clk), .Q(ram[1373]) );
  DFF_X1 ram_reg_85__12_ ( .D(n12143), .CK(clk), .Q(ram[1372]) );
  DFF_X1 ram_reg_85__11_ ( .D(n12142), .CK(clk), .Q(ram[1371]) );
  DFF_X1 ram_reg_85__10_ ( .D(n12141), .CK(clk), .Q(ram[1370]) );
  DFF_X1 ram_reg_85__9_ ( .D(n12140), .CK(clk), .Q(ram[1369]) );
  DFF_X1 ram_reg_85__8_ ( .D(n12139), .CK(clk), .Q(ram[1368]) );
  DFF_X1 ram_reg_85__7_ ( .D(n12138), .CK(clk), .Q(ram[1367]) );
  DFF_X1 ram_reg_85__6_ ( .D(n12137), .CK(clk), .Q(ram[1366]) );
  DFF_X1 ram_reg_85__5_ ( .D(n12136), .CK(clk), .Q(ram[1365]) );
  DFF_X1 ram_reg_85__4_ ( .D(n12135), .CK(clk), .Q(ram[1364]) );
  DFF_X1 ram_reg_85__3_ ( .D(n12134), .CK(clk), .Q(ram[1363]) );
  DFF_X1 ram_reg_85__2_ ( .D(n12133), .CK(clk), .Q(ram[1362]) );
  DFF_X1 ram_reg_85__1_ ( .D(n12132), .CK(clk), .Q(ram[1361]) );
  DFF_X1 ram_reg_85__0_ ( .D(n12131), .CK(clk), .Q(ram[1360]) );
  DFF_X1 ram_reg_84__15_ ( .D(n12163), .CK(clk), .Q(ram[1359]) );
  DFF_X1 ram_reg_84__14_ ( .D(n12162), .CK(clk), .Q(ram[1358]) );
  DFF_X1 ram_reg_84__13_ ( .D(n12161), .CK(clk), .Q(ram[1357]) );
  DFF_X1 ram_reg_84__12_ ( .D(n12160), .CK(clk), .Q(ram[1356]) );
  DFF_X1 ram_reg_84__11_ ( .D(n12159), .CK(clk), .Q(ram[1355]) );
  DFF_X1 ram_reg_84__10_ ( .D(n12158), .CK(clk), .Q(ram[1354]) );
  DFF_X1 ram_reg_84__9_ ( .D(n12157), .CK(clk), .Q(ram[1353]) );
  DFF_X1 ram_reg_84__8_ ( .D(n12156), .CK(clk), .Q(ram[1352]) );
  DFF_X1 ram_reg_84__7_ ( .D(n12155), .CK(clk), .Q(ram[1351]) );
  DFF_X1 ram_reg_84__6_ ( .D(n12154), .CK(clk), .Q(ram[1350]) );
  DFF_X1 ram_reg_84__5_ ( .D(n12153), .CK(clk), .Q(ram[1349]) );
  DFF_X1 ram_reg_84__4_ ( .D(n12152), .CK(clk), .Q(ram[1348]) );
  DFF_X1 ram_reg_84__3_ ( .D(n12151), .CK(clk), .Q(ram[1347]) );
  DFF_X1 ram_reg_84__2_ ( .D(n12150), .CK(clk), .Q(ram[1346]) );
  DFF_X1 ram_reg_84__1_ ( .D(n12149), .CK(clk), .Q(ram[1345]) );
  DFF_X1 ram_reg_84__0_ ( .D(n12148), .CK(clk), .Q(ram[1344]) );
  DFF_X1 ram_reg_83__15_ ( .D(n12180), .CK(clk), .Q(ram[1343]) );
  DFF_X1 ram_reg_83__14_ ( .D(n12179), .CK(clk), .Q(ram[1342]) );
  DFF_X1 ram_reg_83__13_ ( .D(n12178), .CK(clk), .Q(ram[1341]) );
  DFF_X1 ram_reg_83__12_ ( .D(n12177), .CK(clk), .Q(ram[1340]) );
  DFF_X1 ram_reg_83__11_ ( .D(n12176), .CK(clk), .Q(ram[1339]) );
  DFF_X1 ram_reg_83__10_ ( .D(n12175), .CK(clk), .Q(ram[1338]) );
  DFF_X1 ram_reg_83__9_ ( .D(n12174), .CK(clk), .Q(ram[1337]) );
  DFF_X1 ram_reg_83__8_ ( .D(n12173), .CK(clk), .Q(ram[1336]) );
  DFF_X1 ram_reg_83__7_ ( .D(n12172), .CK(clk), .Q(ram[1335]) );
  DFF_X1 ram_reg_83__6_ ( .D(n12171), .CK(clk), .Q(ram[1334]) );
  DFF_X1 ram_reg_83__5_ ( .D(n12170), .CK(clk), .Q(ram[1333]) );
  DFF_X1 ram_reg_83__4_ ( .D(n12169), .CK(clk), .Q(ram[1332]) );
  DFF_X1 ram_reg_83__3_ ( .D(n12168), .CK(clk), .Q(ram[1331]) );
  DFF_X1 ram_reg_83__2_ ( .D(n12167), .CK(clk), .Q(ram[1330]) );
  DFF_X1 ram_reg_83__1_ ( .D(n12166), .CK(clk), .Q(ram[1329]) );
  DFF_X1 ram_reg_83__0_ ( .D(n12165), .CK(clk), .Q(ram[1328]) );
  DFF_X1 ram_reg_82__15_ ( .D(n12197), .CK(clk), .Q(ram[1327]) );
  DFF_X1 ram_reg_82__14_ ( .D(n12196), .CK(clk), .Q(ram[1326]) );
  DFF_X1 ram_reg_82__13_ ( .D(n12195), .CK(clk), .Q(ram[1325]) );
  DFF_X1 ram_reg_82__12_ ( .D(n12194), .CK(clk), .Q(ram[1324]) );
  DFF_X1 ram_reg_82__11_ ( .D(n12193), .CK(clk), .Q(ram[1323]) );
  DFF_X1 ram_reg_82__10_ ( .D(n12192), .CK(clk), .Q(ram[1322]) );
  DFF_X1 ram_reg_82__9_ ( .D(n12191), .CK(clk), .Q(ram[1321]) );
  DFF_X1 ram_reg_82__8_ ( .D(n12190), .CK(clk), .Q(ram[1320]) );
  DFF_X1 ram_reg_82__7_ ( .D(n12189), .CK(clk), .Q(ram[1319]) );
  DFF_X1 ram_reg_82__6_ ( .D(n12188), .CK(clk), .Q(ram[1318]) );
  DFF_X1 ram_reg_82__5_ ( .D(n12187), .CK(clk), .Q(ram[1317]) );
  DFF_X1 ram_reg_82__4_ ( .D(n12186), .CK(clk), .Q(ram[1316]) );
  DFF_X1 ram_reg_82__3_ ( .D(n12185), .CK(clk), .Q(ram[1315]) );
  DFF_X1 ram_reg_82__2_ ( .D(n12184), .CK(clk), .Q(ram[1314]) );
  DFF_X1 ram_reg_82__1_ ( .D(n12183), .CK(clk), .Q(ram[1313]) );
  DFF_X1 ram_reg_82__0_ ( .D(n12182), .CK(clk), .Q(ram[1312]) );
  DFF_X1 ram_reg_81__15_ ( .D(n12214), .CK(clk), .Q(ram[1311]) );
  DFF_X1 ram_reg_81__14_ ( .D(n12213), .CK(clk), .Q(ram[1310]) );
  DFF_X1 ram_reg_81__13_ ( .D(n12212), .CK(clk), .Q(ram[1309]) );
  DFF_X1 ram_reg_81__12_ ( .D(n12211), .CK(clk), .Q(ram[1308]) );
  DFF_X1 ram_reg_81__11_ ( .D(n12210), .CK(clk), .Q(ram[1307]) );
  DFF_X1 ram_reg_81__10_ ( .D(n12209), .CK(clk), .Q(ram[1306]) );
  DFF_X1 ram_reg_81__9_ ( .D(n12208), .CK(clk), .Q(ram[1305]) );
  DFF_X1 ram_reg_81__8_ ( .D(n12207), .CK(clk), .Q(ram[1304]) );
  DFF_X1 ram_reg_81__7_ ( .D(n12206), .CK(clk), .Q(ram[1303]) );
  DFF_X1 ram_reg_81__6_ ( .D(n12205), .CK(clk), .Q(ram[1302]) );
  DFF_X1 ram_reg_81__5_ ( .D(n12204), .CK(clk), .Q(ram[1301]) );
  DFF_X1 ram_reg_81__4_ ( .D(n12203), .CK(clk), .Q(ram[1300]) );
  DFF_X1 ram_reg_81__3_ ( .D(n12202), .CK(clk), .Q(ram[1299]) );
  DFF_X1 ram_reg_81__2_ ( .D(n12201), .CK(clk), .Q(ram[1298]) );
  DFF_X1 ram_reg_81__1_ ( .D(n12200), .CK(clk), .Q(ram[1297]) );
  DFF_X1 ram_reg_81__0_ ( .D(n12199), .CK(clk), .Q(ram[1296]) );
  DFF_X1 ram_reg_80__15_ ( .D(n12231), .CK(clk), .Q(ram[1295]) );
  DFF_X1 ram_reg_80__14_ ( .D(n12230), .CK(clk), .Q(ram[1294]) );
  DFF_X1 ram_reg_80__13_ ( .D(n12229), .CK(clk), .Q(ram[1293]) );
  DFF_X1 ram_reg_80__12_ ( .D(n12228), .CK(clk), .Q(ram[1292]) );
  DFF_X1 ram_reg_80__11_ ( .D(n12227), .CK(clk), .Q(ram[1291]) );
  DFF_X1 ram_reg_80__10_ ( .D(n12226), .CK(clk), .Q(ram[1290]) );
  DFF_X1 ram_reg_80__9_ ( .D(n12225), .CK(clk), .Q(ram[1289]) );
  DFF_X1 ram_reg_80__8_ ( .D(n12224), .CK(clk), .Q(ram[1288]) );
  DFF_X1 ram_reg_80__7_ ( .D(n12223), .CK(clk), .Q(ram[1287]) );
  DFF_X1 ram_reg_80__6_ ( .D(n12222), .CK(clk), .Q(ram[1286]) );
  DFF_X1 ram_reg_80__5_ ( .D(n12221), .CK(clk), .Q(ram[1285]) );
  DFF_X1 ram_reg_80__4_ ( .D(n12220), .CK(clk), .Q(ram[1284]) );
  DFF_X1 ram_reg_80__3_ ( .D(n12219), .CK(clk), .Q(ram[1283]) );
  DFF_X1 ram_reg_80__2_ ( .D(n12218), .CK(clk), .Q(ram[1282]) );
  DFF_X1 ram_reg_80__1_ ( .D(n12217), .CK(clk), .Q(ram[1281]) );
  DFF_X1 ram_reg_80__0_ ( .D(n12216), .CK(clk), .Q(ram[1280]) );
  DFF_X1 ram_reg_79__15_ ( .D(n12248), .CK(clk), .Q(ram[1279]) );
  DFF_X1 ram_reg_79__14_ ( .D(n12247), .CK(clk), .Q(ram[1278]) );
  DFF_X1 ram_reg_79__13_ ( .D(n12246), .CK(clk), .Q(ram[1277]) );
  DFF_X1 ram_reg_79__12_ ( .D(n12245), .CK(clk), .Q(ram[1276]) );
  DFF_X1 ram_reg_79__11_ ( .D(n12244), .CK(clk), .Q(ram[1275]) );
  DFF_X1 ram_reg_79__10_ ( .D(n12243), .CK(clk), .Q(ram[1274]) );
  DFF_X1 ram_reg_79__9_ ( .D(n12242), .CK(clk), .Q(ram[1273]) );
  DFF_X1 ram_reg_79__8_ ( .D(n12241), .CK(clk), .Q(ram[1272]) );
  DFF_X1 ram_reg_79__7_ ( .D(n12240), .CK(clk), .Q(ram[1271]) );
  DFF_X1 ram_reg_79__6_ ( .D(n12239), .CK(clk), .Q(ram[1270]) );
  DFF_X1 ram_reg_79__5_ ( .D(n12238), .CK(clk), .Q(ram[1269]) );
  DFF_X1 ram_reg_79__4_ ( .D(n12237), .CK(clk), .Q(ram[1268]) );
  DFF_X1 ram_reg_79__3_ ( .D(n12236), .CK(clk), .Q(ram[1267]) );
  DFF_X1 ram_reg_79__2_ ( .D(n12235), .CK(clk), .Q(ram[1266]) );
  DFF_X1 ram_reg_79__1_ ( .D(n12234), .CK(clk), .Q(ram[1265]) );
  DFF_X1 ram_reg_79__0_ ( .D(n12233), .CK(clk), .Q(ram[1264]) );
  DFF_X1 ram_reg_78__15_ ( .D(n12265), .CK(clk), .Q(ram[1263]) );
  DFF_X1 ram_reg_78__14_ ( .D(n12264), .CK(clk), .Q(ram[1262]) );
  DFF_X1 ram_reg_78__13_ ( .D(n12263), .CK(clk), .Q(ram[1261]) );
  DFF_X1 ram_reg_78__12_ ( .D(n12262), .CK(clk), .Q(ram[1260]) );
  DFF_X1 ram_reg_78__11_ ( .D(n12261), .CK(clk), .Q(ram[1259]) );
  DFF_X1 ram_reg_78__10_ ( .D(n12260), .CK(clk), .Q(ram[1258]) );
  DFF_X1 ram_reg_78__9_ ( .D(n12259), .CK(clk), .Q(ram[1257]) );
  DFF_X1 ram_reg_78__8_ ( .D(n12258), .CK(clk), .Q(ram[1256]) );
  DFF_X1 ram_reg_78__7_ ( .D(n12257), .CK(clk), .Q(ram[1255]) );
  DFF_X1 ram_reg_78__6_ ( .D(n12256), .CK(clk), .Q(ram[1254]) );
  DFF_X1 ram_reg_78__5_ ( .D(n12255), .CK(clk), .Q(ram[1253]) );
  DFF_X1 ram_reg_78__4_ ( .D(n12254), .CK(clk), .Q(ram[1252]) );
  DFF_X1 ram_reg_78__3_ ( .D(n12253), .CK(clk), .Q(ram[1251]) );
  DFF_X1 ram_reg_78__2_ ( .D(n12252), .CK(clk), .Q(ram[1250]) );
  DFF_X1 ram_reg_78__1_ ( .D(n12251), .CK(clk), .Q(ram[1249]) );
  DFF_X1 ram_reg_78__0_ ( .D(n12250), .CK(clk), .Q(ram[1248]) );
  DFF_X1 ram_reg_77__15_ ( .D(n12282), .CK(clk), .Q(ram[1247]) );
  DFF_X1 ram_reg_77__14_ ( .D(n12281), .CK(clk), .Q(ram[1246]) );
  DFF_X1 ram_reg_77__13_ ( .D(n12280), .CK(clk), .Q(ram[1245]) );
  DFF_X1 ram_reg_77__12_ ( .D(n12279), .CK(clk), .Q(ram[1244]) );
  DFF_X1 ram_reg_77__11_ ( .D(n12278), .CK(clk), .Q(ram[1243]) );
  DFF_X1 ram_reg_77__10_ ( .D(n12277), .CK(clk), .Q(ram[1242]) );
  DFF_X1 ram_reg_77__9_ ( .D(n12276), .CK(clk), .Q(ram[1241]) );
  DFF_X1 ram_reg_77__8_ ( .D(n12275), .CK(clk), .Q(ram[1240]) );
  DFF_X1 ram_reg_77__7_ ( .D(n12274), .CK(clk), .Q(ram[1239]) );
  DFF_X1 ram_reg_77__6_ ( .D(n12273), .CK(clk), .Q(ram[1238]) );
  DFF_X1 ram_reg_77__5_ ( .D(n12272), .CK(clk), .Q(ram[1237]) );
  DFF_X1 ram_reg_77__4_ ( .D(n12271), .CK(clk), .Q(ram[1236]) );
  DFF_X1 ram_reg_77__3_ ( .D(n12270), .CK(clk), .Q(ram[1235]) );
  DFF_X1 ram_reg_77__2_ ( .D(n12269), .CK(clk), .Q(ram[1234]) );
  DFF_X1 ram_reg_77__1_ ( .D(n12268), .CK(clk), .Q(ram[1233]) );
  DFF_X1 ram_reg_77__0_ ( .D(n12267), .CK(clk), .Q(ram[1232]) );
  DFF_X1 ram_reg_76__15_ ( .D(n12299), .CK(clk), .Q(ram[1231]) );
  DFF_X1 ram_reg_76__14_ ( .D(n12298), .CK(clk), .Q(ram[1230]) );
  DFF_X1 ram_reg_76__13_ ( .D(n12297), .CK(clk), .Q(ram[1229]) );
  DFF_X1 ram_reg_76__12_ ( .D(n12296), .CK(clk), .Q(ram[1228]) );
  DFF_X1 ram_reg_76__11_ ( .D(n12295), .CK(clk), .Q(ram[1227]) );
  DFF_X1 ram_reg_76__10_ ( .D(n12294), .CK(clk), .Q(ram[1226]) );
  DFF_X1 ram_reg_76__9_ ( .D(n12293), .CK(clk), .Q(ram[1225]) );
  DFF_X1 ram_reg_76__8_ ( .D(n12292), .CK(clk), .Q(ram[1224]) );
  DFF_X1 ram_reg_76__7_ ( .D(n12291), .CK(clk), .Q(ram[1223]) );
  DFF_X1 ram_reg_76__6_ ( .D(n12290), .CK(clk), .Q(ram[1222]) );
  DFF_X1 ram_reg_76__5_ ( .D(n12289), .CK(clk), .Q(ram[1221]) );
  DFF_X1 ram_reg_76__4_ ( .D(n12288), .CK(clk), .Q(ram[1220]) );
  DFF_X1 ram_reg_76__3_ ( .D(n12287), .CK(clk), .Q(ram[1219]) );
  DFF_X1 ram_reg_76__2_ ( .D(n12286), .CK(clk), .Q(ram[1218]) );
  DFF_X1 ram_reg_76__1_ ( .D(n12285), .CK(clk), .Q(ram[1217]) );
  DFF_X1 ram_reg_76__0_ ( .D(n12284), .CK(clk), .Q(ram[1216]) );
  DFF_X1 ram_reg_75__15_ ( .D(n12316), .CK(clk), .Q(ram[1215]) );
  DFF_X1 ram_reg_75__14_ ( .D(n12315), .CK(clk), .Q(ram[1214]) );
  DFF_X1 ram_reg_75__13_ ( .D(n12314), .CK(clk), .Q(ram[1213]) );
  DFF_X1 ram_reg_75__12_ ( .D(n12313), .CK(clk), .Q(ram[1212]) );
  DFF_X1 ram_reg_75__11_ ( .D(n12312), .CK(clk), .Q(ram[1211]) );
  DFF_X1 ram_reg_75__10_ ( .D(n12311), .CK(clk), .Q(ram[1210]) );
  DFF_X1 ram_reg_75__9_ ( .D(n12310), .CK(clk), .Q(ram[1209]) );
  DFF_X1 ram_reg_75__8_ ( .D(n12309), .CK(clk), .Q(ram[1208]) );
  DFF_X1 ram_reg_75__7_ ( .D(n12308), .CK(clk), .Q(ram[1207]) );
  DFF_X1 ram_reg_75__6_ ( .D(n12307), .CK(clk), .Q(ram[1206]) );
  DFF_X1 ram_reg_75__5_ ( .D(n12306), .CK(clk), .Q(ram[1205]) );
  DFF_X1 ram_reg_75__4_ ( .D(n12305), .CK(clk), .Q(ram[1204]) );
  DFF_X1 ram_reg_75__3_ ( .D(n12304), .CK(clk), .Q(ram[1203]) );
  DFF_X1 ram_reg_75__2_ ( .D(n12303), .CK(clk), .Q(ram[1202]) );
  DFF_X1 ram_reg_75__1_ ( .D(n12302), .CK(clk), .Q(ram[1201]) );
  DFF_X1 ram_reg_75__0_ ( .D(n12301), .CK(clk), .Q(ram[1200]) );
  DFF_X1 ram_reg_74__15_ ( .D(n12333), .CK(clk), .Q(ram[1199]) );
  DFF_X1 ram_reg_74__14_ ( .D(n12332), .CK(clk), .Q(ram[1198]) );
  DFF_X1 ram_reg_74__13_ ( .D(n12331), .CK(clk), .Q(ram[1197]) );
  DFF_X1 ram_reg_74__12_ ( .D(n12330), .CK(clk), .Q(ram[1196]) );
  DFF_X1 ram_reg_74__11_ ( .D(n12329), .CK(clk), .Q(ram[1195]) );
  DFF_X1 ram_reg_74__10_ ( .D(n12328), .CK(clk), .Q(ram[1194]) );
  DFF_X1 ram_reg_74__9_ ( .D(n12327), .CK(clk), .Q(ram[1193]) );
  DFF_X1 ram_reg_74__8_ ( .D(n12326), .CK(clk), .Q(ram[1192]) );
  DFF_X1 ram_reg_74__7_ ( .D(n12325), .CK(clk), .Q(ram[1191]) );
  DFF_X1 ram_reg_74__6_ ( .D(n12324), .CK(clk), .Q(ram[1190]) );
  DFF_X1 ram_reg_74__5_ ( .D(n12323), .CK(clk), .Q(ram[1189]) );
  DFF_X1 ram_reg_74__4_ ( .D(n12322), .CK(clk), .Q(ram[1188]) );
  DFF_X1 ram_reg_74__3_ ( .D(n12321), .CK(clk), .Q(ram[1187]) );
  DFF_X1 ram_reg_74__2_ ( .D(n12320), .CK(clk), .Q(ram[1186]) );
  DFF_X1 ram_reg_74__1_ ( .D(n12319), .CK(clk), .Q(ram[1185]) );
  DFF_X1 ram_reg_74__0_ ( .D(n12318), .CK(clk), .Q(ram[1184]) );
  DFF_X1 ram_reg_73__15_ ( .D(n12350), .CK(clk), .Q(ram[1183]) );
  DFF_X1 ram_reg_73__14_ ( .D(n12349), .CK(clk), .Q(ram[1182]) );
  DFF_X1 ram_reg_73__13_ ( .D(n12348), .CK(clk), .Q(ram[1181]) );
  DFF_X1 ram_reg_73__12_ ( .D(n12347), .CK(clk), .Q(ram[1180]) );
  DFF_X1 ram_reg_73__11_ ( .D(n12346), .CK(clk), .Q(ram[1179]) );
  DFF_X1 ram_reg_73__10_ ( .D(n12345), .CK(clk), .Q(ram[1178]) );
  DFF_X1 ram_reg_73__9_ ( .D(n12344), .CK(clk), .Q(ram[1177]) );
  DFF_X1 ram_reg_73__8_ ( .D(n12343), .CK(clk), .Q(ram[1176]) );
  DFF_X1 ram_reg_73__7_ ( .D(n12342), .CK(clk), .Q(ram[1175]) );
  DFF_X1 ram_reg_73__6_ ( .D(n12341), .CK(clk), .Q(ram[1174]) );
  DFF_X1 ram_reg_73__5_ ( .D(n12340), .CK(clk), .Q(ram[1173]) );
  DFF_X1 ram_reg_73__4_ ( .D(n12339), .CK(clk), .Q(ram[1172]) );
  DFF_X1 ram_reg_73__3_ ( .D(n12338), .CK(clk), .Q(ram[1171]) );
  DFF_X1 ram_reg_73__2_ ( .D(n12337), .CK(clk), .Q(ram[1170]) );
  DFF_X1 ram_reg_73__1_ ( .D(n12336), .CK(clk), .Q(ram[1169]) );
  DFF_X1 ram_reg_73__0_ ( .D(n12335), .CK(clk), .Q(ram[1168]) );
  DFF_X1 ram_reg_72__15_ ( .D(n12367), .CK(clk), .Q(ram[1167]) );
  DFF_X1 ram_reg_72__14_ ( .D(n12366), .CK(clk), .Q(ram[1166]) );
  DFF_X1 ram_reg_72__13_ ( .D(n12365), .CK(clk), .Q(ram[1165]) );
  DFF_X1 ram_reg_72__12_ ( .D(n12364), .CK(clk), .Q(ram[1164]) );
  DFF_X1 ram_reg_72__11_ ( .D(n12363), .CK(clk), .Q(ram[1163]) );
  DFF_X1 ram_reg_72__10_ ( .D(n12362), .CK(clk), .Q(ram[1162]) );
  DFF_X1 ram_reg_72__9_ ( .D(n12361), .CK(clk), .Q(ram[1161]) );
  DFF_X1 ram_reg_72__8_ ( .D(n12360), .CK(clk), .Q(ram[1160]) );
  DFF_X1 ram_reg_72__7_ ( .D(n12359), .CK(clk), .Q(ram[1159]) );
  DFF_X1 ram_reg_72__6_ ( .D(n12358), .CK(clk), .Q(ram[1158]) );
  DFF_X1 ram_reg_72__5_ ( .D(n12357), .CK(clk), .Q(ram[1157]) );
  DFF_X1 ram_reg_72__4_ ( .D(n12356), .CK(clk), .Q(ram[1156]) );
  DFF_X1 ram_reg_72__3_ ( .D(n12355), .CK(clk), .Q(ram[1155]) );
  DFF_X1 ram_reg_72__2_ ( .D(n12354), .CK(clk), .Q(ram[1154]) );
  DFF_X1 ram_reg_72__1_ ( .D(n12353), .CK(clk), .Q(ram[1153]) );
  DFF_X1 ram_reg_72__0_ ( .D(n12352), .CK(clk), .Q(ram[1152]) );
  DFF_X1 ram_reg_71__15_ ( .D(n12384), .CK(clk), .Q(ram[1151]) );
  DFF_X1 ram_reg_71__14_ ( .D(n12383), .CK(clk), .Q(ram[1150]) );
  DFF_X1 ram_reg_71__13_ ( .D(n12382), .CK(clk), .Q(ram[1149]) );
  DFF_X1 ram_reg_71__12_ ( .D(n12381), .CK(clk), .Q(ram[1148]) );
  DFF_X1 ram_reg_71__11_ ( .D(n12380), .CK(clk), .Q(ram[1147]) );
  DFF_X1 ram_reg_71__10_ ( .D(n12379), .CK(clk), .Q(ram[1146]) );
  DFF_X1 ram_reg_71__9_ ( .D(n12378), .CK(clk), .Q(ram[1145]) );
  DFF_X1 ram_reg_71__8_ ( .D(n12377), .CK(clk), .Q(ram[1144]) );
  DFF_X1 ram_reg_71__7_ ( .D(n12376), .CK(clk), .Q(ram[1143]) );
  DFF_X1 ram_reg_71__6_ ( .D(n12375), .CK(clk), .Q(ram[1142]) );
  DFF_X1 ram_reg_71__5_ ( .D(n12374), .CK(clk), .Q(ram[1141]) );
  DFF_X1 ram_reg_71__4_ ( .D(n12373), .CK(clk), .Q(ram[1140]) );
  DFF_X1 ram_reg_71__3_ ( .D(n12372), .CK(clk), .Q(ram[1139]) );
  DFF_X1 ram_reg_71__2_ ( .D(n12371), .CK(clk), .Q(ram[1138]) );
  DFF_X1 ram_reg_71__1_ ( .D(n12370), .CK(clk), .Q(ram[1137]) );
  DFF_X1 ram_reg_71__0_ ( .D(n12369), .CK(clk), .Q(ram[1136]) );
  DFF_X1 ram_reg_70__15_ ( .D(n12401), .CK(clk), .Q(ram[1135]) );
  DFF_X1 ram_reg_70__14_ ( .D(n12400), .CK(clk), .Q(ram[1134]) );
  DFF_X1 ram_reg_70__13_ ( .D(n12399), .CK(clk), .Q(ram[1133]) );
  DFF_X1 ram_reg_70__12_ ( .D(n12398), .CK(clk), .Q(ram[1132]) );
  DFF_X1 ram_reg_70__11_ ( .D(n12397), .CK(clk), .Q(ram[1131]) );
  DFF_X1 ram_reg_70__10_ ( .D(n12396), .CK(clk), .Q(ram[1130]) );
  DFF_X1 ram_reg_70__9_ ( .D(n12395), .CK(clk), .Q(ram[1129]) );
  DFF_X1 ram_reg_70__8_ ( .D(n12394), .CK(clk), .Q(ram[1128]) );
  DFF_X1 ram_reg_70__7_ ( .D(n12393), .CK(clk), .Q(ram[1127]) );
  DFF_X1 ram_reg_70__6_ ( .D(n12392), .CK(clk), .Q(ram[1126]) );
  DFF_X1 ram_reg_70__5_ ( .D(n12391), .CK(clk), .Q(ram[1125]) );
  DFF_X1 ram_reg_70__4_ ( .D(n12390), .CK(clk), .Q(ram[1124]) );
  DFF_X1 ram_reg_70__3_ ( .D(n12389), .CK(clk), .Q(ram[1123]) );
  DFF_X1 ram_reg_70__2_ ( .D(n12388), .CK(clk), .Q(ram[1122]) );
  DFF_X1 ram_reg_70__1_ ( .D(n12387), .CK(clk), .Q(ram[1121]) );
  DFF_X1 ram_reg_70__0_ ( .D(n12386), .CK(clk), .Q(ram[1120]) );
  DFF_X1 ram_reg_69__15_ ( .D(n12418), .CK(clk), .Q(ram[1119]) );
  DFF_X1 ram_reg_69__14_ ( .D(n12417), .CK(clk), .Q(ram[1118]) );
  DFF_X1 ram_reg_69__13_ ( .D(n12416), .CK(clk), .Q(ram[1117]) );
  DFF_X1 ram_reg_69__12_ ( .D(n12415), .CK(clk), .Q(ram[1116]) );
  DFF_X1 ram_reg_69__11_ ( .D(n12414), .CK(clk), .Q(ram[1115]) );
  DFF_X1 ram_reg_69__10_ ( .D(n12413), .CK(clk), .Q(ram[1114]) );
  DFF_X1 ram_reg_69__9_ ( .D(n12412), .CK(clk), .Q(ram[1113]) );
  DFF_X1 ram_reg_69__8_ ( .D(n12411), .CK(clk), .Q(ram[1112]) );
  DFF_X1 ram_reg_69__7_ ( .D(n12410), .CK(clk), .Q(ram[1111]) );
  DFF_X1 ram_reg_69__6_ ( .D(n12409), .CK(clk), .Q(ram[1110]) );
  DFF_X1 ram_reg_69__5_ ( .D(n12408), .CK(clk), .Q(ram[1109]) );
  DFF_X1 ram_reg_69__4_ ( .D(n12407), .CK(clk), .Q(ram[1108]) );
  DFF_X1 ram_reg_69__3_ ( .D(n12406), .CK(clk), .Q(ram[1107]) );
  DFF_X1 ram_reg_69__2_ ( .D(n12405), .CK(clk), .Q(ram[1106]) );
  DFF_X1 ram_reg_69__1_ ( .D(n12404), .CK(clk), .Q(ram[1105]) );
  DFF_X1 ram_reg_69__0_ ( .D(n12403), .CK(clk), .Q(ram[1104]) );
  DFF_X1 ram_reg_68__15_ ( .D(n12435), .CK(clk), .Q(ram[1103]) );
  DFF_X1 ram_reg_68__14_ ( .D(n12434), .CK(clk), .Q(ram[1102]) );
  DFF_X1 ram_reg_68__13_ ( .D(n12433), .CK(clk), .Q(ram[1101]) );
  DFF_X1 ram_reg_68__12_ ( .D(n12432), .CK(clk), .Q(ram[1100]) );
  DFF_X1 ram_reg_68__11_ ( .D(n12431), .CK(clk), .Q(ram[1099]) );
  DFF_X1 ram_reg_68__10_ ( .D(n12430), .CK(clk), .Q(ram[1098]) );
  DFF_X1 ram_reg_68__9_ ( .D(n12429), .CK(clk), .Q(ram[1097]) );
  DFF_X1 ram_reg_68__8_ ( .D(n12428), .CK(clk), .Q(ram[1096]) );
  DFF_X1 ram_reg_68__7_ ( .D(n12427), .CK(clk), .Q(ram[1095]) );
  DFF_X1 ram_reg_68__6_ ( .D(n12426), .CK(clk), .Q(ram[1094]) );
  DFF_X1 ram_reg_68__5_ ( .D(n12425), .CK(clk), .Q(ram[1093]) );
  DFF_X1 ram_reg_68__4_ ( .D(n12424), .CK(clk), .Q(ram[1092]) );
  DFF_X1 ram_reg_68__3_ ( .D(n12423), .CK(clk), .Q(ram[1091]) );
  DFF_X1 ram_reg_68__2_ ( .D(n12422), .CK(clk), .Q(ram[1090]) );
  DFF_X1 ram_reg_68__1_ ( .D(n12421), .CK(clk), .Q(ram[1089]) );
  DFF_X1 ram_reg_68__0_ ( .D(n12420), .CK(clk), .Q(ram[1088]) );
  DFF_X1 ram_reg_67__15_ ( .D(n12452), .CK(clk), .Q(ram[1087]) );
  DFF_X1 ram_reg_67__14_ ( .D(n12451), .CK(clk), .Q(ram[1086]) );
  DFF_X1 ram_reg_67__13_ ( .D(n12450), .CK(clk), .Q(ram[1085]) );
  DFF_X1 ram_reg_67__12_ ( .D(n12449), .CK(clk), .Q(ram[1084]) );
  DFF_X1 ram_reg_67__11_ ( .D(n12448), .CK(clk), .Q(ram[1083]) );
  DFF_X1 ram_reg_67__10_ ( .D(n12447), .CK(clk), .Q(ram[1082]) );
  DFF_X1 ram_reg_67__9_ ( .D(n12446), .CK(clk), .Q(ram[1081]) );
  DFF_X1 ram_reg_67__8_ ( .D(n12445), .CK(clk), .Q(ram[1080]) );
  DFF_X1 ram_reg_67__7_ ( .D(n12444), .CK(clk), .Q(ram[1079]) );
  DFF_X1 ram_reg_67__6_ ( .D(n12443), .CK(clk), .Q(ram[1078]) );
  DFF_X1 ram_reg_67__5_ ( .D(n12442), .CK(clk), .Q(ram[1077]) );
  DFF_X1 ram_reg_67__4_ ( .D(n12441), .CK(clk), .Q(ram[1076]) );
  DFF_X1 ram_reg_67__3_ ( .D(n12440), .CK(clk), .Q(ram[1075]) );
  DFF_X1 ram_reg_67__2_ ( .D(n12439), .CK(clk), .Q(ram[1074]) );
  DFF_X1 ram_reg_67__1_ ( .D(n12438), .CK(clk), .Q(ram[1073]) );
  DFF_X1 ram_reg_67__0_ ( .D(n12437), .CK(clk), .Q(ram[1072]) );
  DFF_X1 ram_reg_66__15_ ( .D(n12469), .CK(clk), .Q(ram[1071]) );
  DFF_X1 ram_reg_66__14_ ( .D(n12468), .CK(clk), .Q(ram[1070]) );
  DFF_X1 ram_reg_66__13_ ( .D(n12467), .CK(clk), .Q(ram[1069]) );
  DFF_X1 ram_reg_66__12_ ( .D(n12466), .CK(clk), .Q(ram[1068]) );
  DFF_X1 ram_reg_66__11_ ( .D(n12465), .CK(clk), .Q(ram[1067]) );
  DFF_X1 ram_reg_66__10_ ( .D(n12464), .CK(clk), .Q(ram[1066]) );
  DFF_X1 ram_reg_66__9_ ( .D(n12463), .CK(clk), .Q(ram[1065]) );
  DFF_X1 ram_reg_66__8_ ( .D(n12462), .CK(clk), .Q(ram[1064]) );
  DFF_X1 ram_reg_66__7_ ( .D(n12461), .CK(clk), .Q(ram[1063]) );
  DFF_X1 ram_reg_66__6_ ( .D(n12460), .CK(clk), .Q(ram[1062]) );
  DFF_X1 ram_reg_66__5_ ( .D(n12459), .CK(clk), .Q(ram[1061]) );
  DFF_X1 ram_reg_66__4_ ( .D(n12458), .CK(clk), .Q(ram[1060]) );
  DFF_X1 ram_reg_66__3_ ( .D(n12457), .CK(clk), .Q(ram[1059]) );
  DFF_X1 ram_reg_66__2_ ( .D(n12456), .CK(clk), .Q(ram[1058]) );
  DFF_X1 ram_reg_66__1_ ( .D(n12455), .CK(clk), .Q(ram[1057]) );
  DFF_X1 ram_reg_66__0_ ( .D(n12454), .CK(clk), .Q(ram[1056]) );
  DFF_X1 ram_reg_65__15_ ( .D(n12486), .CK(clk), .Q(ram[1055]) );
  DFF_X1 ram_reg_65__14_ ( .D(n12485), .CK(clk), .Q(ram[1054]) );
  DFF_X1 ram_reg_65__13_ ( .D(n12484), .CK(clk), .Q(ram[1053]) );
  DFF_X1 ram_reg_65__12_ ( .D(n12483), .CK(clk), .Q(ram[1052]) );
  DFF_X1 ram_reg_65__11_ ( .D(n12482), .CK(clk), .Q(ram[1051]) );
  DFF_X1 ram_reg_65__10_ ( .D(n12481), .CK(clk), .Q(ram[1050]) );
  DFF_X1 ram_reg_65__9_ ( .D(n12480), .CK(clk), .Q(ram[1049]) );
  DFF_X1 ram_reg_65__8_ ( .D(n12479), .CK(clk), .Q(ram[1048]) );
  DFF_X1 ram_reg_65__7_ ( .D(n12478), .CK(clk), .Q(ram[1047]) );
  DFF_X1 ram_reg_65__6_ ( .D(n12477), .CK(clk), .Q(ram[1046]) );
  DFF_X1 ram_reg_65__5_ ( .D(n12476), .CK(clk), .Q(ram[1045]) );
  DFF_X1 ram_reg_65__4_ ( .D(n12475), .CK(clk), .Q(ram[1044]) );
  DFF_X1 ram_reg_65__3_ ( .D(n12474), .CK(clk), .Q(ram[1043]) );
  DFF_X1 ram_reg_65__2_ ( .D(n12473), .CK(clk), .Q(ram[1042]) );
  DFF_X1 ram_reg_65__1_ ( .D(n12472), .CK(clk), .Q(ram[1041]) );
  DFF_X1 ram_reg_65__0_ ( .D(n12471), .CK(clk), .Q(ram[1040]) );
  DFF_X1 ram_reg_64__15_ ( .D(n12503), .CK(clk), .Q(ram[1039]) );
  DFF_X1 ram_reg_64__14_ ( .D(n12502), .CK(clk), .Q(ram[1038]) );
  DFF_X1 ram_reg_64__13_ ( .D(n12501), .CK(clk), .Q(ram[1037]) );
  DFF_X1 ram_reg_64__12_ ( .D(n12500), .CK(clk), .Q(ram[1036]) );
  DFF_X1 ram_reg_64__11_ ( .D(n12499), .CK(clk), .Q(ram[1035]) );
  DFF_X1 ram_reg_64__10_ ( .D(n12498), .CK(clk), .Q(ram[1034]) );
  DFF_X1 ram_reg_64__9_ ( .D(n12497), .CK(clk), .Q(ram[1033]) );
  DFF_X1 ram_reg_64__8_ ( .D(n12496), .CK(clk), .Q(ram[1032]) );
  DFF_X1 ram_reg_64__7_ ( .D(n12495), .CK(clk), .Q(ram[1031]) );
  DFF_X1 ram_reg_64__6_ ( .D(n12494), .CK(clk), .Q(ram[1030]) );
  DFF_X1 ram_reg_64__5_ ( .D(n12493), .CK(clk), .Q(ram[1029]) );
  DFF_X1 ram_reg_64__4_ ( .D(n12492), .CK(clk), .Q(ram[1028]) );
  DFF_X1 ram_reg_64__3_ ( .D(n12491), .CK(clk), .Q(ram[1027]) );
  DFF_X1 ram_reg_64__2_ ( .D(n12490), .CK(clk), .Q(ram[1026]) );
  DFF_X1 ram_reg_64__1_ ( .D(n12489), .CK(clk), .Q(ram[1025]) );
  DFF_X1 ram_reg_64__0_ ( .D(n12488), .CK(clk), .Q(ram[1024]) );
  DFF_X1 ram_reg_63__15_ ( .D(n12520), .CK(clk), .Q(ram[1023]) );
  DFF_X1 ram_reg_63__14_ ( .D(n12519), .CK(clk), .Q(ram[1022]) );
  DFF_X1 ram_reg_63__13_ ( .D(n12518), .CK(clk), .Q(ram[1021]) );
  DFF_X1 ram_reg_63__12_ ( .D(n12517), .CK(clk), .Q(ram[1020]) );
  DFF_X1 ram_reg_63__11_ ( .D(n12516), .CK(clk), .Q(ram[1019]) );
  DFF_X1 ram_reg_63__10_ ( .D(n12515), .CK(clk), .Q(ram[1018]) );
  DFF_X1 ram_reg_63__9_ ( .D(n12514), .CK(clk), .Q(ram[1017]) );
  DFF_X1 ram_reg_63__8_ ( .D(n12513), .CK(clk), .Q(ram[1016]) );
  DFF_X1 ram_reg_63__7_ ( .D(n12512), .CK(clk), .Q(ram[1015]) );
  DFF_X1 ram_reg_63__6_ ( .D(n12511), .CK(clk), .Q(ram[1014]) );
  DFF_X1 ram_reg_63__5_ ( .D(n12510), .CK(clk), .Q(ram[1013]) );
  DFF_X1 ram_reg_63__4_ ( .D(n12509), .CK(clk), .Q(ram[1012]) );
  DFF_X1 ram_reg_63__3_ ( .D(n12508), .CK(clk), .Q(ram[1011]) );
  DFF_X1 ram_reg_63__2_ ( .D(n12507), .CK(clk), .Q(ram[1010]) );
  DFF_X1 ram_reg_63__1_ ( .D(n12506), .CK(clk), .Q(ram[1009]) );
  DFF_X1 ram_reg_63__0_ ( .D(n12505), .CK(clk), .Q(ram[1008]) );
  DFF_X1 ram_reg_62__15_ ( .D(n12537), .CK(clk), .Q(ram[1007]) );
  DFF_X1 ram_reg_62__14_ ( .D(n12536), .CK(clk), .Q(ram[1006]) );
  DFF_X1 ram_reg_62__13_ ( .D(n12535), .CK(clk), .Q(ram[1005]) );
  DFF_X1 ram_reg_62__12_ ( .D(n12534), .CK(clk), .Q(ram[1004]) );
  DFF_X1 ram_reg_62__11_ ( .D(n12533), .CK(clk), .Q(ram[1003]) );
  DFF_X1 ram_reg_62__10_ ( .D(n12532), .CK(clk), .Q(ram[1002]) );
  DFF_X1 ram_reg_62__9_ ( .D(n12531), .CK(clk), .Q(ram[1001]) );
  DFF_X1 ram_reg_62__8_ ( .D(n12530), .CK(clk), .Q(ram[1000]) );
  DFF_X1 ram_reg_62__7_ ( .D(n12529), .CK(clk), .Q(ram[999]) );
  DFF_X1 ram_reg_62__6_ ( .D(n12528), .CK(clk), .Q(ram[998]) );
  DFF_X1 ram_reg_62__5_ ( .D(n12527), .CK(clk), .Q(ram[997]) );
  DFF_X1 ram_reg_62__4_ ( .D(n12526), .CK(clk), .Q(ram[996]) );
  DFF_X1 ram_reg_62__3_ ( .D(n12525), .CK(clk), .Q(ram[995]) );
  DFF_X1 ram_reg_62__2_ ( .D(n12524), .CK(clk), .Q(ram[994]) );
  DFF_X1 ram_reg_62__1_ ( .D(n12523), .CK(clk), .Q(ram[993]) );
  DFF_X1 ram_reg_62__0_ ( .D(n12522), .CK(clk), .Q(ram[992]) );
  DFF_X1 ram_reg_61__15_ ( .D(n12554), .CK(clk), .Q(ram[991]) );
  DFF_X1 ram_reg_61__14_ ( .D(n12553), .CK(clk), .Q(ram[990]) );
  DFF_X1 ram_reg_61__13_ ( .D(n12552), .CK(clk), .Q(ram[989]) );
  DFF_X1 ram_reg_61__12_ ( .D(n12551), .CK(clk), .Q(ram[988]) );
  DFF_X1 ram_reg_61__11_ ( .D(n12550), .CK(clk), .Q(ram[987]) );
  DFF_X1 ram_reg_61__10_ ( .D(n12549), .CK(clk), .Q(ram[986]) );
  DFF_X1 ram_reg_61__9_ ( .D(n12548), .CK(clk), .Q(ram[985]) );
  DFF_X1 ram_reg_61__8_ ( .D(n12547), .CK(clk), .Q(ram[984]) );
  DFF_X1 ram_reg_61__7_ ( .D(n12546), .CK(clk), .Q(ram[983]) );
  DFF_X1 ram_reg_61__6_ ( .D(n12545), .CK(clk), .Q(ram[982]) );
  DFF_X1 ram_reg_61__5_ ( .D(n12544), .CK(clk), .Q(ram[981]) );
  DFF_X1 ram_reg_61__4_ ( .D(n12543), .CK(clk), .Q(ram[980]) );
  DFF_X1 ram_reg_61__3_ ( .D(n12542), .CK(clk), .Q(ram[979]) );
  DFF_X1 ram_reg_61__2_ ( .D(n12541), .CK(clk), .Q(ram[978]) );
  DFF_X1 ram_reg_61__1_ ( .D(n12540), .CK(clk), .Q(ram[977]) );
  DFF_X1 ram_reg_61__0_ ( .D(n12539), .CK(clk), .Q(ram[976]) );
  DFF_X1 ram_reg_60__15_ ( .D(n12571), .CK(clk), .Q(ram[975]) );
  DFF_X1 ram_reg_60__14_ ( .D(n12570), .CK(clk), .Q(ram[974]) );
  DFF_X1 ram_reg_60__13_ ( .D(n12569), .CK(clk), .Q(ram[973]) );
  DFF_X1 ram_reg_60__12_ ( .D(n12568), .CK(clk), .Q(ram[972]) );
  DFF_X1 ram_reg_60__11_ ( .D(n12567), .CK(clk), .Q(ram[971]) );
  DFF_X1 ram_reg_60__10_ ( .D(n12566), .CK(clk), .Q(ram[970]) );
  DFF_X1 ram_reg_60__9_ ( .D(n12565), .CK(clk), .Q(ram[969]) );
  DFF_X1 ram_reg_60__8_ ( .D(n12564), .CK(clk), .Q(ram[968]) );
  DFF_X1 ram_reg_60__7_ ( .D(n12563), .CK(clk), .Q(ram[967]) );
  DFF_X1 ram_reg_60__6_ ( .D(n12562), .CK(clk), .Q(ram[966]) );
  DFF_X1 ram_reg_60__5_ ( .D(n12561), .CK(clk), .Q(ram[965]) );
  DFF_X1 ram_reg_60__4_ ( .D(n12560), .CK(clk), .Q(ram[964]) );
  DFF_X1 ram_reg_60__3_ ( .D(n12559), .CK(clk), .Q(ram[963]) );
  DFF_X1 ram_reg_60__2_ ( .D(n12558), .CK(clk), .Q(ram[962]) );
  DFF_X1 ram_reg_60__1_ ( .D(n12557), .CK(clk), .Q(ram[961]) );
  DFF_X1 ram_reg_60__0_ ( .D(n12556), .CK(clk), .Q(ram[960]) );
  DFF_X1 ram_reg_59__15_ ( .D(n12588), .CK(clk), .Q(ram[959]) );
  DFF_X1 ram_reg_59__14_ ( .D(n12587), .CK(clk), .Q(ram[958]) );
  DFF_X1 ram_reg_59__13_ ( .D(n12586), .CK(clk), .Q(ram[957]) );
  DFF_X1 ram_reg_59__12_ ( .D(n12585), .CK(clk), .Q(ram[956]) );
  DFF_X1 ram_reg_59__11_ ( .D(n12584), .CK(clk), .Q(ram[955]) );
  DFF_X1 ram_reg_59__10_ ( .D(n12583), .CK(clk), .Q(ram[954]) );
  DFF_X1 ram_reg_59__9_ ( .D(n12582), .CK(clk), .Q(ram[953]) );
  DFF_X1 ram_reg_59__8_ ( .D(n12581), .CK(clk), .Q(ram[952]) );
  DFF_X1 ram_reg_59__7_ ( .D(n12580), .CK(clk), .Q(ram[951]) );
  DFF_X1 ram_reg_59__6_ ( .D(n12579), .CK(clk), .Q(ram[950]) );
  DFF_X1 ram_reg_59__5_ ( .D(n12578), .CK(clk), .Q(ram[949]) );
  DFF_X1 ram_reg_59__4_ ( .D(n12577), .CK(clk), .Q(ram[948]) );
  DFF_X1 ram_reg_59__3_ ( .D(n12576), .CK(clk), .Q(ram[947]) );
  DFF_X1 ram_reg_59__2_ ( .D(n12575), .CK(clk), .Q(ram[946]) );
  DFF_X1 ram_reg_59__1_ ( .D(n12574), .CK(clk), .Q(ram[945]) );
  DFF_X1 ram_reg_59__0_ ( .D(n12573), .CK(clk), .Q(ram[944]) );
  DFF_X1 ram_reg_58__15_ ( .D(n12605), .CK(clk), .Q(ram[943]) );
  DFF_X1 ram_reg_58__14_ ( .D(n12604), .CK(clk), .Q(ram[942]) );
  DFF_X1 ram_reg_58__13_ ( .D(n12603), .CK(clk), .Q(ram[941]) );
  DFF_X1 ram_reg_58__12_ ( .D(n12602), .CK(clk), .Q(ram[940]) );
  DFF_X1 ram_reg_58__11_ ( .D(n12601), .CK(clk), .Q(ram[939]) );
  DFF_X1 ram_reg_58__10_ ( .D(n12600), .CK(clk), .Q(ram[938]) );
  DFF_X1 ram_reg_58__9_ ( .D(n12599), .CK(clk), .Q(ram[937]) );
  DFF_X1 ram_reg_58__8_ ( .D(n12598), .CK(clk), .Q(ram[936]) );
  DFF_X1 ram_reg_58__7_ ( .D(n12597), .CK(clk), .Q(ram[935]) );
  DFF_X1 ram_reg_58__6_ ( .D(n12596), .CK(clk), .Q(ram[934]) );
  DFF_X1 ram_reg_58__5_ ( .D(n12595), .CK(clk), .Q(ram[933]) );
  DFF_X1 ram_reg_58__4_ ( .D(n12594), .CK(clk), .Q(ram[932]) );
  DFF_X1 ram_reg_58__3_ ( .D(n12593), .CK(clk), .Q(ram[931]) );
  DFF_X1 ram_reg_58__2_ ( .D(n12592), .CK(clk), .Q(ram[930]) );
  DFF_X1 ram_reg_58__1_ ( .D(n12591), .CK(clk), .Q(ram[929]) );
  DFF_X1 ram_reg_58__0_ ( .D(n12590), .CK(clk), .Q(ram[928]) );
  DFF_X1 ram_reg_57__15_ ( .D(n12622), .CK(clk), .Q(ram[927]) );
  DFF_X1 ram_reg_57__14_ ( .D(n12621), .CK(clk), .Q(ram[926]) );
  DFF_X1 ram_reg_57__13_ ( .D(n12620), .CK(clk), .Q(ram[925]) );
  DFF_X1 ram_reg_57__12_ ( .D(n12619), .CK(clk), .Q(ram[924]) );
  DFF_X1 ram_reg_57__11_ ( .D(n12618), .CK(clk), .Q(ram[923]) );
  DFF_X1 ram_reg_57__10_ ( .D(n12617), .CK(clk), .Q(ram[922]) );
  DFF_X1 ram_reg_57__9_ ( .D(n12616), .CK(clk), .Q(ram[921]) );
  DFF_X1 ram_reg_57__8_ ( .D(n12615), .CK(clk), .Q(ram[920]) );
  DFF_X1 ram_reg_57__7_ ( .D(n12614), .CK(clk), .Q(ram[919]) );
  DFF_X1 ram_reg_57__6_ ( .D(n12613), .CK(clk), .Q(ram[918]) );
  DFF_X1 ram_reg_57__5_ ( .D(n12612), .CK(clk), .Q(ram[917]) );
  DFF_X1 ram_reg_57__4_ ( .D(n12611), .CK(clk), .Q(ram[916]) );
  DFF_X1 ram_reg_57__3_ ( .D(n12610), .CK(clk), .Q(ram[915]) );
  DFF_X1 ram_reg_57__2_ ( .D(n12609), .CK(clk), .Q(ram[914]) );
  DFF_X1 ram_reg_57__1_ ( .D(n12608), .CK(clk), .Q(ram[913]) );
  DFF_X1 ram_reg_57__0_ ( .D(n12607), .CK(clk), .Q(ram[912]) );
  DFF_X1 ram_reg_56__15_ ( .D(n12639), .CK(clk), .Q(ram[911]) );
  DFF_X1 ram_reg_56__14_ ( .D(n12638), .CK(clk), .Q(ram[910]) );
  DFF_X1 ram_reg_56__13_ ( .D(n12637), .CK(clk), .Q(ram[909]) );
  DFF_X1 ram_reg_56__12_ ( .D(n12636), .CK(clk), .Q(ram[908]) );
  DFF_X1 ram_reg_56__11_ ( .D(n12635), .CK(clk), .Q(ram[907]) );
  DFF_X1 ram_reg_56__10_ ( .D(n12634), .CK(clk), .Q(ram[906]) );
  DFF_X1 ram_reg_56__9_ ( .D(n12633), .CK(clk), .Q(ram[905]) );
  DFF_X1 ram_reg_56__8_ ( .D(n12632), .CK(clk), .Q(ram[904]) );
  DFF_X1 ram_reg_56__7_ ( .D(n12631), .CK(clk), .Q(ram[903]) );
  DFF_X1 ram_reg_56__6_ ( .D(n12630), .CK(clk), .Q(ram[902]) );
  DFF_X1 ram_reg_56__5_ ( .D(n12629), .CK(clk), .Q(ram[901]) );
  DFF_X1 ram_reg_56__4_ ( .D(n12628), .CK(clk), .Q(ram[900]) );
  DFF_X1 ram_reg_56__3_ ( .D(n12627), .CK(clk), .Q(ram[899]) );
  DFF_X1 ram_reg_56__2_ ( .D(n12626), .CK(clk), .Q(ram[898]) );
  DFF_X1 ram_reg_56__1_ ( .D(n12625), .CK(clk), .Q(ram[897]) );
  DFF_X1 ram_reg_56__0_ ( .D(n12624), .CK(clk), .Q(ram[896]) );
  DFF_X1 ram_reg_55__15_ ( .D(n12656), .CK(clk), .Q(ram[895]) );
  DFF_X1 ram_reg_55__14_ ( .D(n12655), .CK(clk), .Q(ram[894]) );
  DFF_X1 ram_reg_55__13_ ( .D(n12654), .CK(clk), .Q(ram[893]) );
  DFF_X1 ram_reg_55__12_ ( .D(n12653), .CK(clk), .Q(ram[892]) );
  DFF_X1 ram_reg_55__11_ ( .D(n12652), .CK(clk), .Q(ram[891]) );
  DFF_X1 ram_reg_55__10_ ( .D(n12651), .CK(clk), .Q(ram[890]) );
  DFF_X1 ram_reg_55__9_ ( .D(n12650), .CK(clk), .Q(ram[889]) );
  DFF_X1 ram_reg_55__8_ ( .D(n12649), .CK(clk), .Q(ram[888]) );
  DFF_X1 ram_reg_55__7_ ( .D(n12648), .CK(clk), .Q(ram[887]) );
  DFF_X1 ram_reg_55__6_ ( .D(n12647), .CK(clk), .Q(ram[886]) );
  DFF_X1 ram_reg_55__5_ ( .D(n12646), .CK(clk), .Q(ram[885]) );
  DFF_X1 ram_reg_55__4_ ( .D(n12645), .CK(clk), .Q(ram[884]) );
  DFF_X1 ram_reg_55__3_ ( .D(n12644), .CK(clk), .Q(ram[883]) );
  DFF_X1 ram_reg_55__2_ ( .D(n12643), .CK(clk), .Q(ram[882]) );
  DFF_X1 ram_reg_55__1_ ( .D(n12642), .CK(clk), .Q(ram[881]) );
  DFF_X1 ram_reg_55__0_ ( .D(n12641), .CK(clk), .Q(ram[880]) );
  DFF_X1 ram_reg_54__15_ ( .D(n12673), .CK(clk), .Q(ram[879]) );
  DFF_X1 ram_reg_54__14_ ( .D(n12672), .CK(clk), .Q(ram[878]) );
  DFF_X1 ram_reg_54__13_ ( .D(n12671), .CK(clk), .Q(ram[877]) );
  DFF_X1 ram_reg_54__12_ ( .D(n12670), .CK(clk), .Q(ram[876]) );
  DFF_X1 ram_reg_54__11_ ( .D(n12669), .CK(clk), .Q(ram[875]) );
  DFF_X1 ram_reg_54__10_ ( .D(n12668), .CK(clk), .Q(ram[874]) );
  DFF_X1 ram_reg_54__9_ ( .D(n12667), .CK(clk), .Q(ram[873]) );
  DFF_X1 ram_reg_54__8_ ( .D(n12666), .CK(clk), .Q(ram[872]) );
  DFF_X1 ram_reg_54__7_ ( .D(n12665), .CK(clk), .Q(ram[871]) );
  DFF_X1 ram_reg_54__6_ ( .D(n12664), .CK(clk), .Q(ram[870]) );
  DFF_X1 ram_reg_54__5_ ( .D(n12663), .CK(clk), .Q(ram[869]) );
  DFF_X1 ram_reg_54__4_ ( .D(n12662), .CK(clk), .Q(ram[868]) );
  DFF_X1 ram_reg_54__3_ ( .D(n12661), .CK(clk), .Q(ram[867]) );
  DFF_X1 ram_reg_54__2_ ( .D(n12660), .CK(clk), .Q(ram[866]) );
  DFF_X1 ram_reg_54__1_ ( .D(n12659), .CK(clk), .Q(ram[865]) );
  DFF_X1 ram_reg_54__0_ ( .D(n12658), .CK(clk), .Q(ram[864]) );
  DFF_X1 ram_reg_53__15_ ( .D(n12690), .CK(clk), .Q(ram[863]) );
  DFF_X1 ram_reg_53__14_ ( .D(n12689), .CK(clk), .Q(ram[862]) );
  DFF_X1 ram_reg_53__13_ ( .D(n12688), .CK(clk), .Q(ram[861]) );
  DFF_X1 ram_reg_53__12_ ( .D(n12687), .CK(clk), .Q(ram[860]) );
  DFF_X1 ram_reg_53__11_ ( .D(n12686), .CK(clk), .Q(ram[859]) );
  DFF_X1 ram_reg_53__10_ ( .D(n12685), .CK(clk), .Q(ram[858]) );
  DFF_X1 ram_reg_53__9_ ( .D(n12684), .CK(clk), .Q(ram[857]) );
  DFF_X1 ram_reg_53__8_ ( .D(n12683), .CK(clk), .Q(ram[856]) );
  DFF_X1 ram_reg_53__7_ ( .D(n12682), .CK(clk), .Q(ram[855]) );
  DFF_X1 ram_reg_53__6_ ( .D(n12681), .CK(clk), .Q(ram[854]) );
  DFF_X1 ram_reg_53__5_ ( .D(n12680), .CK(clk), .Q(ram[853]) );
  DFF_X1 ram_reg_53__4_ ( .D(n12679), .CK(clk), .Q(ram[852]) );
  DFF_X1 ram_reg_53__3_ ( .D(n12678), .CK(clk), .Q(ram[851]) );
  DFF_X1 ram_reg_53__2_ ( .D(n12677), .CK(clk), .Q(ram[850]) );
  DFF_X1 ram_reg_53__1_ ( .D(n12676), .CK(clk), .Q(ram[849]) );
  DFF_X1 ram_reg_53__0_ ( .D(n12675), .CK(clk), .Q(ram[848]) );
  DFF_X1 ram_reg_52__15_ ( .D(n12707), .CK(clk), .Q(ram[847]) );
  DFF_X1 ram_reg_52__14_ ( .D(n12706), .CK(clk), .Q(ram[846]) );
  DFF_X1 ram_reg_52__13_ ( .D(n12705), .CK(clk), .Q(ram[845]) );
  DFF_X1 ram_reg_52__12_ ( .D(n12704), .CK(clk), .Q(ram[844]) );
  DFF_X1 ram_reg_52__11_ ( .D(n12703), .CK(clk), .Q(ram[843]) );
  DFF_X1 ram_reg_52__10_ ( .D(n12702), .CK(clk), .Q(ram[842]) );
  DFF_X1 ram_reg_52__9_ ( .D(n12701), .CK(clk), .Q(ram[841]) );
  DFF_X1 ram_reg_52__8_ ( .D(n12700), .CK(clk), .Q(ram[840]) );
  DFF_X1 ram_reg_52__7_ ( .D(n12699), .CK(clk), .Q(ram[839]) );
  DFF_X1 ram_reg_52__6_ ( .D(n12698), .CK(clk), .Q(ram[838]) );
  DFF_X1 ram_reg_52__5_ ( .D(n12697), .CK(clk), .Q(ram[837]) );
  DFF_X1 ram_reg_52__4_ ( .D(n12696), .CK(clk), .Q(ram[836]) );
  DFF_X1 ram_reg_52__3_ ( .D(n12695), .CK(clk), .Q(ram[835]) );
  DFF_X1 ram_reg_52__2_ ( .D(n12694), .CK(clk), .Q(ram[834]) );
  DFF_X1 ram_reg_52__1_ ( .D(n12693), .CK(clk), .Q(ram[833]) );
  DFF_X1 ram_reg_52__0_ ( .D(n12692), .CK(clk), .Q(ram[832]) );
  DFF_X1 ram_reg_51__15_ ( .D(n12724), .CK(clk), .Q(ram[831]) );
  DFF_X1 ram_reg_51__14_ ( .D(n12723), .CK(clk), .Q(ram[830]) );
  DFF_X1 ram_reg_51__13_ ( .D(n12722), .CK(clk), .Q(ram[829]) );
  DFF_X1 ram_reg_51__12_ ( .D(n12721), .CK(clk), .Q(ram[828]) );
  DFF_X1 ram_reg_51__11_ ( .D(n12720), .CK(clk), .Q(ram[827]) );
  DFF_X1 ram_reg_51__10_ ( .D(n12719), .CK(clk), .Q(ram[826]) );
  DFF_X1 ram_reg_51__9_ ( .D(n12718), .CK(clk), .Q(ram[825]) );
  DFF_X1 ram_reg_51__8_ ( .D(n12717), .CK(clk), .Q(ram[824]) );
  DFF_X1 ram_reg_51__7_ ( .D(n12716), .CK(clk), .Q(ram[823]) );
  DFF_X1 ram_reg_51__6_ ( .D(n12715), .CK(clk), .Q(ram[822]) );
  DFF_X1 ram_reg_51__5_ ( .D(n12714), .CK(clk), .Q(ram[821]) );
  DFF_X1 ram_reg_51__4_ ( .D(n12713), .CK(clk), .Q(ram[820]) );
  DFF_X1 ram_reg_51__3_ ( .D(n12712), .CK(clk), .Q(ram[819]) );
  DFF_X1 ram_reg_51__2_ ( .D(n12711), .CK(clk), .Q(ram[818]) );
  DFF_X1 ram_reg_51__1_ ( .D(n12710), .CK(clk), .Q(ram[817]) );
  DFF_X1 ram_reg_51__0_ ( .D(n12709), .CK(clk), .Q(ram[816]) );
  DFF_X1 ram_reg_50__15_ ( .D(n12741), .CK(clk), .Q(ram[815]) );
  DFF_X1 ram_reg_50__14_ ( .D(n12740), .CK(clk), .Q(ram[814]) );
  DFF_X1 ram_reg_50__13_ ( .D(n12739), .CK(clk), .Q(ram[813]) );
  DFF_X1 ram_reg_50__12_ ( .D(n12738), .CK(clk), .Q(ram[812]) );
  DFF_X1 ram_reg_50__11_ ( .D(n12737), .CK(clk), .Q(ram[811]) );
  DFF_X1 ram_reg_50__10_ ( .D(n12736), .CK(clk), .Q(ram[810]) );
  DFF_X1 ram_reg_50__9_ ( .D(n12735), .CK(clk), .Q(ram[809]) );
  DFF_X1 ram_reg_50__8_ ( .D(n12734), .CK(clk), .Q(ram[808]) );
  DFF_X1 ram_reg_50__7_ ( .D(n12733), .CK(clk), .Q(ram[807]) );
  DFF_X1 ram_reg_50__6_ ( .D(n12732), .CK(clk), .Q(ram[806]) );
  DFF_X1 ram_reg_50__5_ ( .D(n12731), .CK(clk), .Q(ram[805]) );
  DFF_X1 ram_reg_50__4_ ( .D(n12730), .CK(clk), .Q(ram[804]) );
  DFF_X1 ram_reg_50__3_ ( .D(n12729), .CK(clk), .Q(ram[803]) );
  DFF_X1 ram_reg_50__2_ ( .D(n12728), .CK(clk), .Q(ram[802]) );
  DFF_X1 ram_reg_50__1_ ( .D(n12727), .CK(clk), .Q(ram[801]) );
  DFF_X1 ram_reg_50__0_ ( .D(n12726), .CK(clk), .Q(ram[800]) );
  DFF_X1 ram_reg_49__15_ ( .D(n12758), .CK(clk), .Q(ram[799]) );
  DFF_X1 ram_reg_49__14_ ( .D(n12757), .CK(clk), .Q(ram[798]) );
  DFF_X1 ram_reg_49__13_ ( .D(n12756), .CK(clk), .Q(ram[797]) );
  DFF_X1 ram_reg_49__12_ ( .D(n12755), .CK(clk), .Q(ram[796]) );
  DFF_X1 ram_reg_49__11_ ( .D(n12754), .CK(clk), .Q(ram[795]) );
  DFF_X1 ram_reg_49__10_ ( .D(n12753), .CK(clk), .Q(ram[794]) );
  DFF_X1 ram_reg_49__9_ ( .D(n12752), .CK(clk), .Q(ram[793]) );
  DFF_X1 ram_reg_49__8_ ( .D(n12751), .CK(clk), .Q(ram[792]) );
  DFF_X1 ram_reg_49__7_ ( .D(n12750), .CK(clk), .Q(ram[791]) );
  DFF_X1 ram_reg_49__6_ ( .D(n12749), .CK(clk), .Q(ram[790]) );
  DFF_X1 ram_reg_49__5_ ( .D(n12748), .CK(clk), .Q(ram[789]) );
  DFF_X1 ram_reg_49__4_ ( .D(n12747), .CK(clk), .Q(ram[788]) );
  DFF_X1 ram_reg_49__3_ ( .D(n12746), .CK(clk), .Q(ram[787]) );
  DFF_X1 ram_reg_49__2_ ( .D(n12745), .CK(clk), .Q(ram[786]) );
  DFF_X1 ram_reg_49__1_ ( .D(n12744), .CK(clk), .Q(ram[785]) );
  DFF_X1 ram_reg_49__0_ ( .D(n12743), .CK(clk), .Q(ram[784]) );
  DFF_X1 ram_reg_48__15_ ( .D(n12775), .CK(clk), .Q(ram[783]) );
  DFF_X1 ram_reg_48__14_ ( .D(n12774), .CK(clk), .Q(ram[782]) );
  DFF_X1 ram_reg_48__13_ ( .D(n12773), .CK(clk), .Q(ram[781]) );
  DFF_X1 ram_reg_48__12_ ( .D(n12772), .CK(clk), .Q(ram[780]) );
  DFF_X1 ram_reg_48__11_ ( .D(n12771), .CK(clk), .Q(ram[779]) );
  DFF_X1 ram_reg_48__10_ ( .D(n12770), .CK(clk), .Q(ram[778]) );
  DFF_X1 ram_reg_48__9_ ( .D(n12769), .CK(clk), .Q(ram[777]) );
  DFF_X1 ram_reg_48__8_ ( .D(n12768), .CK(clk), .Q(ram[776]) );
  DFF_X1 ram_reg_48__7_ ( .D(n12767), .CK(clk), .Q(ram[775]) );
  DFF_X1 ram_reg_48__6_ ( .D(n12766), .CK(clk), .Q(ram[774]) );
  DFF_X1 ram_reg_48__5_ ( .D(n12765), .CK(clk), .Q(ram[773]) );
  DFF_X1 ram_reg_48__4_ ( .D(n12764), .CK(clk), .Q(ram[772]) );
  DFF_X1 ram_reg_48__3_ ( .D(n12763), .CK(clk), .Q(ram[771]) );
  DFF_X1 ram_reg_48__2_ ( .D(n12762), .CK(clk), .Q(ram[770]) );
  DFF_X1 ram_reg_48__1_ ( .D(n12761), .CK(clk), .Q(ram[769]) );
  DFF_X1 ram_reg_48__0_ ( .D(n12760), .CK(clk), .Q(ram[768]) );
  DFF_X1 ram_reg_47__15_ ( .D(n12792), .CK(clk), .Q(ram[767]) );
  DFF_X1 ram_reg_47__14_ ( .D(n12791), .CK(clk), .Q(ram[766]) );
  DFF_X1 ram_reg_47__13_ ( .D(n12790), .CK(clk), .Q(ram[765]) );
  DFF_X1 ram_reg_47__12_ ( .D(n12789), .CK(clk), .Q(ram[764]) );
  DFF_X1 ram_reg_47__11_ ( .D(n12788), .CK(clk), .Q(ram[763]) );
  DFF_X1 ram_reg_47__10_ ( .D(n12787), .CK(clk), .Q(ram[762]) );
  DFF_X1 ram_reg_47__9_ ( .D(n12786), .CK(clk), .Q(ram[761]) );
  DFF_X1 ram_reg_47__8_ ( .D(n12785), .CK(clk), .Q(ram[760]) );
  DFF_X1 ram_reg_47__7_ ( .D(n12784), .CK(clk), .Q(ram[759]) );
  DFF_X1 ram_reg_47__6_ ( .D(n12783), .CK(clk), .Q(ram[758]) );
  DFF_X1 ram_reg_47__5_ ( .D(n12782), .CK(clk), .Q(ram[757]) );
  DFF_X1 ram_reg_47__4_ ( .D(n12781), .CK(clk), .Q(ram[756]) );
  DFF_X1 ram_reg_47__3_ ( .D(n12780), .CK(clk), .Q(ram[755]) );
  DFF_X1 ram_reg_47__2_ ( .D(n12779), .CK(clk), .Q(ram[754]) );
  DFF_X1 ram_reg_47__1_ ( .D(n12778), .CK(clk), .Q(ram[753]) );
  DFF_X1 ram_reg_47__0_ ( .D(n12777), .CK(clk), .Q(ram[752]) );
  DFF_X1 ram_reg_46__15_ ( .D(n12809), .CK(clk), .Q(ram[751]) );
  DFF_X1 ram_reg_46__14_ ( .D(n12808), .CK(clk), .Q(ram[750]) );
  DFF_X1 ram_reg_46__13_ ( .D(n12807), .CK(clk), .Q(ram[749]) );
  DFF_X1 ram_reg_46__12_ ( .D(n12806), .CK(clk), .Q(ram[748]) );
  DFF_X1 ram_reg_46__11_ ( .D(n12805), .CK(clk), .Q(ram[747]) );
  DFF_X1 ram_reg_46__10_ ( .D(n12804), .CK(clk), .Q(ram[746]) );
  DFF_X1 ram_reg_46__9_ ( .D(n12803), .CK(clk), .Q(ram[745]) );
  DFF_X1 ram_reg_46__8_ ( .D(n12802), .CK(clk), .Q(ram[744]) );
  DFF_X1 ram_reg_46__7_ ( .D(n12801), .CK(clk), .Q(ram[743]) );
  DFF_X1 ram_reg_46__6_ ( .D(n12800), .CK(clk), .Q(ram[742]) );
  DFF_X1 ram_reg_46__5_ ( .D(n12799), .CK(clk), .Q(ram[741]) );
  DFF_X1 ram_reg_46__4_ ( .D(n12798), .CK(clk), .Q(ram[740]) );
  DFF_X1 ram_reg_46__3_ ( .D(n12797), .CK(clk), .Q(ram[739]) );
  DFF_X1 ram_reg_46__2_ ( .D(n12796), .CK(clk), .Q(ram[738]) );
  DFF_X1 ram_reg_46__1_ ( .D(n12795), .CK(clk), .Q(ram[737]) );
  DFF_X1 ram_reg_46__0_ ( .D(n12794), .CK(clk), .Q(ram[736]) );
  DFF_X1 ram_reg_45__15_ ( .D(n12826), .CK(clk), .Q(ram[735]) );
  DFF_X1 ram_reg_45__14_ ( .D(n12825), .CK(clk), .Q(ram[734]) );
  DFF_X1 ram_reg_45__13_ ( .D(n12824), .CK(clk), .Q(ram[733]) );
  DFF_X1 ram_reg_45__12_ ( .D(n12823), .CK(clk), .Q(ram[732]) );
  DFF_X1 ram_reg_45__11_ ( .D(n12822), .CK(clk), .Q(ram[731]) );
  DFF_X1 ram_reg_45__10_ ( .D(n12821), .CK(clk), .Q(ram[730]) );
  DFF_X1 ram_reg_45__9_ ( .D(n12820), .CK(clk), .Q(ram[729]) );
  DFF_X1 ram_reg_45__8_ ( .D(n12819), .CK(clk), .Q(ram[728]) );
  DFF_X1 ram_reg_45__7_ ( .D(n12818), .CK(clk), .Q(ram[727]) );
  DFF_X1 ram_reg_45__6_ ( .D(n12817), .CK(clk), .Q(ram[726]) );
  DFF_X1 ram_reg_45__5_ ( .D(n12816), .CK(clk), .Q(ram[725]) );
  DFF_X1 ram_reg_45__4_ ( .D(n12815), .CK(clk), .Q(ram[724]) );
  DFF_X1 ram_reg_45__3_ ( .D(n12814), .CK(clk), .Q(ram[723]) );
  DFF_X1 ram_reg_45__2_ ( .D(n12813), .CK(clk), .Q(ram[722]) );
  DFF_X1 ram_reg_45__1_ ( .D(n12812), .CK(clk), .Q(ram[721]) );
  DFF_X1 ram_reg_45__0_ ( .D(n12811), .CK(clk), .Q(ram[720]) );
  DFF_X1 ram_reg_44__15_ ( .D(n12843), .CK(clk), .Q(ram[719]) );
  DFF_X1 ram_reg_44__14_ ( .D(n12842), .CK(clk), .Q(ram[718]) );
  DFF_X1 ram_reg_44__13_ ( .D(n12841), .CK(clk), .Q(ram[717]) );
  DFF_X1 ram_reg_44__12_ ( .D(n12840), .CK(clk), .Q(ram[716]) );
  DFF_X1 ram_reg_44__11_ ( .D(n12839), .CK(clk), .Q(ram[715]) );
  DFF_X1 ram_reg_44__10_ ( .D(n12838), .CK(clk), .Q(ram[714]) );
  DFF_X1 ram_reg_44__9_ ( .D(n12837), .CK(clk), .Q(ram[713]) );
  DFF_X1 ram_reg_44__8_ ( .D(n12836), .CK(clk), .Q(ram[712]) );
  DFF_X1 ram_reg_44__7_ ( .D(n12835), .CK(clk), .Q(ram[711]) );
  DFF_X1 ram_reg_44__6_ ( .D(n12834), .CK(clk), .Q(ram[710]) );
  DFF_X1 ram_reg_44__5_ ( .D(n12833), .CK(clk), .Q(ram[709]) );
  DFF_X1 ram_reg_44__4_ ( .D(n12832), .CK(clk), .Q(ram[708]) );
  DFF_X1 ram_reg_44__3_ ( .D(n12831), .CK(clk), .Q(ram[707]) );
  DFF_X1 ram_reg_44__2_ ( .D(n12830), .CK(clk), .Q(ram[706]) );
  DFF_X1 ram_reg_44__1_ ( .D(n12829), .CK(clk), .Q(ram[705]) );
  DFF_X1 ram_reg_44__0_ ( .D(n12828), .CK(clk), .Q(ram[704]) );
  DFF_X1 ram_reg_43__15_ ( .D(n12860), .CK(clk), .Q(ram[703]) );
  DFF_X1 ram_reg_43__14_ ( .D(n12859), .CK(clk), .Q(ram[702]) );
  DFF_X1 ram_reg_43__13_ ( .D(n12858), .CK(clk), .Q(ram[701]) );
  DFF_X1 ram_reg_43__12_ ( .D(n12857), .CK(clk), .Q(ram[700]) );
  DFF_X1 ram_reg_43__11_ ( .D(n12856), .CK(clk), .Q(ram[699]) );
  DFF_X1 ram_reg_43__10_ ( .D(n12855), .CK(clk), .Q(ram[698]) );
  DFF_X1 ram_reg_43__9_ ( .D(n12854), .CK(clk), .Q(ram[697]) );
  DFF_X1 ram_reg_43__8_ ( .D(n12853), .CK(clk), .Q(ram[696]) );
  DFF_X1 ram_reg_43__7_ ( .D(n12852), .CK(clk), .Q(ram[695]) );
  DFF_X1 ram_reg_43__6_ ( .D(n12851), .CK(clk), .Q(ram[694]) );
  DFF_X1 ram_reg_43__5_ ( .D(n12850), .CK(clk), .Q(ram[693]) );
  DFF_X1 ram_reg_43__4_ ( .D(n12849), .CK(clk), .Q(ram[692]) );
  DFF_X1 ram_reg_43__3_ ( .D(n12848), .CK(clk), .Q(ram[691]) );
  DFF_X1 ram_reg_43__2_ ( .D(n12847), .CK(clk), .Q(ram[690]) );
  DFF_X1 ram_reg_43__1_ ( .D(n12846), .CK(clk), .Q(ram[689]) );
  DFF_X1 ram_reg_43__0_ ( .D(n12845), .CK(clk), .Q(ram[688]) );
  DFF_X1 ram_reg_42__15_ ( .D(n12877), .CK(clk), .Q(ram[687]) );
  DFF_X1 ram_reg_42__14_ ( .D(n12876), .CK(clk), .Q(ram[686]) );
  DFF_X1 ram_reg_42__13_ ( .D(n12875), .CK(clk), .Q(ram[685]) );
  DFF_X1 ram_reg_42__12_ ( .D(n12874), .CK(clk), .Q(ram[684]) );
  DFF_X1 ram_reg_42__11_ ( .D(n12873), .CK(clk), .Q(ram[683]) );
  DFF_X1 ram_reg_42__10_ ( .D(n12872), .CK(clk), .Q(ram[682]) );
  DFF_X1 ram_reg_42__9_ ( .D(n12871), .CK(clk), .Q(ram[681]) );
  DFF_X1 ram_reg_42__8_ ( .D(n12870), .CK(clk), .Q(ram[680]) );
  DFF_X1 ram_reg_42__7_ ( .D(n12869), .CK(clk), .Q(ram[679]) );
  DFF_X1 ram_reg_42__6_ ( .D(n12868), .CK(clk), .Q(ram[678]) );
  DFF_X1 ram_reg_42__5_ ( .D(n12867), .CK(clk), .Q(ram[677]) );
  DFF_X1 ram_reg_42__4_ ( .D(n12866), .CK(clk), .Q(ram[676]) );
  DFF_X1 ram_reg_42__3_ ( .D(n12865), .CK(clk), .Q(ram[675]) );
  DFF_X1 ram_reg_42__2_ ( .D(n12864), .CK(clk), .Q(ram[674]) );
  DFF_X1 ram_reg_42__1_ ( .D(n12863), .CK(clk), .Q(ram[673]) );
  DFF_X1 ram_reg_42__0_ ( .D(n12862), .CK(clk), .Q(ram[672]) );
  DFF_X1 ram_reg_41__15_ ( .D(n12894), .CK(clk), .Q(ram[671]) );
  DFF_X1 ram_reg_41__14_ ( .D(n12893), .CK(clk), .Q(ram[670]) );
  DFF_X1 ram_reg_41__13_ ( .D(n12892), .CK(clk), .Q(ram[669]) );
  DFF_X1 ram_reg_41__12_ ( .D(n12891), .CK(clk), .Q(ram[668]) );
  DFF_X1 ram_reg_41__11_ ( .D(n12890), .CK(clk), .Q(ram[667]) );
  DFF_X1 ram_reg_41__10_ ( .D(n12889), .CK(clk), .Q(ram[666]) );
  DFF_X1 ram_reg_41__9_ ( .D(n12888), .CK(clk), .Q(ram[665]) );
  DFF_X1 ram_reg_41__8_ ( .D(n12887), .CK(clk), .Q(ram[664]) );
  DFF_X1 ram_reg_41__7_ ( .D(n12886), .CK(clk), .Q(ram[663]) );
  DFF_X1 ram_reg_41__6_ ( .D(n12885), .CK(clk), .Q(ram[662]) );
  DFF_X1 ram_reg_41__5_ ( .D(n12884), .CK(clk), .Q(ram[661]) );
  DFF_X1 ram_reg_41__4_ ( .D(n12883), .CK(clk), .Q(ram[660]) );
  DFF_X1 ram_reg_41__3_ ( .D(n12882), .CK(clk), .Q(ram[659]) );
  DFF_X1 ram_reg_41__2_ ( .D(n12881), .CK(clk), .Q(ram[658]) );
  DFF_X1 ram_reg_41__1_ ( .D(n12880), .CK(clk), .Q(ram[657]) );
  DFF_X1 ram_reg_41__0_ ( .D(n12879), .CK(clk), .Q(ram[656]) );
  DFF_X1 ram_reg_40__15_ ( .D(n12911), .CK(clk), .Q(ram[655]) );
  DFF_X1 ram_reg_40__14_ ( .D(n12910), .CK(clk), .Q(ram[654]) );
  DFF_X1 ram_reg_40__13_ ( .D(n12909), .CK(clk), .Q(ram[653]) );
  DFF_X1 ram_reg_40__12_ ( .D(n12908), .CK(clk), .Q(ram[652]) );
  DFF_X1 ram_reg_40__11_ ( .D(n12907), .CK(clk), .Q(ram[651]) );
  DFF_X1 ram_reg_40__10_ ( .D(n12906), .CK(clk), .Q(ram[650]) );
  DFF_X1 ram_reg_40__9_ ( .D(n12905), .CK(clk), .Q(ram[649]) );
  DFF_X1 ram_reg_40__8_ ( .D(n12904), .CK(clk), .Q(ram[648]) );
  DFF_X1 ram_reg_40__7_ ( .D(n12903), .CK(clk), .Q(ram[647]) );
  DFF_X1 ram_reg_40__6_ ( .D(n12902), .CK(clk), .Q(ram[646]) );
  DFF_X1 ram_reg_40__5_ ( .D(n12901), .CK(clk), .Q(ram[645]) );
  DFF_X1 ram_reg_40__4_ ( .D(n12900), .CK(clk), .Q(ram[644]) );
  DFF_X1 ram_reg_40__3_ ( .D(n12899), .CK(clk), .Q(ram[643]) );
  DFF_X1 ram_reg_40__2_ ( .D(n12898), .CK(clk), .Q(ram[642]) );
  DFF_X1 ram_reg_40__1_ ( .D(n12897), .CK(clk), .Q(ram[641]) );
  DFF_X1 ram_reg_40__0_ ( .D(n12896), .CK(clk), .Q(ram[640]) );
  DFF_X1 ram_reg_39__15_ ( .D(n12928), .CK(clk), .Q(ram[639]) );
  DFF_X1 ram_reg_39__14_ ( .D(n12927), .CK(clk), .Q(ram[638]) );
  DFF_X1 ram_reg_39__13_ ( .D(n12926), .CK(clk), .Q(ram[637]) );
  DFF_X1 ram_reg_39__12_ ( .D(n12925), .CK(clk), .Q(ram[636]) );
  DFF_X1 ram_reg_39__11_ ( .D(n12924), .CK(clk), .Q(ram[635]) );
  DFF_X1 ram_reg_39__10_ ( .D(n12923), .CK(clk), .Q(ram[634]) );
  DFF_X1 ram_reg_39__9_ ( .D(n12922), .CK(clk), .Q(ram[633]) );
  DFF_X1 ram_reg_39__8_ ( .D(n12921), .CK(clk), .Q(ram[632]) );
  DFF_X1 ram_reg_39__7_ ( .D(n12920), .CK(clk), .Q(ram[631]) );
  DFF_X1 ram_reg_39__6_ ( .D(n12919), .CK(clk), .Q(ram[630]) );
  DFF_X1 ram_reg_39__5_ ( .D(n12918), .CK(clk), .Q(ram[629]) );
  DFF_X1 ram_reg_39__4_ ( .D(n12917), .CK(clk), .Q(ram[628]) );
  DFF_X1 ram_reg_39__3_ ( .D(n12916), .CK(clk), .Q(ram[627]) );
  DFF_X1 ram_reg_39__2_ ( .D(n12915), .CK(clk), .Q(ram[626]) );
  DFF_X1 ram_reg_39__1_ ( .D(n12914), .CK(clk), .Q(ram[625]) );
  DFF_X1 ram_reg_39__0_ ( .D(n12913), .CK(clk), .Q(ram[624]) );
  DFF_X1 ram_reg_38__15_ ( .D(n12945), .CK(clk), .Q(ram[623]) );
  DFF_X1 ram_reg_38__14_ ( .D(n12944), .CK(clk), .Q(ram[622]) );
  DFF_X1 ram_reg_38__13_ ( .D(n12943), .CK(clk), .Q(ram[621]) );
  DFF_X1 ram_reg_38__12_ ( .D(n12942), .CK(clk), .Q(ram[620]) );
  DFF_X1 ram_reg_38__11_ ( .D(n12941), .CK(clk), .Q(ram[619]) );
  DFF_X1 ram_reg_38__10_ ( .D(n12940), .CK(clk), .Q(ram[618]) );
  DFF_X1 ram_reg_38__9_ ( .D(n12939), .CK(clk), .Q(ram[617]) );
  DFF_X1 ram_reg_38__8_ ( .D(n12938), .CK(clk), .Q(ram[616]) );
  DFF_X1 ram_reg_38__7_ ( .D(n12937), .CK(clk), .Q(ram[615]) );
  DFF_X1 ram_reg_38__6_ ( .D(n12936), .CK(clk), .Q(ram[614]) );
  DFF_X1 ram_reg_38__5_ ( .D(n12935), .CK(clk), .Q(ram[613]) );
  DFF_X1 ram_reg_38__4_ ( .D(n12934), .CK(clk), .Q(ram[612]) );
  DFF_X1 ram_reg_38__3_ ( .D(n12933), .CK(clk), .Q(ram[611]) );
  DFF_X1 ram_reg_38__2_ ( .D(n12932), .CK(clk), .Q(ram[610]) );
  DFF_X1 ram_reg_38__1_ ( .D(n12931), .CK(clk), .Q(ram[609]) );
  DFF_X1 ram_reg_38__0_ ( .D(n12930), .CK(clk), .Q(ram[608]) );
  DFF_X1 ram_reg_37__15_ ( .D(n12962), .CK(clk), .Q(ram[607]) );
  DFF_X1 ram_reg_37__14_ ( .D(n12961), .CK(clk), .Q(ram[606]) );
  DFF_X1 ram_reg_37__13_ ( .D(n12960), .CK(clk), .Q(ram[605]) );
  DFF_X1 ram_reg_37__12_ ( .D(n12959), .CK(clk), .Q(ram[604]) );
  DFF_X1 ram_reg_37__11_ ( .D(n12958), .CK(clk), .Q(ram[603]) );
  DFF_X1 ram_reg_37__10_ ( .D(n12957), .CK(clk), .Q(ram[602]) );
  DFF_X1 ram_reg_37__9_ ( .D(n12956), .CK(clk), .Q(ram[601]) );
  DFF_X1 ram_reg_37__8_ ( .D(n12955), .CK(clk), .Q(ram[600]) );
  DFF_X1 ram_reg_37__7_ ( .D(n12954), .CK(clk), .Q(ram[599]) );
  DFF_X1 ram_reg_37__6_ ( .D(n12953), .CK(clk), .Q(ram[598]) );
  DFF_X1 ram_reg_37__5_ ( .D(n12952), .CK(clk), .Q(ram[597]) );
  DFF_X1 ram_reg_37__4_ ( .D(n12951), .CK(clk), .Q(ram[596]) );
  DFF_X1 ram_reg_37__3_ ( .D(n12950), .CK(clk), .Q(ram[595]) );
  DFF_X1 ram_reg_37__2_ ( .D(n12949), .CK(clk), .Q(ram[594]) );
  DFF_X1 ram_reg_37__1_ ( .D(n12948), .CK(clk), .Q(ram[593]) );
  DFF_X1 ram_reg_37__0_ ( .D(n12947), .CK(clk), .Q(ram[592]) );
  DFF_X1 ram_reg_36__15_ ( .D(n12979), .CK(clk), .Q(ram[591]) );
  DFF_X1 ram_reg_36__14_ ( .D(n12978), .CK(clk), .Q(ram[590]) );
  DFF_X1 ram_reg_36__13_ ( .D(n12977), .CK(clk), .Q(ram[589]) );
  DFF_X1 ram_reg_36__12_ ( .D(n12976), .CK(clk), .Q(ram[588]) );
  DFF_X1 ram_reg_36__11_ ( .D(n12975), .CK(clk), .Q(ram[587]) );
  DFF_X1 ram_reg_36__10_ ( .D(n12974), .CK(clk), .Q(ram[586]) );
  DFF_X1 ram_reg_36__9_ ( .D(n12973), .CK(clk), .Q(ram[585]) );
  DFF_X1 ram_reg_36__8_ ( .D(n12972), .CK(clk), .Q(ram[584]) );
  DFF_X1 ram_reg_36__7_ ( .D(n12971), .CK(clk), .Q(ram[583]) );
  DFF_X1 ram_reg_36__6_ ( .D(n12970), .CK(clk), .Q(ram[582]) );
  DFF_X1 ram_reg_36__5_ ( .D(n12969), .CK(clk), .Q(ram[581]) );
  DFF_X1 ram_reg_36__4_ ( .D(n12968), .CK(clk), .Q(ram[580]) );
  DFF_X1 ram_reg_36__3_ ( .D(n12967), .CK(clk), .Q(ram[579]) );
  DFF_X1 ram_reg_36__2_ ( .D(n12966), .CK(clk), .Q(ram[578]) );
  DFF_X1 ram_reg_36__1_ ( .D(n12965), .CK(clk), .Q(ram[577]) );
  DFF_X1 ram_reg_36__0_ ( .D(n12964), .CK(clk), .Q(ram[576]) );
  DFF_X1 ram_reg_35__15_ ( .D(n12996), .CK(clk), .Q(ram[575]) );
  DFF_X1 ram_reg_35__14_ ( .D(n12995), .CK(clk), .Q(ram[574]) );
  DFF_X1 ram_reg_35__13_ ( .D(n12994), .CK(clk), .Q(ram[573]) );
  DFF_X1 ram_reg_35__12_ ( .D(n12993), .CK(clk), .Q(ram[572]) );
  DFF_X1 ram_reg_35__11_ ( .D(n12992), .CK(clk), .Q(ram[571]) );
  DFF_X1 ram_reg_35__10_ ( .D(n12991), .CK(clk), .Q(ram[570]) );
  DFF_X1 ram_reg_35__9_ ( .D(n12990), .CK(clk), .Q(ram[569]) );
  DFF_X1 ram_reg_35__8_ ( .D(n12989), .CK(clk), .Q(ram[568]) );
  DFF_X1 ram_reg_35__7_ ( .D(n12988), .CK(clk), .Q(ram[567]) );
  DFF_X1 ram_reg_35__6_ ( .D(n12987), .CK(clk), .Q(ram[566]) );
  DFF_X1 ram_reg_35__5_ ( .D(n12986), .CK(clk), .Q(ram[565]) );
  DFF_X1 ram_reg_35__4_ ( .D(n12985), .CK(clk), .Q(ram[564]) );
  DFF_X1 ram_reg_35__3_ ( .D(n12984), .CK(clk), .Q(ram[563]) );
  DFF_X1 ram_reg_35__2_ ( .D(n12983), .CK(clk), .Q(ram[562]) );
  DFF_X1 ram_reg_35__1_ ( .D(n12982), .CK(clk), .Q(ram[561]) );
  DFF_X1 ram_reg_35__0_ ( .D(n12981), .CK(clk), .Q(ram[560]) );
  DFF_X1 ram_reg_34__15_ ( .D(n13013), .CK(clk), .Q(ram[559]) );
  DFF_X1 ram_reg_34__14_ ( .D(n13012), .CK(clk), .Q(ram[558]) );
  DFF_X1 ram_reg_34__13_ ( .D(n13011), .CK(clk), .Q(ram[557]) );
  DFF_X1 ram_reg_34__12_ ( .D(n13010), .CK(clk), .Q(ram[556]) );
  DFF_X1 ram_reg_34__11_ ( .D(n13009), .CK(clk), .Q(ram[555]) );
  DFF_X1 ram_reg_34__10_ ( .D(n13008), .CK(clk), .Q(ram[554]) );
  DFF_X1 ram_reg_34__9_ ( .D(n13007), .CK(clk), .Q(ram[553]) );
  DFF_X1 ram_reg_34__8_ ( .D(n13006), .CK(clk), .Q(ram[552]) );
  DFF_X1 ram_reg_34__7_ ( .D(n13005), .CK(clk), .Q(ram[551]) );
  DFF_X1 ram_reg_34__6_ ( .D(n13004), .CK(clk), .Q(ram[550]) );
  DFF_X1 ram_reg_34__5_ ( .D(n13003), .CK(clk), .Q(ram[549]) );
  DFF_X1 ram_reg_34__4_ ( .D(n13002), .CK(clk), .Q(ram[548]) );
  DFF_X1 ram_reg_34__3_ ( .D(n13001), .CK(clk), .Q(ram[547]) );
  DFF_X1 ram_reg_34__2_ ( .D(n13000), .CK(clk), .Q(ram[546]) );
  DFF_X1 ram_reg_34__1_ ( .D(n12999), .CK(clk), .Q(ram[545]) );
  DFF_X1 ram_reg_34__0_ ( .D(n12998), .CK(clk), .Q(ram[544]) );
  DFF_X1 ram_reg_33__15_ ( .D(n13030), .CK(clk), .Q(ram[543]) );
  DFF_X1 ram_reg_33__14_ ( .D(n13029), .CK(clk), .Q(ram[542]) );
  DFF_X1 ram_reg_33__13_ ( .D(n13028), .CK(clk), .Q(ram[541]) );
  DFF_X1 ram_reg_33__12_ ( .D(n13027), .CK(clk), .Q(ram[540]) );
  DFF_X1 ram_reg_33__11_ ( .D(n13026), .CK(clk), .Q(ram[539]) );
  DFF_X1 ram_reg_33__10_ ( .D(n13025), .CK(clk), .Q(ram[538]) );
  DFF_X1 ram_reg_33__9_ ( .D(n13024), .CK(clk), .Q(ram[537]) );
  DFF_X1 ram_reg_33__8_ ( .D(n13023), .CK(clk), .Q(ram[536]) );
  DFF_X1 ram_reg_33__7_ ( .D(n13022), .CK(clk), .Q(ram[535]) );
  DFF_X1 ram_reg_33__6_ ( .D(n13021), .CK(clk), .Q(ram[534]) );
  DFF_X1 ram_reg_33__5_ ( .D(n13020), .CK(clk), .Q(ram[533]) );
  DFF_X1 ram_reg_33__4_ ( .D(n13019), .CK(clk), .Q(ram[532]) );
  DFF_X1 ram_reg_33__3_ ( .D(n13018), .CK(clk), .Q(ram[531]) );
  DFF_X1 ram_reg_33__2_ ( .D(n13017), .CK(clk), .Q(ram[530]) );
  DFF_X1 ram_reg_33__1_ ( .D(n13016), .CK(clk), .Q(ram[529]) );
  DFF_X1 ram_reg_33__0_ ( .D(n13015), .CK(clk), .Q(ram[528]) );
  DFF_X1 ram_reg_32__15_ ( .D(n13047), .CK(clk), .Q(ram[527]) );
  DFF_X1 ram_reg_32__14_ ( .D(n13046), .CK(clk), .Q(ram[526]) );
  DFF_X1 ram_reg_32__13_ ( .D(n13045), .CK(clk), .Q(ram[525]) );
  DFF_X1 ram_reg_32__12_ ( .D(n13044), .CK(clk), .Q(ram[524]) );
  DFF_X1 ram_reg_32__11_ ( .D(n13043), .CK(clk), .Q(ram[523]) );
  DFF_X1 ram_reg_32__10_ ( .D(n13042), .CK(clk), .Q(ram[522]) );
  DFF_X1 ram_reg_32__9_ ( .D(n13041), .CK(clk), .Q(ram[521]) );
  DFF_X1 ram_reg_32__8_ ( .D(n13040), .CK(clk), .Q(ram[520]) );
  DFF_X1 ram_reg_32__7_ ( .D(n13039), .CK(clk), .Q(ram[519]) );
  DFF_X1 ram_reg_32__6_ ( .D(n13038), .CK(clk), .Q(ram[518]) );
  DFF_X1 ram_reg_32__5_ ( .D(n13037), .CK(clk), .Q(ram[517]) );
  DFF_X1 ram_reg_32__4_ ( .D(n13036), .CK(clk), .Q(ram[516]) );
  DFF_X1 ram_reg_32__3_ ( .D(n13035), .CK(clk), .Q(ram[515]) );
  DFF_X1 ram_reg_32__2_ ( .D(n13034), .CK(clk), .Q(ram[514]) );
  DFF_X1 ram_reg_32__1_ ( .D(n13033), .CK(clk), .Q(ram[513]) );
  DFF_X1 ram_reg_32__0_ ( .D(n13032), .CK(clk), .Q(ram[512]) );
  DFF_X1 ram_reg_31__15_ ( .D(n13064), .CK(clk), .Q(ram[511]) );
  DFF_X1 ram_reg_31__14_ ( .D(n13063), .CK(clk), .Q(ram[510]) );
  DFF_X1 ram_reg_31__13_ ( .D(n13062), .CK(clk), .Q(ram[509]) );
  DFF_X1 ram_reg_31__12_ ( .D(n13061), .CK(clk), .Q(ram[508]) );
  DFF_X1 ram_reg_31__11_ ( .D(n13060), .CK(clk), .Q(ram[507]) );
  DFF_X1 ram_reg_31__10_ ( .D(n13059), .CK(clk), .Q(ram[506]) );
  DFF_X1 ram_reg_31__9_ ( .D(n13058), .CK(clk), .Q(ram[505]) );
  DFF_X1 ram_reg_31__8_ ( .D(n13057), .CK(clk), .Q(ram[504]) );
  DFF_X1 ram_reg_31__7_ ( .D(n13056), .CK(clk), .Q(ram[503]) );
  DFF_X1 ram_reg_31__6_ ( .D(n13055), .CK(clk), .Q(ram[502]) );
  DFF_X1 ram_reg_31__5_ ( .D(n13054), .CK(clk), .Q(ram[501]) );
  DFF_X1 ram_reg_31__4_ ( .D(n13053), .CK(clk), .Q(ram[500]) );
  DFF_X1 ram_reg_31__3_ ( .D(n13052), .CK(clk), .Q(ram[499]) );
  DFF_X1 ram_reg_31__2_ ( .D(n13051), .CK(clk), .Q(ram[498]) );
  DFF_X1 ram_reg_31__1_ ( .D(n13050), .CK(clk), .Q(ram[497]) );
  DFF_X1 ram_reg_31__0_ ( .D(n13049), .CK(clk), .Q(ram[496]) );
  DFF_X1 ram_reg_30__15_ ( .D(n13081), .CK(clk), .Q(ram[495]) );
  DFF_X1 ram_reg_30__14_ ( .D(n13080), .CK(clk), .Q(ram[494]) );
  DFF_X1 ram_reg_30__13_ ( .D(n13079), .CK(clk), .Q(ram[493]) );
  DFF_X1 ram_reg_30__12_ ( .D(n13078), .CK(clk), .Q(ram[492]) );
  DFF_X1 ram_reg_30__11_ ( .D(n13077), .CK(clk), .Q(ram[491]) );
  DFF_X1 ram_reg_30__10_ ( .D(n13076), .CK(clk), .Q(ram[490]) );
  DFF_X1 ram_reg_30__9_ ( .D(n13075), .CK(clk), .Q(ram[489]) );
  DFF_X1 ram_reg_30__8_ ( .D(n13074), .CK(clk), .Q(ram[488]) );
  DFF_X1 ram_reg_30__7_ ( .D(n13073), .CK(clk), .Q(ram[487]) );
  DFF_X1 ram_reg_30__6_ ( .D(n13072), .CK(clk), .Q(ram[486]) );
  DFF_X1 ram_reg_30__5_ ( .D(n13071), .CK(clk), .Q(ram[485]) );
  DFF_X1 ram_reg_30__4_ ( .D(n13070), .CK(clk), .Q(ram[484]) );
  DFF_X1 ram_reg_30__3_ ( .D(n13069), .CK(clk), .Q(ram[483]) );
  DFF_X1 ram_reg_30__2_ ( .D(n13068), .CK(clk), .Q(ram[482]) );
  DFF_X1 ram_reg_30__1_ ( .D(n13067), .CK(clk), .Q(ram[481]) );
  DFF_X1 ram_reg_30__0_ ( .D(n13066), .CK(clk), .Q(ram[480]) );
  DFF_X1 ram_reg_29__15_ ( .D(n13098), .CK(clk), .Q(ram[479]) );
  DFF_X1 ram_reg_29__14_ ( .D(n13097), .CK(clk), .Q(ram[478]) );
  DFF_X1 ram_reg_29__13_ ( .D(n13096), .CK(clk), .Q(ram[477]) );
  DFF_X1 ram_reg_29__12_ ( .D(n13095), .CK(clk), .Q(ram[476]) );
  DFF_X1 ram_reg_29__11_ ( .D(n13094), .CK(clk), .Q(ram[475]) );
  DFF_X1 ram_reg_29__10_ ( .D(n13093), .CK(clk), .Q(ram[474]) );
  DFF_X1 ram_reg_29__9_ ( .D(n13092), .CK(clk), .Q(ram[473]) );
  DFF_X1 ram_reg_29__8_ ( .D(n13091), .CK(clk), .Q(ram[472]) );
  DFF_X1 ram_reg_29__7_ ( .D(n13090), .CK(clk), .Q(ram[471]) );
  DFF_X1 ram_reg_29__6_ ( .D(n13089), .CK(clk), .Q(ram[470]) );
  DFF_X1 ram_reg_29__5_ ( .D(n13088), .CK(clk), .Q(ram[469]) );
  DFF_X1 ram_reg_29__4_ ( .D(n13087), .CK(clk), .Q(ram[468]) );
  DFF_X1 ram_reg_29__3_ ( .D(n13086), .CK(clk), .Q(ram[467]) );
  DFF_X1 ram_reg_29__2_ ( .D(n13085), .CK(clk), .Q(ram[466]) );
  DFF_X1 ram_reg_29__1_ ( .D(n13084), .CK(clk), .Q(ram[465]) );
  DFF_X1 ram_reg_29__0_ ( .D(n13083), .CK(clk), .Q(ram[464]) );
  DFF_X1 ram_reg_28__15_ ( .D(n13115), .CK(clk), .Q(ram[463]) );
  DFF_X1 ram_reg_28__14_ ( .D(n13114), .CK(clk), .Q(ram[462]) );
  DFF_X1 ram_reg_28__13_ ( .D(n13113), .CK(clk), .Q(ram[461]) );
  DFF_X1 ram_reg_28__12_ ( .D(n13112), .CK(clk), .Q(ram[460]) );
  DFF_X1 ram_reg_28__11_ ( .D(n13111), .CK(clk), .Q(ram[459]) );
  DFF_X1 ram_reg_28__10_ ( .D(n13110), .CK(clk), .Q(ram[458]) );
  DFF_X1 ram_reg_28__9_ ( .D(n13109), .CK(clk), .Q(ram[457]) );
  DFF_X1 ram_reg_28__8_ ( .D(n13108), .CK(clk), .Q(ram[456]) );
  DFF_X1 ram_reg_28__7_ ( .D(n13107), .CK(clk), .Q(ram[455]) );
  DFF_X1 ram_reg_28__6_ ( .D(n13106), .CK(clk), .Q(ram[454]) );
  DFF_X1 ram_reg_28__5_ ( .D(n13105), .CK(clk), .Q(ram[453]) );
  DFF_X1 ram_reg_28__4_ ( .D(n13104), .CK(clk), .Q(ram[452]) );
  DFF_X1 ram_reg_28__3_ ( .D(n13103), .CK(clk), .Q(ram[451]) );
  DFF_X1 ram_reg_28__2_ ( .D(n13102), .CK(clk), .Q(ram[450]) );
  DFF_X1 ram_reg_28__1_ ( .D(n13101), .CK(clk), .Q(ram[449]) );
  DFF_X1 ram_reg_28__0_ ( .D(n13100), .CK(clk), .Q(ram[448]) );
  DFF_X1 ram_reg_27__15_ ( .D(n13132), .CK(clk), .Q(ram[447]) );
  DFF_X1 ram_reg_27__14_ ( .D(n13131), .CK(clk), .Q(ram[446]) );
  DFF_X1 ram_reg_27__13_ ( .D(n13130), .CK(clk), .Q(ram[445]) );
  DFF_X1 ram_reg_27__12_ ( .D(n13129), .CK(clk), .Q(ram[444]) );
  DFF_X1 ram_reg_27__11_ ( .D(n13128), .CK(clk), .Q(ram[443]) );
  DFF_X1 ram_reg_27__10_ ( .D(n13127), .CK(clk), .Q(ram[442]) );
  DFF_X1 ram_reg_27__9_ ( .D(n13126), .CK(clk), .Q(ram[441]) );
  DFF_X1 ram_reg_27__8_ ( .D(n13125), .CK(clk), .Q(ram[440]) );
  DFF_X1 ram_reg_27__7_ ( .D(n13124), .CK(clk), .Q(ram[439]) );
  DFF_X1 ram_reg_27__6_ ( .D(n13123), .CK(clk), .Q(ram[438]) );
  DFF_X1 ram_reg_27__5_ ( .D(n13122), .CK(clk), .Q(ram[437]) );
  DFF_X1 ram_reg_27__4_ ( .D(n13121), .CK(clk), .Q(ram[436]) );
  DFF_X1 ram_reg_27__3_ ( .D(n13120), .CK(clk), .Q(ram[435]) );
  DFF_X1 ram_reg_27__2_ ( .D(n13119), .CK(clk), .Q(ram[434]) );
  DFF_X1 ram_reg_27__1_ ( .D(n13118), .CK(clk), .Q(ram[433]) );
  DFF_X1 ram_reg_27__0_ ( .D(n13117), .CK(clk), .Q(ram[432]) );
  DFF_X1 ram_reg_26__15_ ( .D(n13149), .CK(clk), .Q(ram[431]) );
  DFF_X1 ram_reg_26__14_ ( .D(n13148), .CK(clk), .Q(ram[430]) );
  DFF_X1 ram_reg_26__13_ ( .D(n13147), .CK(clk), .Q(ram[429]) );
  DFF_X1 ram_reg_26__12_ ( .D(n13146), .CK(clk), .Q(ram[428]) );
  DFF_X1 ram_reg_26__11_ ( .D(n13145), .CK(clk), .Q(ram[427]) );
  DFF_X1 ram_reg_26__10_ ( .D(n13144), .CK(clk), .Q(ram[426]) );
  DFF_X1 ram_reg_26__9_ ( .D(n13143), .CK(clk), .Q(ram[425]) );
  DFF_X1 ram_reg_26__8_ ( .D(n13142), .CK(clk), .Q(ram[424]) );
  DFF_X1 ram_reg_26__7_ ( .D(n13141), .CK(clk), .Q(ram[423]) );
  DFF_X1 ram_reg_26__6_ ( .D(n13140), .CK(clk), .Q(ram[422]) );
  DFF_X1 ram_reg_26__5_ ( .D(n13139), .CK(clk), .Q(ram[421]) );
  DFF_X1 ram_reg_26__4_ ( .D(n13138), .CK(clk), .Q(ram[420]) );
  DFF_X1 ram_reg_26__3_ ( .D(n13137), .CK(clk), .Q(ram[419]) );
  DFF_X1 ram_reg_26__2_ ( .D(n13136), .CK(clk), .Q(ram[418]) );
  DFF_X1 ram_reg_26__1_ ( .D(n13135), .CK(clk), .Q(ram[417]) );
  DFF_X1 ram_reg_26__0_ ( .D(n13134), .CK(clk), .Q(ram[416]) );
  DFF_X1 ram_reg_25__15_ ( .D(n13166), .CK(clk), .Q(ram[415]) );
  DFF_X1 ram_reg_25__14_ ( .D(n13165), .CK(clk), .Q(ram[414]) );
  DFF_X1 ram_reg_25__13_ ( .D(n13164), .CK(clk), .Q(ram[413]) );
  DFF_X1 ram_reg_25__12_ ( .D(n13163), .CK(clk), .Q(ram[412]) );
  DFF_X1 ram_reg_25__11_ ( .D(n13162), .CK(clk), .Q(ram[411]) );
  DFF_X1 ram_reg_25__10_ ( .D(n13161), .CK(clk), .Q(ram[410]) );
  DFF_X1 ram_reg_25__9_ ( .D(n13160), .CK(clk), .Q(ram[409]) );
  DFF_X1 ram_reg_25__8_ ( .D(n13159), .CK(clk), .Q(ram[408]) );
  DFF_X1 ram_reg_25__7_ ( .D(n13158), .CK(clk), .Q(ram[407]) );
  DFF_X1 ram_reg_25__6_ ( .D(n13157), .CK(clk), .Q(ram[406]) );
  DFF_X1 ram_reg_25__5_ ( .D(n13156), .CK(clk), .Q(ram[405]) );
  DFF_X1 ram_reg_25__4_ ( .D(n13155), .CK(clk), .Q(ram[404]) );
  DFF_X1 ram_reg_25__3_ ( .D(n13154), .CK(clk), .Q(ram[403]) );
  DFF_X1 ram_reg_25__2_ ( .D(n13153), .CK(clk), .Q(ram[402]) );
  DFF_X1 ram_reg_25__1_ ( .D(n13152), .CK(clk), .Q(ram[401]) );
  DFF_X1 ram_reg_25__0_ ( .D(n13151), .CK(clk), .Q(ram[400]) );
  DFF_X1 ram_reg_24__15_ ( .D(n13183), .CK(clk), .Q(ram[399]) );
  DFF_X1 ram_reg_24__14_ ( .D(n13182), .CK(clk), .Q(ram[398]) );
  DFF_X1 ram_reg_24__13_ ( .D(n13181), .CK(clk), .Q(ram[397]) );
  DFF_X1 ram_reg_24__12_ ( .D(n13180), .CK(clk), .Q(ram[396]) );
  DFF_X1 ram_reg_24__11_ ( .D(n13179), .CK(clk), .Q(ram[395]) );
  DFF_X1 ram_reg_24__10_ ( .D(n13178), .CK(clk), .Q(ram[394]) );
  DFF_X1 ram_reg_24__9_ ( .D(n13177), .CK(clk), .Q(ram[393]) );
  DFF_X1 ram_reg_24__8_ ( .D(n13176), .CK(clk), .Q(ram[392]) );
  DFF_X1 ram_reg_24__7_ ( .D(n13175), .CK(clk), .Q(ram[391]) );
  DFF_X1 ram_reg_24__6_ ( .D(n13174), .CK(clk), .Q(ram[390]) );
  DFF_X1 ram_reg_24__5_ ( .D(n13173), .CK(clk), .Q(ram[389]) );
  DFF_X1 ram_reg_24__4_ ( .D(n13172), .CK(clk), .Q(ram[388]) );
  DFF_X1 ram_reg_24__3_ ( .D(n13171), .CK(clk), .Q(ram[387]) );
  DFF_X1 ram_reg_24__2_ ( .D(n13170), .CK(clk), .Q(ram[386]) );
  DFF_X1 ram_reg_24__1_ ( .D(n13169), .CK(clk), .Q(ram[385]) );
  DFF_X1 ram_reg_24__0_ ( .D(n13168), .CK(clk), .Q(ram[384]) );
  DFF_X1 ram_reg_23__15_ ( .D(n13200), .CK(clk), .Q(ram[383]) );
  DFF_X1 ram_reg_23__14_ ( .D(n13199), .CK(clk), .Q(ram[382]) );
  DFF_X1 ram_reg_23__13_ ( .D(n13198), .CK(clk), .Q(ram[381]) );
  DFF_X1 ram_reg_23__12_ ( .D(n13197), .CK(clk), .Q(ram[380]) );
  DFF_X1 ram_reg_23__11_ ( .D(n13196), .CK(clk), .Q(ram[379]) );
  DFF_X1 ram_reg_23__10_ ( .D(n13195), .CK(clk), .Q(ram[378]) );
  DFF_X1 ram_reg_23__9_ ( .D(n13194), .CK(clk), .Q(ram[377]) );
  DFF_X1 ram_reg_23__8_ ( .D(n13193), .CK(clk), .Q(ram[376]) );
  DFF_X1 ram_reg_23__7_ ( .D(n13192), .CK(clk), .Q(ram[375]) );
  DFF_X1 ram_reg_23__6_ ( .D(n13191), .CK(clk), .Q(ram[374]) );
  DFF_X1 ram_reg_23__5_ ( .D(n13190), .CK(clk), .Q(ram[373]) );
  DFF_X1 ram_reg_23__4_ ( .D(n13189), .CK(clk), .Q(ram[372]) );
  DFF_X1 ram_reg_23__3_ ( .D(n13188), .CK(clk), .Q(ram[371]) );
  DFF_X1 ram_reg_23__2_ ( .D(n13187), .CK(clk), .Q(ram[370]) );
  DFF_X1 ram_reg_23__1_ ( .D(n13186), .CK(clk), .Q(ram[369]) );
  DFF_X1 ram_reg_23__0_ ( .D(n13185), .CK(clk), .Q(ram[368]) );
  DFF_X1 ram_reg_22__15_ ( .D(n13217), .CK(clk), .Q(ram[367]) );
  DFF_X1 ram_reg_22__14_ ( .D(n13216), .CK(clk), .Q(ram[366]) );
  DFF_X1 ram_reg_22__13_ ( .D(n13215), .CK(clk), .Q(ram[365]) );
  DFF_X1 ram_reg_22__12_ ( .D(n13214), .CK(clk), .Q(ram[364]) );
  DFF_X1 ram_reg_22__11_ ( .D(n13213), .CK(clk), .Q(ram[363]) );
  DFF_X1 ram_reg_22__10_ ( .D(n13212), .CK(clk), .Q(ram[362]) );
  DFF_X1 ram_reg_22__9_ ( .D(n13211), .CK(clk), .Q(ram[361]) );
  DFF_X1 ram_reg_22__8_ ( .D(n13210), .CK(clk), .Q(ram[360]) );
  DFF_X1 ram_reg_22__7_ ( .D(n13209), .CK(clk), .Q(ram[359]) );
  DFF_X1 ram_reg_22__6_ ( .D(n13208), .CK(clk), .Q(ram[358]) );
  DFF_X1 ram_reg_22__5_ ( .D(n13207), .CK(clk), .Q(ram[357]) );
  DFF_X1 ram_reg_22__4_ ( .D(n13206), .CK(clk), .Q(ram[356]) );
  DFF_X1 ram_reg_22__3_ ( .D(n13205), .CK(clk), .Q(ram[355]) );
  DFF_X1 ram_reg_22__2_ ( .D(n13204), .CK(clk), .Q(ram[354]) );
  DFF_X1 ram_reg_22__1_ ( .D(n13203), .CK(clk), .Q(ram[353]) );
  DFF_X1 ram_reg_22__0_ ( .D(n13202), .CK(clk), .Q(ram[352]) );
  DFF_X1 ram_reg_21__15_ ( .D(n13234), .CK(clk), .Q(ram[351]) );
  DFF_X1 ram_reg_21__14_ ( .D(n13233), .CK(clk), .Q(ram[350]) );
  DFF_X1 ram_reg_21__13_ ( .D(n13232), .CK(clk), .Q(ram[349]) );
  DFF_X1 ram_reg_21__12_ ( .D(n13231), .CK(clk), .Q(ram[348]) );
  DFF_X1 ram_reg_21__11_ ( .D(n13230), .CK(clk), .Q(ram[347]) );
  DFF_X1 ram_reg_21__10_ ( .D(n13229), .CK(clk), .Q(ram[346]) );
  DFF_X1 ram_reg_21__9_ ( .D(n13228), .CK(clk), .Q(ram[345]) );
  DFF_X1 ram_reg_21__8_ ( .D(n13227), .CK(clk), .Q(ram[344]) );
  DFF_X1 ram_reg_21__7_ ( .D(n13226), .CK(clk), .Q(ram[343]) );
  DFF_X1 ram_reg_21__6_ ( .D(n13225), .CK(clk), .Q(ram[342]) );
  DFF_X1 ram_reg_21__5_ ( .D(n13224), .CK(clk), .Q(ram[341]) );
  DFF_X1 ram_reg_21__4_ ( .D(n13223), .CK(clk), .Q(ram[340]) );
  DFF_X1 ram_reg_21__3_ ( .D(n13222), .CK(clk), .Q(ram[339]) );
  DFF_X1 ram_reg_21__2_ ( .D(n13221), .CK(clk), .Q(ram[338]) );
  DFF_X1 ram_reg_21__1_ ( .D(n13220), .CK(clk), .Q(ram[337]) );
  DFF_X1 ram_reg_21__0_ ( .D(n13219), .CK(clk), .Q(ram[336]) );
  DFF_X1 ram_reg_20__15_ ( .D(n13251), .CK(clk), .Q(ram[335]) );
  DFF_X1 ram_reg_20__14_ ( .D(n13250), .CK(clk), .Q(ram[334]) );
  DFF_X1 ram_reg_20__13_ ( .D(n13249), .CK(clk), .Q(ram[333]) );
  DFF_X1 ram_reg_20__12_ ( .D(n13248), .CK(clk), .Q(ram[332]) );
  DFF_X1 ram_reg_20__11_ ( .D(n13247), .CK(clk), .Q(ram[331]) );
  DFF_X1 ram_reg_20__10_ ( .D(n13246), .CK(clk), .Q(ram[330]) );
  DFF_X1 ram_reg_20__9_ ( .D(n13245), .CK(clk), .Q(ram[329]) );
  DFF_X1 ram_reg_20__8_ ( .D(n13244), .CK(clk), .Q(ram[328]) );
  DFF_X1 ram_reg_20__7_ ( .D(n13243), .CK(clk), .Q(ram[327]) );
  DFF_X1 ram_reg_20__6_ ( .D(n13242), .CK(clk), .Q(ram[326]) );
  DFF_X1 ram_reg_20__5_ ( .D(n13241), .CK(clk), .Q(ram[325]) );
  DFF_X1 ram_reg_20__4_ ( .D(n13240), .CK(clk), .Q(ram[324]) );
  DFF_X1 ram_reg_20__3_ ( .D(n13239), .CK(clk), .Q(ram[323]) );
  DFF_X1 ram_reg_20__2_ ( .D(n13238), .CK(clk), .Q(ram[322]) );
  DFF_X1 ram_reg_20__1_ ( .D(n13237), .CK(clk), .Q(ram[321]) );
  DFF_X1 ram_reg_20__0_ ( .D(n13236), .CK(clk), .Q(ram[320]) );
  DFF_X1 ram_reg_19__15_ ( .D(n13268), .CK(clk), .Q(ram[319]) );
  DFF_X1 ram_reg_19__14_ ( .D(n13267), .CK(clk), .Q(ram[318]) );
  DFF_X1 ram_reg_19__13_ ( .D(n13266), .CK(clk), .Q(ram[317]) );
  DFF_X1 ram_reg_19__12_ ( .D(n13265), .CK(clk), .Q(ram[316]) );
  DFF_X1 ram_reg_19__11_ ( .D(n13264), .CK(clk), .Q(ram[315]) );
  DFF_X1 ram_reg_19__10_ ( .D(n13263), .CK(clk), .Q(ram[314]) );
  DFF_X1 ram_reg_19__9_ ( .D(n13262), .CK(clk), .Q(ram[313]) );
  DFF_X1 ram_reg_19__8_ ( .D(n13261), .CK(clk), .Q(ram[312]) );
  DFF_X1 ram_reg_19__7_ ( .D(n13260), .CK(clk), .Q(ram[311]) );
  DFF_X1 ram_reg_19__6_ ( .D(n13259), .CK(clk), .Q(ram[310]) );
  DFF_X1 ram_reg_19__5_ ( .D(n13258), .CK(clk), .Q(ram[309]) );
  DFF_X1 ram_reg_19__4_ ( .D(n13257), .CK(clk), .Q(ram[308]) );
  DFF_X1 ram_reg_19__3_ ( .D(n13256), .CK(clk), .Q(ram[307]) );
  DFF_X1 ram_reg_19__2_ ( .D(n13255), .CK(clk), .Q(ram[306]) );
  DFF_X1 ram_reg_19__1_ ( .D(n13254), .CK(clk), .Q(ram[305]) );
  DFF_X1 ram_reg_19__0_ ( .D(n13253), .CK(clk), .Q(ram[304]) );
  DFF_X1 ram_reg_18__15_ ( .D(n13285), .CK(clk), .Q(ram[303]) );
  DFF_X1 ram_reg_18__14_ ( .D(n13284), .CK(clk), .Q(ram[302]) );
  DFF_X1 ram_reg_18__13_ ( .D(n13283), .CK(clk), .Q(ram[301]) );
  DFF_X1 ram_reg_18__12_ ( .D(n13282), .CK(clk), .Q(ram[300]) );
  DFF_X1 ram_reg_18__11_ ( .D(n13281), .CK(clk), .Q(ram[299]) );
  DFF_X1 ram_reg_18__10_ ( .D(n13280), .CK(clk), .Q(ram[298]) );
  DFF_X1 ram_reg_18__9_ ( .D(n13279), .CK(clk), .Q(ram[297]) );
  DFF_X1 ram_reg_18__8_ ( .D(n13278), .CK(clk), .Q(ram[296]) );
  DFF_X1 ram_reg_18__7_ ( .D(n13277), .CK(clk), .Q(ram[295]) );
  DFF_X1 ram_reg_18__6_ ( .D(n13276), .CK(clk), .Q(ram[294]) );
  DFF_X1 ram_reg_18__5_ ( .D(n13275), .CK(clk), .Q(ram[293]) );
  DFF_X1 ram_reg_18__4_ ( .D(n13274), .CK(clk), .Q(ram[292]) );
  DFF_X1 ram_reg_18__3_ ( .D(n13273), .CK(clk), .Q(ram[291]) );
  DFF_X1 ram_reg_18__2_ ( .D(n13272), .CK(clk), .Q(ram[290]) );
  DFF_X1 ram_reg_18__1_ ( .D(n13271), .CK(clk), .Q(ram[289]) );
  DFF_X1 ram_reg_18__0_ ( .D(n13270), .CK(clk), .Q(ram[288]) );
  DFF_X1 ram_reg_17__15_ ( .D(n13302), .CK(clk), .Q(ram[287]) );
  DFF_X1 ram_reg_17__14_ ( .D(n13301), .CK(clk), .Q(ram[286]) );
  DFF_X1 ram_reg_17__13_ ( .D(n13300), .CK(clk), .Q(ram[285]) );
  DFF_X1 ram_reg_17__12_ ( .D(n13299), .CK(clk), .Q(ram[284]) );
  DFF_X1 ram_reg_17__11_ ( .D(n13298), .CK(clk), .Q(ram[283]) );
  DFF_X1 ram_reg_17__10_ ( .D(n13297), .CK(clk), .Q(ram[282]) );
  DFF_X1 ram_reg_17__9_ ( .D(n13296), .CK(clk), .Q(ram[281]) );
  DFF_X1 ram_reg_17__8_ ( .D(n13295), .CK(clk), .Q(ram[280]) );
  DFF_X1 ram_reg_17__7_ ( .D(n13294), .CK(clk), .Q(ram[279]) );
  DFF_X1 ram_reg_17__6_ ( .D(n13293), .CK(clk), .Q(ram[278]) );
  DFF_X1 ram_reg_17__5_ ( .D(n13292), .CK(clk), .Q(ram[277]) );
  DFF_X1 ram_reg_17__4_ ( .D(n13291), .CK(clk), .Q(ram[276]) );
  DFF_X1 ram_reg_17__3_ ( .D(n13290), .CK(clk), .Q(ram[275]) );
  DFF_X1 ram_reg_17__2_ ( .D(n13289), .CK(clk), .Q(ram[274]) );
  DFF_X1 ram_reg_17__1_ ( .D(n13288), .CK(clk), .Q(ram[273]) );
  DFF_X1 ram_reg_17__0_ ( .D(n13287), .CK(clk), .Q(ram[272]) );
  DFF_X1 ram_reg_16__15_ ( .D(n13319), .CK(clk), .Q(ram[271]) );
  DFF_X1 ram_reg_16__14_ ( .D(n13318), .CK(clk), .Q(ram[270]) );
  DFF_X1 ram_reg_16__13_ ( .D(n13317), .CK(clk), .Q(ram[269]) );
  DFF_X1 ram_reg_16__12_ ( .D(n13316), .CK(clk), .Q(ram[268]) );
  DFF_X1 ram_reg_16__11_ ( .D(n13315), .CK(clk), .Q(ram[267]) );
  DFF_X1 ram_reg_16__10_ ( .D(n13314), .CK(clk), .Q(ram[266]) );
  DFF_X1 ram_reg_16__9_ ( .D(n13313), .CK(clk), .Q(ram[265]) );
  DFF_X1 ram_reg_16__8_ ( .D(n13312), .CK(clk), .Q(ram[264]) );
  DFF_X1 ram_reg_16__7_ ( .D(n13311), .CK(clk), .Q(ram[263]) );
  DFF_X1 ram_reg_16__6_ ( .D(n13310), .CK(clk), .Q(ram[262]) );
  DFF_X1 ram_reg_16__5_ ( .D(n13309), .CK(clk), .Q(ram[261]) );
  DFF_X1 ram_reg_16__4_ ( .D(n13308), .CK(clk), .Q(ram[260]) );
  DFF_X1 ram_reg_16__3_ ( .D(n13307), .CK(clk), .Q(ram[259]) );
  DFF_X1 ram_reg_16__2_ ( .D(n13306), .CK(clk), .Q(ram[258]) );
  DFF_X1 ram_reg_16__1_ ( .D(n13305), .CK(clk), .Q(ram[257]) );
  DFF_X1 ram_reg_16__0_ ( .D(n13304), .CK(clk), .Q(ram[256]) );
  DFF_X1 ram_reg_15__15_ ( .D(n13336), .CK(clk), .Q(ram[255]) );
  DFF_X1 ram_reg_15__14_ ( .D(n13335), .CK(clk), .Q(ram[254]) );
  DFF_X1 ram_reg_15__13_ ( .D(n13334), .CK(clk), .Q(ram[253]) );
  DFF_X1 ram_reg_15__12_ ( .D(n13333), .CK(clk), .Q(ram[252]) );
  DFF_X1 ram_reg_15__11_ ( .D(n13332), .CK(clk), .Q(ram[251]) );
  DFF_X1 ram_reg_15__10_ ( .D(n13331), .CK(clk), .Q(ram[250]) );
  DFF_X1 ram_reg_15__9_ ( .D(n13330), .CK(clk), .Q(ram[249]) );
  DFF_X1 ram_reg_15__8_ ( .D(n13329), .CK(clk), .Q(ram[248]) );
  DFF_X1 ram_reg_15__7_ ( .D(n13328), .CK(clk), .Q(ram[247]) );
  DFF_X1 ram_reg_15__6_ ( .D(n13327), .CK(clk), .Q(ram[246]) );
  DFF_X1 ram_reg_15__5_ ( .D(n13326), .CK(clk), .Q(ram[245]) );
  DFF_X1 ram_reg_15__4_ ( .D(n13325), .CK(clk), .Q(ram[244]) );
  DFF_X1 ram_reg_15__3_ ( .D(n13324), .CK(clk), .Q(ram[243]) );
  DFF_X1 ram_reg_15__2_ ( .D(n13323), .CK(clk), .Q(ram[242]) );
  DFF_X1 ram_reg_15__1_ ( .D(n13322), .CK(clk), .Q(ram[241]) );
  DFF_X1 ram_reg_15__0_ ( .D(n13321), .CK(clk), .Q(ram[240]) );
  DFF_X1 ram_reg_14__15_ ( .D(n13353), .CK(clk), .Q(ram[239]) );
  DFF_X1 ram_reg_14__14_ ( .D(n13352), .CK(clk), .Q(ram[238]) );
  DFF_X1 ram_reg_14__13_ ( .D(n13351), .CK(clk), .Q(ram[237]) );
  DFF_X1 ram_reg_14__12_ ( .D(n13350), .CK(clk), .Q(ram[236]) );
  DFF_X1 ram_reg_14__11_ ( .D(n13349), .CK(clk), .Q(ram[235]) );
  DFF_X1 ram_reg_14__10_ ( .D(n13348), .CK(clk), .Q(ram[234]) );
  DFF_X1 ram_reg_14__9_ ( .D(n13347), .CK(clk), .Q(ram[233]) );
  DFF_X1 ram_reg_14__8_ ( .D(n13346), .CK(clk), .Q(ram[232]) );
  DFF_X1 ram_reg_14__7_ ( .D(n13345), .CK(clk), .Q(ram[231]) );
  DFF_X1 ram_reg_14__6_ ( .D(n13344), .CK(clk), .Q(ram[230]) );
  DFF_X1 ram_reg_14__5_ ( .D(n13343), .CK(clk), .Q(ram[229]) );
  DFF_X1 ram_reg_14__4_ ( .D(n13342), .CK(clk), .Q(ram[228]) );
  DFF_X1 ram_reg_14__3_ ( .D(n13341), .CK(clk), .Q(ram[227]) );
  DFF_X1 ram_reg_14__2_ ( .D(n13340), .CK(clk), .Q(ram[226]) );
  DFF_X1 ram_reg_14__1_ ( .D(n13339), .CK(clk), .Q(ram[225]) );
  DFF_X1 ram_reg_14__0_ ( .D(n13338), .CK(clk), .Q(ram[224]) );
  DFF_X1 ram_reg_13__15_ ( .D(n13370), .CK(clk), .Q(ram[223]) );
  DFF_X1 ram_reg_13__14_ ( .D(n13369), .CK(clk), .Q(ram[222]) );
  DFF_X1 ram_reg_13__13_ ( .D(n13368), .CK(clk), .Q(ram[221]) );
  DFF_X1 ram_reg_13__12_ ( .D(n13367), .CK(clk), .Q(ram[220]) );
  DFF_X1 ram_reg_13__11_ ( .D(n13366), .CK(clk), .Q(ram[219]) );
  DFF_X1 ram_reg_13__10_ ( .D(n13365), .CK(clk), .Q(ram[218]) );
  DFF_X1 ram_reg_13__9_ ( .D(n13364), .CK(clk), .Q(ram[217]) );
  DFF_X1 ram_reg_13__8_ ( .D(n13363), .CK(clk), .Q(ram[216]) );
  DFF_X1 ram_reg_13__7_ ( .D(n13362), .CK(clk), .Q(ram[215]) );
  DFF_X1 ram_reg_13__6_ ( .D(n13361), .CK(clk), .Q(ram[214]) );
  DFF_X1 ram_reg_13__5_ ( .D(n13360), .CK(clk), .Q(ram[213]) );
  DFF_X1 ram_reg_13__4_ ( .D(n13359), .CK(clk), .Q(ram[212]) );
  DFF_X1 ram_reg_13__3_ ( .D(n13358), .CK(clk), .Q(ram[211]) );
  DFF_X1 ram_reg_13__2_ ( .D(n13357), .CK(clk), .Q(ram[210]) );
  DFF_X1 ram_reg_13__1_ ( .D(n13356), .CK(clk), .Q(ram[209]) );
  DFF_X1 ram_reg_13__0_ ( .D(n13355), .CK(clk), .Q(ram[208]) );
  DFF_X1 ram_reg_12__15_ ( .D(n13387), .CK(clk), .Q(ram[207]) );
  DFF_X1 ram_reg_12__14_ ( .D(n13386), .CK(clk), .Q(ram[206]) );
  DFF_X1 ram_reg_12__13_ ( .D(n13385), .CK(clk), .Q(ram[205]) );
  DFF_X1 ram_reg_12__12_ ( .D(n13384), .CK(clk), .Q(ram[204]) );
  DFF_X1 ram_reg_12__11_ ( .D(n13383), .CK(clk), .Q(ram[203]) );
  DFF_X1 ram_reg_12__10_ ( .D(n13382), .CK(clk), .Q(ram[202]) );
  DFF_X1 ram_reg_12__9_ ( .D(n13381), .CK(clk), .Q(ram[201]) );
  DFF_X1 ram_reg_12__8_ ( .D(n13380), .CK(clk), .Q(ram[200]) );
  DFF_X1 ram_reg_12__7_ ( .D(n13379), .CK(clk), .Q(ram[199]) );
  DFF_X1 ram_reg_12__6_ ( .D(n13378), .CK(clk), .Q(ram[198]) );
  DFF_X1 ram_reg_12__5_ ( .D(n13377), .CK(clk), .Q(ram[197]) );
  DFF_X1 ram_reg_12__4_ ( .D(n13376), .CK(clk), .Q(ram[196]) );
  DFF_X1 ram_reg_12__3_ ( .D(n13375), .CK(clk), .Q(ram[195]) );
  DFF_X1 ram_reg_12__2_ ( .D(n13374), .CK(clk), .Q(ram[194]) );
  DFF_X1 ram_reg_12__1_ ( .D(n13373), .CK(clk), .Q(ram[193]) );
  DFF_X1 ram_reg_12__0_ ( .D(n13372), .CK(clk), .Q(ram[192]) );
  DFF_X1 ram_reg_11__15_ ( .D(n13404), .CK(clk), .Q(ram[191]) );
  DFF_X1 ram_reg_11__14_ ( .D(n13403), .CK(clk), .Q(ram[190]) );
  DFF_X1 ram_reg_11__13_ ( .D(n13402), .CK(clk), .Q(ram[189]) );
  DFF_X1 ram_reg_11__12_ ( .D(n13401), .CK(clk), .Q(ram[188]) );
  DFF_X1 ram_reg_11__11_ ( .D(n13400), .CK(clk), .Q(ram[187]) );
  DFF_X1 ram_reg_11__10_ ( .D(n13399), .CK(clk), .Q(ram[186]) );
  DFF_X1 ram_reg_11__9_ ( .D(n13398), .CK(clk), .Q(ram[185]) );
  DFF_X1 ram_reg_11__8_ ( .D(n13397), .CK(clk), .Q(ram[184]) );
  DFF_X1 ram_reg_11__7_ ( .D(n13396), .CK(clk), .Q(ram[183]) );
  DFF_X1 ram_reg_11__6_ ( .D(n13395), .CK(clk), .Q(ram[182]) );
  DFF_X1 ram_reg_11__5_ ( .D(n13394), .CK(clk), .Q(ram[181]) );
  DFF_X1 ram_reg_11__4_ ( .D(n13393), .CK(clk), .Q(ram[180]) );
  DFF_X1 ram_reg_11__3_ ( .D(n13392), .CK(clk), .Q(ram[179]) );
  DFF_X1 ram_reg_11__2_ ( .D(n13391), .CK(clk), .Q(ram[178]) );
  DFF_X1 ram_reg_11__1_ ( .D(n13390), .CK(clk), .Q(ram[177]) );
  DFF_X1 ram_reg_11__0_ ( .D(n13389), .CK(clk), .Q(ram[176]) );
  DFF_X1 ram_reg_10__15_ ( .D(n13421), .CK(clk), .Q(ram[175]) );
  DFF_X1 ram_reg_10__14_ ( .D(n13420), .CK(clk), .Q(ram[174]) );
  DFF_X1 ram_reg_10__13_ ( .D(n13419), .CK(clk), .Q(ram[173]) );
  DFF_X1 ram_reg_10__12_ ( .D(n13418), .CK(clk), .Q(ram[172]) );
  DFF_X1 ram_reg_10__11_ ( .D(n13417), .CK(clk), .Q(ram[171]) );
  DFF_X1 ram_reg_10__10_ ( .D(n13416), .CK(clk), .Q(ram[170]) );
  DFF_X1 ram_reg_10__9_ ( .D(n13415), .CK(clk), .Q(ram[169]) );
  DFF_X1 ram_reg_10__8_ ( .D(n13414), .CK(clk), .Q(ram[168]) );
  DFF_X1 ram_reg_10__7_ ( .D(n13413), .CK(clk), .Q(ram[167]) );
  DFF_X1 ram_reg_10__6_ ( .D(n13412), .CK(clk), .Q(ram[166]) );
  DFF_X1 ram_reg_10__5_ ( .D(n13411), .CK(clk), .Q(ram[165]) );
  DFF_X1 ram_reg_10__4_ ( .D(n13410), .CK(clk), .Q(ram[164]) );
  DFF_X1 ram_reg_10__3_ ( .D(n13409), .CK(clk), .Q(ram[163]) );
  DFF_X1 ram_reg_10__2_ ( .D(n13408), .CK(clk), .Q(ram[162]) );
  DFF_X1 ram_reg_10__1_ ( .D(n13407), .CK(clk), .Q(ram[161]) );
  DFF_X1 ram_reg_10__0_ ( .D(n13406), .CK(clk), .Q(ram[160]) );
  DFF_X1 ram_reg_9__15_ ( .D(n13438), .CK(clk), .Q(ram[159]) );
  DFF_X1 ram_reg_9__14_ ( .D(n13437), .CK(clk), .Q(ram[158]) );
  DFF_X1 ram_reg_9__13_ ( .D(n13436), .CK(clk), .Q(ram[157]) );
  DFF_X1 ram_reg_9__12_ ( .D(n13435), .CK(clk), .Q(ram[156]) );
  DFF_X1 ram_reg_9__11_ ( .D(n13434), .CK(clk), .Q(ram[155]) );
  DFF_X1 ram_reg_9__10_ ( .D(n13433), .CK(clk), .Q(ram[154]) );
  DFF_X1 ram_reg_9__9_ ( .D(n13432), .CK(clk), .Q(ram[153]) );
  DFF_X1 ram_reg_9__8_ ( .D(n13431), .CK(clk), .Q(ram[152]) );
  DFF_X1 ram_reg_9__7_ ( .D(n13430), .CK(clk), .Q(ram[151]) );
  DFF_X1 ram_reg_9__6_ ( .D(n13429), .CK(clk), .Q(ram[150]) );
  DFF_X1 ram_reg_9__5_ ( .D(n13428), .CK(clk), .Q(ram[149]) );
  DFF_X1 ram_reg_9__4_ ( .D(n13427), .CK(clk), .Q(ram[148]) );
  DFF_X1 ram_reg_9__3_ ( .D(n13426), .CK(clk), .Q(ram[147]) );
  DFF_X1 ram_reg_9__2_ ( .D(n13425), .CK(clk), .Q(ram[146]) );
  DFF_X1 ram_reg_9__1_ ( .D(n13424), .CK(clk), .Q(ram[145]) );
  DFF_X1 ram_reg_9__0_ ( .D(n13423), .CK(clk), .Q(ram[144]) );
  DFF_X1 ram_reg_8__15_ ( .D(n13455), .CK(clk), .Q(ram[143]) );
  DFF_X1 ram_reg_8__14_ ( .D(n13454), .CK(clk), .Q(ram[142]) );
  DFF_X1 ram_reg_8__13_ ( .D(n13453), .CK(clk), .Q(ram[141]) );
  DFF_X1 ram_reg_8__12_ ( .D(n13452), .CK(clk), .Q(ram[140]) );
  DFF_X1 ram_reg_8__11_ ( .D(n13451), .CK(clk), .Q(ram[139]) );
  DFF_X1 ram_reg_8__10_ ( .D(n13450), .CK(clk), .Q(ram[138]) );
  DFF_X1 ram_reg_8__9_ ( .D(n13449), .CK(clk), .Q(ram[137]) );
  DFF_X1 ram_reg_8__8_ ( .D(n13448), .CK(clk), .Q(ram[136]) );
  DFF_X1 ram_reg_8__7_ ( .D(n13447), .CK(clk), .Q(ram[135]) );
  DFF_X1 ram_reg_8__6_ ( .D(n13446), .CK(clk), .Q(ram[134]) );
  DFF_X1 ram_reg_8__5_ ( .D(n13445), .CK(clk), .Q(ram[133]) );
  DFF_X1 ram_reg_8__4_ ( .D(n13444), .CK(clk), .Q(ram[132]) );
  DFF_X1 ram_reg_8__3_ ( .D(n13443), .CK(clk), .Q(ram[131]) );
  DFF_X1 ram_reg_8__2_ ( .D(n13442), .CK(clk), .Q(ram[130]) );
  DFF_X1 ram_reg_8__1_ ( .D(n13441), .CK(clk), .Q(ram[129]) );
  DFF_X1 ram_reg_8__0_ ( .D(n13440), .CK(clk), .Q(ram[128]) );
  DFF_X1 ram_reg_7__15_ ( .D(n13472), .CK(clk), .Q(ram[127]) );
  DFF_X1 ram_reg_7__14_ ( .D(n13471), .CK(clk), .Q(ram[126]) );
  DFF_X1 ram_reg_7__13_ ( .D(n13470), .CK(clk), .Q(ram[125]) );
  DFF_X1 ram_reg_7__12_ ( .D(n13469), .CK(clk), .Q(ram[124]) );
  DFF_X1 ram_reg_7__11_ ( .D(n13468), .CK(clk), .Q(ram[123]) );
  DFF_X1 ram_reg_7__10_ ( .D(n13467), .CK(clk), .Q(ram[122]) );
  DFF_X1 ram_reg_7__9_ ( .D(n13466), .CK(clk), .Q(ram[121]) );
  DFF_X1 ram_reg_7__8_ ( .D(n13465), .CK(clk), .Q(ram[120]) );
  DFF_X1 ram_reg_7__7_ ( .D(n13464), .CK(clk), .Q(ram[119]) );
  DFF_X1 ram_reg_7__6_ ( .D(n13463), .CK(clk), .Q(ram[118]) );
  DFF_X1 ram_reg_7__5_ ( .D(n13462), .CK(clk), .Q(ram[117]) );
  DFF_X1 ram_reg_7__4_ ( .D(n13461), .CK(clk), .Q(ram[116]) );
  DFF_X1 ram_reg_7__3_ ( .D(n13460), .CK(clk), .Q(ram[115]) );
  DFF_X1 ram_reg_7__2_ ( .D(n13459), .CK(clk), .Q(ram[114]) );
  DFF_X1 ram_reg_7__1_ ( .D(n13458), .CK(clk), .Q(ram[113]) );
  DFF_X1 ram_reg_7__0_ ( .D(n13457), .CK(clk), .Q(ram[112]) );
  DFF_X1 ram_reg_6__15_ ( .D(n13489), .CK(clk), .Q(ram[111]) );
  DFF_X1 ram_reg_6__14_ ( .D(n13488), .CK(clk), .Q(ram[110]) );
  DFF_X1 ram_reg_6__13_ ( .D(n13487), .CK(clk), .Q(ram[109]) );
  DFF_X1 ram_reg_6__12_ ( .D(n13486), .CK(clk), .Q(ram[108]) );
  DFF_X1 ram_reg_6__11_ ( .D(n13485), .CK(clk), .Q(ram[107]) );
  DFF_X1 ram_reg_6__10_ ( .D(n13484), .CK(clk), .Q(ram[106]) );
  DFF_X1 ram_reg_6__9_ ( .D(n13483), .CK(clk), .Q(ram[105]) );
  DFF_X1 ram_reg_6__8_ ( .D(n13482), .CK(clk), .Q(ram[104]) );
  DFF_X1 ram_reg_6__7_ ( .D(n13481), .CK(clk), .Q(ram[103]) );
  DFF_X1 ram_reg_6__6_ ( .D(n13480), .CK(clk), .Q(ram[102]) );
  DFF_X1 ram_reg_6__5_ ( .D(n13479), .CK(clk), .Q(ram[101]) );
  DFF_X1 ram_reg_6__4_ ( .D(n13478), .CK(clk), .Q(ram[100]) );
  DFF_X1 ram_reg_6__3_ ( .D(n13477), .CK(clk), .Q(ram[99]) );
  DFF_X1 ram_reg_6__2_ ( .D(n13476), .CK(clk), .Q(ram[98]) );
  DFF_X1 ram_reg_6__1_ ( .D(n13475), .CK(clk), .Q(ram[97]) );
  DFF_X1 ram_reg_6__0_ ( .D(n13474), .CK(clk), .Q(ram[96]) );
  DFF_X1 ram_reg_5__15_ ( .D(n13506), .CK(clk), .Q(ram[95]) );
  DFF_X1 ram_reg_5__14_ ( .D(n13505), .CK(clk), .Q(ram[94]) );
  DFF_X1 ram_reg_5__13_ ( .D(n13504), .CK(clk), .Q(ram[93]) );
  DFF_X1 ram_reg_5__12_ ( .D(n13503), .CK(clk), .Q(ram[92]) );
  DFF_X1 ram_reg_5__11_ ( .D(n13502), .CK(clk), .Q(ram[91]) );
  DFF_X1 ram_reg_5__10_ ( .D(n13501), .CK(clk), .Q(ram[90]) );
  DFF_X1 ram_reg_5__9_ ( .D(n13500), .CK(clk), .Q(ram[89]) );
  DFF_X1 ram_reg_5__8_ ( .D(n13499), .CK(clk), .Q(ram[88]) );
  DFF_X1 ram_reg_5__7_ ( .D(n13498), .CK(clk), .Q(ram[87]) );
  DFF_X1 ram_reg_5__6_ ( .D(n13497), .CK(clk), .Q(ram[86]) );
  DFF_X1 ram_reg_5__5_ ( .D(n13496), .CK(clk), .Q(ram[85]) );
  DFF_X1 ram_reg_5__4_ ( .D(n13495), .CK(clk), .Q(ram[84]) );
  DFF_X1 ram_reg_5__3_ ( .D(n13494), .CK(clk), .Q(ram[83]) );
  DFF_X1 ram_reg_5__2_ ( .D(n13493), .CK(clk), .Q(ram[82]) );
  DFF_X1 ram_reg_5__1_ ( .D(n13492), .CK(clk), .Q(ram[81]) );
  DFF_X1 ram_reg_5__0_ ( .D(n13491), .CK(clk), .Q(ram[80]) );
  DFF_X1 ram_reg_4__15_ ( .D(n13523), .CK(clk), .Q(ram[79]) );
  DFF_X1 ram_reg_4__14_ ( .D(n13522), .CK(clk), .Q(ram[78]) );
  DFF_X1 ram_reg_4__13_ ( .D(n13521), .CK(clk), .Q(ram[77]) );
  DFF_X1 ram_reg_4__12_ ( .D(n13520), .CK(clk), .Q(ram[76]) );
  DFF_X1 ram_reg_4__11_ ( .D(n13519), .CK(clk), .Q(ram[75]) );
  DFF_X1 ram_reg_4__10_ ( .D(n13518), .CK(clk), .Q(ram[74]) );
  DFF_X1 ram_reg_4__9_ ( .D(n13517), .CK(clk), .Q(ram[73]) );
  DFF_X1 ram_reg_4__8_ ( .D(n13516), .CK(clk), .Q(ram[72]) );
  DFF_X1 ram_reg_4__7_ ( .D(n13515), .CK(clk), .Q(ram[71]) );
  DFF_X1 ram_reg_4__6_ ( .D(n13514), .CK(clk), .Q(ram[70]) );
  DFF_X1 ram_reg_4__5_ ( .D(n13513), .CK(clk), .Q(ram[69]) );
  DFF_X1 ram_reg_4__4_ ( .D(n13512), .CK(clk), .Q(ram[68]) );
  DFF_X1 ram_reg_4__3_ ( .D(n13511), .CK(clk), .Q(ram[67]) );
  DFF_X1 ram_reg_4__2_ ( .D(n13510), .CK(clk), .Q(ram[66]) );
  DFF_X1 ram_reg_4__1_ ( .D(n13509), .CK(clk), .Q(ram[65]) );
  DFF_X1 ram_reg_4__0_ ( .D(n13508), .CK(clk), .Q(ram[64]) );
  DFF_X1 ram_reg_3__15_ ( .D(n13540), .CK(clk), .Q(ram[63]) );
  DFF_X1 ram_reg_3__14_ ( .D(n13539), .CK(clk), .Q(ram[62]) );
  DFF_X1 ram_reg_3__13_ ( .D(n13538), .CK(clk), .Q(ram[61]) );
  DFF_X1 ram_reg_3__12_ ( .D(n13537), .CK(clk), .Q(ram[60]) );
  DFF_X1 ram_reg_3__11_ ( .D(n13536), .CK(clk), .Q(ram[59]) );
  DFF_X1 ram_reg_3__10_ ( .D(n13535), .CK(clk), .Q(ram[58]) );
  DFF_X1 ram_reg_3__9_ ( .D(n13534), .CK(clk), .Q(ram[57]) );
  DFF_X1 ram_reg_3__8_ ( .D(n13533), .CK(clk), .Q(ram[56]) );
  DFF_X1 ram_reg_3__7_ ( .D(n13532), .CK(clk), .Q(ram[55]) );
  DFF_X1 ram_reg_3__6_ ( .D(n13531), .CK(clk), .Q(ram[54]) );
  DFF_X1 ram_reg_3__5_ ( .D(n13530), .CK(clk), .Q(ram[53]) );
  DFF_X1 ram_reg_3__4_ ( .D(n13529), .CK(clk), .Q(ram[52]) );
  DFF_X1 ram_reg_3__3_ ( .D(n13528), .CK(clk), .Q(ram[51]) );
  DFF_X1 ram_reg_3__2_ ( .D(n13527), .CK(clk), .Q(ram[50]) );
  DFF_X1 ram_reg_3__1_ ( .D(n13526), .CK(clk), .Q(ram[49]) );
  DFF_X1 ram_reg_3__0_ ( .D(n13525), .CK(clk), .Q(ram[48]) );
  DFF_X1 ram_reg_2__15_ ( .D(n13557), .CK(clk), .Q(ram[47]) );
  DFF_X1 ram_reg_2__14_ ( .D(n13556), .CK(clk), .Q(ram[46]) );
  DFF_X1 ram_reg_2__13_ ( .D(n13555), .CK(clk), .Q(ram[45]) );
  DFF_X1 ram_reg_2__12_ ( .D(n13554), .CK(clk), .Q(ram[44]) );
  DFF_X1 ram_reg_2__11_ ( .D(n13553), .CK(clk), .Q(ram[43]) );
  DFF_X1 ram_reg_2__10_ ( .D(n13552), .CK(clk), .Q(ram[42]) );
  DFF_X1 ram_reg_2__9_ ( .D(n13551), .CK(clk), .Q(ram[41]) );
  DFF_X1 ram_reg_2__8_ ( .D(n13550), .CK(clk), .Q(ram[40]) );
  DFF_X1 ram_reg_2__7_ ( .D(n13549), .CK(clk), .Q(ram[39]) );
  DFF_X1 ram_reg_2__6_ ( .D(n13548), .CK(clk), .Q(ram[38]) );
  DFF_X1 ram_reg_2__5_ ( .D(n13547), .CK(clk), .Q(ram[37]) );
  DFF_X1 ram_reg_2__4_ ( .D(n13546), .CK(clk), .Q(ram[36]) );
  DFF_X1 ram_reg_2__3_ ( .D(n13545), .CK(clk), .Q(ram[35]) );
  DFF_X1 ram_reg_2__2_ ( .D(n13544), .CK(clk), .Q(ram[34]) );
  DFF_X1 ram_reg_2__1_ ( .D(n13543), .CK(clk), .Q(ram[33]) );
  DFF_X1 ram_reg_2__0_ ( .D(n13542), .CK(clk), .Q(ram[32]) );
  DFF_X1 ram_reg_1__15_ ( .D(n13574), .CK(clk), .Q(ram[31]) );
  DFF_X1 ram_reg_1__14_ ( .D(n13573), .CK(clk), .Q(ram[30]) );
  DFF_X1 ram_reg_1__13_ ( .D(n13572), .CK(clk), .Q(ram[29]) );
  DFF_X1 ram_reg_1__12_ ( .D(n13571), .CK(clk), .Q(ram[28]) );
  DFF_X1 ram_reg_1__11_ ( .D(n13570), .CK(clk), .Q(ram[27]) );
  DFF_X1 ram_reg_1__10_ ( .D(n13569), .CK(clk), .Q(ram[26]) );
  DFF_X1 ram_reg_1__9_ ( .D(n13568), .CK(clk), .Q(ram[25]) );
  DFF_X1 ram_reg_1__8_ ( .D(n13567), .CK(clk), .Q(ram[24]) );
  DFF_X1 ram_reg_1__7_ ( .D(n13566), .CK(clk), .Q(ram[23]) );
  DFF_X1 ram_reg_1__6_ ( .D(n13565), .CK(clk), .Q(ram[22]) );
  DFF_X1 ram_reg_1__5_ ( .D(n13564), .CK(clk), .Q(ram[21]) );
  DFF_X1 ram_reg_1__4_ ( .D(n13563), .CK(clk), .Q(ram[20]) );
  DFF_X1 ram_reg_1__3_ ( .D(n13562), .CK(clk), .Q(ram[19]) );
  DFF_X1 ram_reg_1__2_ ( .D(n13561), .CK(clk), .Q(ram[18]) );
  DFF_X1 ram_reg_1__1_ ( .D(n13560), .CK(clk), .Q(ram[17]) );
  DFF_X1 ram_reg_1__0_ ( .D(n13559), .CK(clk), .Q(ram[16]) );
  DFF_X1 ram_reg_0__15_ ( .D(n13591), .CK(clk), .Q(ram[15]) );
  DFF_X1 ram_reg_0__14_ ( .D(n13590), .CK(clk), .Q(ram[14]) );
  DFF_X1 ram_reg_0__13_ ( .D(n13589), .CK(clk), .Q(ram[13]) );
  DFF_X1 ram_reg_0__12_ ( .D(n13588), .CK(clk), .Q(ram[12]) );
  DFF_X1 ram_reg_0__11_ ( .D(n13587), .CK(clk), .Q(ram[11]) );
  DFF_X1 ram_reg_0__10_ ( .D(n13586), .CK(clk), .Q(ram[10]) );
  DFF_X1 ram_reg_0__9_ ( .D(n13585), .CK(clk), .Q(ram[9]) );
  DFF_X1 ram_reg_0__8_ ( .D(n13584), .CK(clk), .Q(ram[8]) );
  DFF_X1 ram_reg_0__7_ ( .D(n13583), .CK(clk), .Q(ram[7]) );
  DFF_X1 ram_reg_0__6_ ( .D(n13582), .CK(clk), .Q(ram[6]) );
  DFF_X1 ram_reg_0__5_ ( .D(n13581), .CK(clk), .Q(ram[5]) );
  DFF_X1 ram_reg_0__4_ ( .D(n13580), .CK(clk), .Q(ram[4]) );
  DFF_X1 ram_reg_0__3_ ( .D(n13579), .CK(clk), .Q(ram[3]) );
  DFF_X1 ram_reg_0__2_ ( .D(n13578), .CK(clk), .Q(ram[2]) );
  DFF_X1 ram_reg_0__1_ ( .D(n13577), .CK(clk), .Q(ram[1]) );
  DFF_X1 ram_reg_0__0_ ( .D(n13576), .CK(clk), .Q(ram[0]) );
  BUF_X1 U2 ( .A(n4278), .Z(n4283) );
  BUF_X1 U3 ( .A(n4278), .Z(n4282) );
  BUF_X1 U4 ( .A(n4278), .Z(n4281) );
  BUF_X1 U5 ( .A(n4278), .Z(n4280) );
  BUF_X1 U6 ( .A(n4277), .Z(n4293) );
  BUF_X1 U7 ( .A(n4277), .Z(n4292) );
  BUF_X1 U8 ( .A(n4277), .Z(n4291) );
  BUF_X1 U9 ( .A(n4277), .Z(n4290) );
  BUF_X1 U10 ( .A(n4276), .Z(n4304) );
  BUF_X1 U11 ( .A(n4276), .Z(n4303) );
  BUF_X1 U12 ( .A(n4276), .Z(n4302) );
  BUF_X1 U13 ( .A(n4276), .Z(n4301) );
  BUF_X1 U14 ( .A(n4275), .Z(n4315) );
  BUF_X1 U15 ( .A(n4275), .Z(n4314) );
  BUF_X1 U16 ( .A(n4275), .Z(n4313) );
  BUF_X1 U17 ( .A(n4275), .Z(n4312) );
  BUF_X1 U18 ( .A(n4274), .Z(n4326) );
  BUF_X1 U19 ( .A(n4274), .Z(n4325) );
  BUF_X1 U20 ( .A(n4274), .Z(n4324) );
  BUF_X1 U21 ( .A(n4274), .Z(n4323) );
  BUF_X1 U22 ( .A(n4273), .Z(n4337) );
  BUF_X1 U23 ( .A(n4273), .Z(n4336) );
  BUF_X1 U24 ( .A(n4273), .Z(n4335) );
  BUF_X1 U25 ( .A(n4273), .Z(n4334) );
  BUF_X1 U26 ( .A(n4272), .Z(n4348) );
  BUF_X1 U27 ( .A(n4272), .Z(n4347) );
  BUF_X1 U28 ( .A(n4272), .Z(n4346) );
  BUF_X1 U29 ( .A(n4272), .Z(n4345) );
  BUF_X1 U30 ( .A(n4271), .Z(n8759) );
  BUF_X1 U31 ( .A(n4271), .Z(n8758) );
  BUF_X1 U32 ( .A(n4271), .Z(n8757) );
  BUF_X1 U33 ( .A(n4271), .Z(n4356) );
  BUF_X1 U34 ( .A(n4270), .Z(n8770) );
  BUF_X1 U35 ( .A(n4270), .Z(n8769) );
  BUF_X1 U36 ( .A(n4270), .Z(n8768) );
  BUF_X1 U37 ( .A(n4270), .Z(n8767) );
  BUF_X1 U38 ( .A(n4269), .Z(n8781) );
  BUF_X1 U39 ( .A(n4269), .Z(n8780) );
  BUF_X1 U40 ( .A(n4269), .Z(n8779) );
  BUF_X1 U41 ( .A(n4269), .Z(n8778) );
  BUF_X1 U42 ( .A(n4268), .Z(n8792) );
  BUF_X1 U43 ( .A(n4268), .Z(n8791) );
  BUF_X1 U44 ( .A(n4268), .Z(n8790) );
  BUF_X1 U45 ( .A(n4268), .Z(n8789) );
  BUF_X1 U46 ( .A(n4267), .Z(n8803) );
  BUF_X1 U47 ( .A(n4267), .Z(n8802) );
  BUF_X1 U48 ( .A(n4267), .Z(n8801) );
  BUF_X1 U49 ( .A(n4267), .Z(n8800) );
  BUF_X1 U50 ( .A(n4266), .Z(n8814) );
  BUF_X1 U51 ( .A(n4266), .Z(n8813) );
  BUF_X1 U52 ( .A(n4266), .Z(n8812) );
  BUF_X1 U53 ( .A(n4266), .Z(n8811) );
  BUF_X1 U54 ( .A(n4265), .Z(n8825) );
  BUF_X1 U55 ( .A(n4265), .Z(n8824) );
  BUF_X1 U56 ( .A(n4265), .Z(n8823) );
  BUF_X1 U57 ( .A(n4265), .Z(n8822) );
  BUF_X1 U58 ( .A(n4264), .Z(n8836) );
  BUF_X1 U59 ( .A(n4264), .Z(n8835) );
  BUF_X1 U60 ( .A(n4264), .Z(n8834) );
  BUF_X1 U61 ( .A(n4264), .Z(n8833) );
  BUF_X1 U62 ( .A(n4263), .Z(n8849) );
  BUF_X1 U63 ( .A(n4263), .Z(n8848) );
  BUF_X1 U64 ( .A(n4263), .Z(n8847) );
  BUF_X1 U65 ( .A(n4263), .Z(n8846) );
  BUF_X1 U66 ( .A(n4263), .Z(n8845) );
  BUF_X1 U67 ( .A(n4263), .Z(n8844) );
  BUF_X1 U68 ( .A(n4119), .Z(n4122) );
  BUF_X1 U69 ( .A(n4119), .Z(n4121) );
  BUF_X1 U70 ( .A(n4119), .Z(n4124) );
  BUF_X1 U71 ( .A(n4119), .Z(n4123) );
  BUF_X1 U72 ( .A(n4118), .Z(n4127) );
  BUF_X1 U73 ( .A(n4118), .Z(n4126) );
  BUF_X1 U74 ( .A(n4118), .Z(n4125) );
  BUF_X1 U75 ( .A(n4117), .Z(n4130) );
  BUF_X1 U76 ( .A(n4118), .Z(n4129) );
  BUF_X1 U77 ( .A(n4118), .Z(n4128) );
  BUF_X1 U78 ( .A(n4117), .Z(n4132) );
  BUF_X1 U79 ( .A(n4117), .Z(n4131) );
  BUF_X1 U80 ( .A(n4116), .Z(n4135) );
  BUF_X1 U81 ( .A(n4117), .Z(n4134) );
  BUF_X1 U82 ( .A(n4117), .Z(n4133) );
  BUF_X1 U83 ( .A(n4116), .Z(n4138) );
  BUF_X1 U84 ( .A(n4116), .Z(n4137) );
  BUF_X1 U85 ( .A(n4116), .Z(n4136) );
  BUF_X1 U86 ( .A(n4115), .Z(n4140) );
  BUF_X1 U87 ( .A(n4116), .Z(n4139) );
  BUF_X1 U88 ( .A(n4115), .Z(n4143) );
  BUF_X1 U89 ( .A(n4115), .Z(n4142) );
  BUF_X1 U90 ( .A(n4115), .Z(n4141) );
  BUF_X1 U91 ( .A(n4114), .Z(n4146) );
  BUF_X1 U92 ( .A(n4114), .Z(n4145) );
  BUF_X1 U93 ( .A(n4115), .Z(n4144) );
  BUF_X1 U94 ( .A(n4114), .Z(n4148) );
  BUF_X1 U95 ( .A(n4114), .Z(n4147) );
  BUF_X1 U96 ( .A(n4113), .Z(n4151) );
  BUF_X1 U97 ( .A(n4113), .Z(n4150) );
  BUF_X1 U98 ( .A(n4114), .Z(n4149) );
  BUF_X1 U99 ( .A(n4113), .Z(n4154) );
  BUF_X1 U100 ( .A(n4113), .Z(n4153) );
  BUF_X1 U101 ( .A(n4113), .Z(n4152) );
  BUF_X1 U102 ( .A(n4112), .Z(n4156) );
  BUF_X1 U103 ( .A(n4112), .Z(n4155) );
  BUF_X1 U104 ( .A(n4112), .Z(n4159) );
  BUF_X1 U105 ( .A(n4112), .Z(n4158) );
  BUF_X1 U106 ( .A(n4112), .Z(n4157) );
  BUF_X1 U107 ( .A(n4111), .Z(n4162) );
  BUF_X1 U108 ( .A(n4111), .Z(n4161) );
  BUF_X1 U109 ( .A(n4111), .Z(n4160) );
  BUF_X1 U110 ( .A(n4163), .Z(n4111) );
  BUF_X1 U111 ( .A(n4165), .Z(n4118) );
  BUF_X1 U112 ( .A(n4165), .Z(n4117) );
  BUF_X1 U113 ( .A(n4164), .Z(n4116) );
  BUF_X1 U114 ( .A(n4164), .Z(n4115) );
  BUF_X1 U115 ( .A(n4164), .Z(n4114) );
  BUF_X1 U116 ( .A(n4163), .Z(n4113) );
  BUF_X1 U117 ( .A(n4163), .Z(n4112) );
  BUF_X1 U118 ( .A(n4165), .Z(n4119) );
  BUF_X1 U119 ( .A(n8851), .Z(n4278) );
  BUF_X1 U120 ( .A(n8851), .Z(n4277) );
  BUF_X1 U121 ( .A(n8851), .Z(n4276) );
  BUF_X1 U122 ( .A(n8851), .Z(n4275) );
  BUF_X1 U123 ( .A(n8851), .Z(n4274) );
  BUF_X1 U124 ( .A(n8851), .Z(n4273) );
  BUF_X1 U125 ( .A(n8851), .Z(n4272) );
  BUF_X1 U126 ( .A(n8851), .Z(n4271) );
  BUF_X1 U127 ( .A(n8851), .Z(n4270) );
  BUF_X1 U128 ( .A(n8851), .Z(n4269) );
  BUF_X1 U129 ( .A(n8851), .Z(n4268) );
  BUF_X1 U130 ( .A(n8851), .Z(n4267) );
  BUF_X1 U131 ( .A(n8850), .Z(n4266) );
  BUF_X1 U132 ( .A(n8850), .Z(n4265) );
  BUF_X1 U133 ( .A(n8850), .Z(n4264) );
  BUF_X1 U134 ( .A(n8850), .Z(n4263) );
  BUF_X1 U135 ( .A(n9238), .Z(n4077) );
  BUF_X1 U136 ( .A(n9238), .Z(n4078) );
  BUF_X1 U137 ( .A(n9238), .Z(n4079) );
  BUF_X1 U138 ( .A(n9238), .Z(n4080) );
  BUF_X1 U139 ( .A(mem_access_addr[8]), .Z(n4066) );
  BUF_X1 U140 ( .A(mem_access_addr[8]), .Z(n4067) );
  BUF_X1 U141 ( .A(n4173), .Z(n4178) );
  BUF_X1 U142 ( .A(n4173), .Z(n4177) );
  BUF_X1 U143 ( .A(n4173), .Z(n4176) );
  BUF_X1 U144 ( .A(n4173), .Z(n4175) );
  BUF_X1 U145 ( .A(n4172), .Z(n4188) );
  BUF_X1 U146 ( .A(n4172), .Z(n4187) );
  BUF_X1 U147 ( .A(n4172), .Z(n4186) );
  BUF_X1 U148 ( .A(n4172), .Z(n4185) );
  BUF_X1 U149 ( .A(n4171), .Z(n4199) );
  BUF_X1 U150 ( .A(n4171), .Z(n4198) );
  BUF_X1 U151 ( .A(n4171), .Z(n4197) );
  BUF_X1 U152 ( .A(n4171), .Z(n4196) );
  BUF_X1 U153 ( .A(n4170), .Z(n4210) );
  BUF_X1 U154 ( .A(n4170), .Z(n4209) );
  BUF_X1 U155 ( .A(n4170), .Z(n4208) );
  BUF_X1 U156 ( .A(n4170), .Z(n4207) );
  BUF_X1 U157 ( .A(n4169), .Z(n4221) );
  BUF_X1 U158 ( .A(n4169), .Z(n4220) );
  BUF_X1 U159 ( .A(n4169), .Z(n4219) );
  BUF_X1 U160 ( .A(n4169), .Z(n4218) );
  BUF_X1 U161 ( .A(n4168), .Z(n4232) );
  BUF_X1 U162 ( .A(n4168), .Z(n4231) );
  BUF_X1 U163 ( .A(n4168), .Z(n4230) );
  BUF_X1 U164 ( .A(n4168), .Z(n4229) );
  BUF_X1 U165 ( .A(n4167), .Z(n4243) );
  BUF_X1 U166 ( .A(n4167), .Z(n4242) );
  BUF_X1 U167 ( .A(n4167), .Z(n4241) );
  BUF_X1 U168 ( .A(n4167), .Z(n4240) );
  BUF_X1 U169 ( .A(n4166), .Z(n4253) );
  BUF_X1 U170 ( .A(n4166), .Z(n4252) );
  BUF_X1 U171 ( .A(n4166), .Z(n4251) );
  BUF_X1 U172 ( .A(n4166), .Z(n4254) );
  BUF_X1 U173 ( .A(mem_access_addr[8]), .Z(n4065) );
  BUF_X1 U174 ( .A(mem_access_addr[4]), .Z(n4165) );
  BUF_X1 U175 ( .A(mem_access_addr[4]), .Z(n4164) );
  BUF_X1 U176 ( .A(mem_access_addr[4]), .Z(n4163) );
  BUF_X1 U177 ( .A(mem_access_addr[2]), .Z(n8851) );
  BUF_X1 U178 ( .A(mem_access_addr[2]), .Z(n8850) );
  AND2_X1 U179 ( .A1(n8494), .A2(n8495), .ZN(n4374) );
  AND2_X1 U180 ( .A1(n8513), .A2(n8494), .ZN(n4393) );
  AND2_X1 U181 ( .A1(n8567), .A2(n8495), .ZN(n4447) );
  AND2_X1 U182 ( .A1(n8567), .A2(n8513), .ZN(n4465) );
  AND2_X1 U183 ( .A1(n8567), .A2(n8531), .ZN(n4483) );
  AND2_X1 U184 ( .A1(n8567), .A2(n8549), .ZN(n4501) );
  AND2_X1 U185 ( .A1(n8531), .A2(n8494), .ZN(n4411) );
  AND2_X1 U186 ( .A1(n8549), .A2(n8494), .ZN(n4429) );
  AND2_X1 U187 ( .A1(n8636), .A2(n8495), .ZN(n4519) );
  AND2_X1 U188 ( .A1(n8636), .A2(n8513), .ZN(n4537) );
  AND2_X1 U189 ( .A1(n8705), .A2(n8495), .ZN(n4591) );
  AND2_X1 U190 ( .A1(n8705), .A2(n8513), .ZN(n4609) );
  AND2_X1 U191 ( .A1(n8636), .A2(n8531), .ZN(n4555) );
  AND2_X1 U192 ( .A1(n8636), .A2(n8549), .ZN(n4573) );
  AND2_X1 U193 ( .A1(n8705), .A2(n8531), .ZN(n4627) );
  AND2_X1 U194 ( .A1(n8705), .A2(n8549), .ZN(n4645) );
  BUF_X1 U195 ( .A(n4109), .Z(n4088) );
  BUF_X1 U196 ( .A(n4109), .Z(n4089) );
  BUF_X1 U197 ( .A(n4109), .Z(n4090) );
  BUF_X1 U198 ( .A(n4109), .Z(n4091) );
  BUF_X1 U199 ( .A(n4110), .Z(n4098) );
  BUF_X1 U200 ( .A(n4110), .Z(n4100) );
  BUF_X1 U201 ( .A(n4110), .Z(n4099) );
  BUF_X1 U202 ( .A(n4110), .Z(n4101) );
  BUF_X1 U203 ( .A(n4074), .Z(n4069) );
  BUF_X1 U204 ( .A(n4074), .Z(n4070) );
  BUF_X1 U205 ( .A(n4075), .Z(n4071) );
  BUF_X1 U206 ( .A(n4075), .Z(n4072) );
  BUF_X1 U207 ( .A(n4075), .Z(n4073) );
  BUF_X1 U208 ( .A(n4262), .Z(n4173) );
  BUF_X1 U209 ( .A(n4262), .Z(n4172) );
  BUF_X1 U210 ( .A(n4262), .Z(n4171) );
  BUF_X1 U211 ( .A(n4261), .Z(n4170) );
  BUF_X1 U212 ( .A(n4261), .Z(n4169) );
  BUF_X1 U213 ( .A(n4261), .Z(n4168) );
  BUF_X1 U214 ( .A(n4260), .Z(n4167) );
  BUF_X1 U215 ( .A(n4260), .Z(n4166) );
  INV_X1 U216 ( .A(n4358), .ZN(n13592) );
  INV_X1 U217 ( .A(n4649), .ZN(n13320) );
  INV_X1 U218 ( .A(n4667), .ZN(n13303) );
  INV_X1 U219 ( .A(n4684), .ZN(n13286) );
  INV_X1 U220 ( .A(n4701), .ZN(n13269) );
  INV_X1 U221 ( .A(n4718), .ZN(n13252) );
  INV_X1 U222 ( .A(n4735), .ZN(n13235) );
  INV_X1 U223 ( .A(n4752), .ZN(n13218) );
  INV_X1 U224 ( .A(n4769), .ZN(n13201) );
  INV_X1 U225 ( .A(n4786), .ZN(n13184) );
  INV_X1 U226 ( .A(n4803), .ZN(n13167) );
  INV_X1 U227 ( .A(n4820), .ZN(n13150) );
  INV_X1 U228 ( .A(n4837), .ZN(n13133) );
  INV_X1 U229 ( .A(n4854), .ZN(n13116) );
  INV_X1 U230 ( .A(n4871), .ZN(n13099) );
  INV_X1 U231 ( .A(n4888), .ZN(n13082) );
  INV_X1 U232 ( .A(n4905), .ZN(n13065) );
  INV_X1 U233 ( .A(n4923), .ZN(n13048) );
  INV_X1 U234 ( .A(n4941), .ZN(n13031) );
  INV_X1 U235 ( .A(n4958), .ZN(n13014) );
  INV_X1 U236 ( .A(n4975), .ZN(n12997) );
  INV_X1 U237 ( .A(n4992), .ZN(n12980) );
  INV_X1 U238 ( .A(n5009), .ZN(n12963) );
  INV_X1 U239 ( .A(n5026), .ZN(n12946) );
  INV_X1 U240 ( .A(n5043), .ZN(n12929) );
  INV_X1 U241 ( .A(n5060), .ZN(n12912) );
  INV_X1 U242 ( .A(n5077), .ZN(n12895) );
  INV_X1 U243 ( .A(n5094), .ZN(n12878) );
  INV_X1 U244 ( .A(n5111), .ZN(n12861) );
  INV_X1 U245 ( .A(n5128), .ZN(n12844) );
  INV_X1 U246 ( .A(n5145), .ZN(n12827) );
  INV_X1 U247 ( .A(n5162), .ZN(n12810) );
  INV_X1 U248 ( .A(n5179), .ZN(n12793) );
  INV_X1 U249 ( .A(n5197), .ZN(n12776) );
  INV_X1 U250 ( .A(n5215), .ZN(n12759) );
  INV_X1 U251 ( .A(n5232), .ZN(n12742) );
  INV_X1 U252 ( .A(n5249), .ZN(n12725) );
  INV_X1 U253 ( .A(n5266), .ZN(n12708) );
  INV_X1 U254 ( .A(n5283), .ZN(n12691) );
  INV_X1 U255 ( .A(n5300), .ZN(n12674) );
  INV_X1 U256 ( .A(n5317), .ZN(n12657) );
  INV_X1 U257 ( .A(n5334), .ZN(n12640) );
  INV_X1 U258 ( .A(n5351), .ZN(n12623) );
  INV_X1 U259 ( .A(n5368), .ZN(n12606) );
  INV_X1 U260 ( .A(n5385), .ZN(n12589) );
  INV_X1 U261 ( .A(n5402), .ZN(n12572) );
  INV_X1 U262 ( .A(n5419), .ZN(n12555) );
  INV_X1 U263 ( .A(n5436), .ZN(n12538) );
  INV_X1 U264 ( .A(n5453), .ZN(n12521) );
  INV_X1 U265 ( .A(n5471), .ZN(n12504) );
  INV_X1 U266 ( .A(n5489), .ZN(n12487) );
  INV_X1 U267 ( .A(n5506), .ZN(n12470) );
  INV_X1 U268 ( .A(n5523), .ZN(n12453) );
  INV_X1 U269 ( .A(n5540), .ZN(n12436) );
  INV_X1 U270 ( .A(n5557), .ZN(n12419) );
  INV_X1 U271 ( .A(n5574), .ZN(n12402) );
  INV_X1 U272 ( .A(n5591), .ZN(n12385) );
  INV_X1 U273 ( .A(n5608), .ZN(n12368) );
  INV_X1 U274 ( .A(n5625), .ZN(n12351) );
  INV_X1 U275 ( .A(n5642), .ZN(n12334) );
  INV_X1 U276 ( .A(n5659), .ZN(n12317) );
  INV_X1 U277 ( .A(n5676), .ZN(n12300) );
  INV_X1 U278 ( .A(n5693), .ZN(n12283) );
  INV_X1 U279 ( .A(n5710), .ZN(n12266) );
  INV_X1 U280 ( .A(n5727), .ZN(n12249) );
  INV_X1 U281 ( .A(n5745), .ZN(n12232) );
  INV_X1 U282 ( .A(n5763), .ZN(n12215) );
  INV_X1 U283 ( .A(n5780), .ZN(n12198) );
  INV_X1 U284 ( .A(n5797), .ZN(n12181) );
  INV_X1 U285 ( .A(n5814), .ZN(n12164) );
  INV_X1 U286 ( .A(n5831), .ZN(n12147) );
  INV_X1 U287 ( .A(n5848), .ZN(n12130) );
  INV_X1 U288 ( .A(n5865), .ZN(n12113) );
  INV_X1 U289 ( .A(n5882), .ZN(n12096) );
  INV_X1 U290 ( .A(n5899), .ZN(n12079) );
  INV_X1 U291 ( .A(n5916), .ZN(n12062) );
  INV_X1 U292 ( .A(n5933), .ZN(n12045) );
  INV_X1 U293 ( .A(n5950), .ZN(n12028) );
  INV_X1 U294 ( .A(n5967), .ZN(n12011) );
  INV_X1 U295 ( .A(n5984), .ZN(n11994) );
  INV_X1 U296 ( .A(n6001), .ZN(n11977) );
  INV_X1 U297 ( .A(n6018), .ZN(n11960) );
  INV_X1 U298 ( .A(n6036), .ZN(n11943) );
  INV_X1 U299 ( .A(n6053), .ZN(n11926) );
  INV_X1 U300 ( .A(n6070), .ZN(n11909) );
  INV_X1 U301 ( .A(n6087), .ZN(n11892) );
  INV_X1 U302 ( .A(n6104), .ZN(n11875) );
  INV_X1 U303 ( .A(n6121), .ZN(n11858) );
  INV_X1 U304 ( .A(n6138), .ZN(n11841) );
  INV_X1 U305 ( .A(n6155), .ZN(n11824) );
  INV_X1 U306 ( .A(n6172), .ZN(n11807) );
  INV_X1 U307 ( .A(n6189), .ZN(n11790) );
  INV_X1 U308 ( .A(n6206), .ZN(n11773) );
  INV_X1 U309 ( .A(n6223), .ZN(n11756) );
  INV_X1 U310 ( .A(n6240), .ZN(n11739) );
  INV_X1 U311 ( .A(n6257), .ZN(n11722) );
  INV_X1 U312 ( .A(n6274), .ZN(n11705) );
  INV_X1 U313 ( .A(n6291), .ZN(n11688) );
  INV_X1 U314 ( .A(n6309), .ZN(n11671) );
  INV_X1 U315 ( .A(n6326), .ZN(n11654) );
  INV_X1 U316 ( .A(n6343), .ZN(n11637) );
  INV_X1 U317 ( .A(n6360), .ZN(n11620) );
  INV_X1 U318 ( .A(n6377), .ZN(n11603) );
  INV_X1 U319 ( .A(n6394), .ZN(n11586) );
  INV_X1 U320 ( .A(n6411), .ZN(n11569) );
  INV_X1 U321 ( .A(n6428), .ZN(n11552) );
  INV_X1 U322 ( .A(n6445), .ZN(n11535) );
  INV_X1 U323 ( .A(n6462), .ZN(n11518) );
  INV_X1 U324 ( .A(n6479), .ZN(n11501) );
  INV_X1 U325 ( .A(n6496), .ZN(n11484) );
  INV_X1 U326 ( .A(n6513), .ZN(n11467) );
  INV_X1 U327 ( .A(n6530), .ZN(n11450) );
  INV_X1 U328 ( .A(n6547), .ZN(n11433) );
  INV_X1 U329 ( .A(n6564), .ZN(n11416) );
  INV_X1 U330 ( .A(n6582), .ZN(n11399) );
  INV_X1 U331 ( .A(n6599), .ZN(n11382) );
  INV_X1 U332 ( .A(n6616), .ZN(n11365) );
  INV_X1 U333 ( .A(n6633), .ZN(n11348) );
  INV_X1 U334 ( .A(n6650), .ZN(n11331) );
  INV_X1 U335 ( .A(n6667), .ZN(n11314) );
  INV_X1 U336 ( .A(n6684), .ZN(n11297) );
  INV_X1 U337 ( .A(n6701), .ZN(n11280) );
  INV_X1 U338 ( .A(n6718), .ZN(n11263) );
  INV_X1 U339 ( .A(n6735), .ZN(n11246) );
  INV_X1 U340 ( .A(n6752), .ZN(n11229) );
  INV_X1 U341 ( .A(n6769), .ZN(n11212) );
  INV_X1 U342 ( .A(n6786), .ZN(n11195) );
  INV_X1 U343 ( .A(n6803), .ZN(n11178) );
  INV_X1 U344 ( .A(n6820), .ZN(n11161) );
  INV_X1 U345 ( .A(n6838), .ZN(n11144) );
  INV_X1 U346 ( .A(n6856), .ZN(n11127) );
  INV_X1 U347 ( .A(n6873), .ZN(n11110) );
  INV_X1 U348 ( .A(n6890), .ZN(n11093) );
  INV_X1 U349 ( .A(n6907), .ZN(n11076) );
  INV_X1 U350 ( .A(n6924), .ZN(n11059) );
  INV_X1 U351 ( .A(n6941), .ZN(n11042) );
  INV_X1 U352 ( .A(n6958), .ZN(n11025) );
  INV_X1 U353 ( .A(n6975), .ZN(n11008) );
  INV_X1 U354 ( .A(n6992), .ZN(n10991) );
  INV_X1 U355 ( .A(n7009), .ZN(n10974) );
  INV_X1 U356 ( .A(n7026), .ZN(n10957) );
  INV_X1 U357 ( .A(n7043), .ZN(n10940) );
  INV_X1 U358 ( .A(n7060), .ZN(n10923) );
  INV_X1 U359 ( .A(n7077), .ZN(n10906) );
  INV_X1 U360 ( .A(n7094), .ZN(n10889) );
  INV_X1 U361 ( .A(n7111), .ZN(n10872) );
  INV_X1 U362 ( .A(n7129), .ZN(n10855) );
  INV_X1 U363 ( .A(n7146), .ZN(n10838) );
  INV_X1 U364 ( .A(n7163), .ZN(n10821) );
  INV_X1 U365 ( .A(n7180), .ZN(n10804) );
  INV_X1 U366 ( .A(n7197), .ZN(n10787) );
  INV_X1 U367 ( .A(n7214), .ZN(n10770) );
  INV_X1 U368 ( .A(n7231), .ZN(n10753) );
  INV_X1 U369 ( .A(n7248), .ZN(n10736) );
  INV_X1 U370 ( .A(n7265), .ZN(n10719) );
  INV_X1 U371 ( .A(n7282), .ZN(n10702) );
  INV_X1 U372 ( .A(n7299), .ZN(n10685) );
  INV_X1 U373 ( .A(n7316), .ZN(n10668) );
  INV_X1 U374 ( .A(n7333), .ZN(n10651) );
  INV_X1 U375 ( .A(n7350), .ZN(n10634) );
  INV_X1 U376 ( .A(n7367), .ZN(n10617) );
  INV_X1 U377 ( .A(n7384), .ZN(n10600) );
  INV_X1 U378 ( .A(n7402), .ZN(n10583) );
  INV_X1 U379 ( .A(n7419), .ZN(n10566) );
  INV_X1 U380 ( .A(n7436), .ZN(n10549) );
  INV_X1 U381 ( .A(n7453), .ZN(n10532) );
  INV_X1 U382 ( .A(n7470), .ZN(n10515) );
  INV_X1 U383 ( .A(n7487), .ZN(n10498) );
  INV_X1 U384 ( .A(n7504), .ZN(n10481) );
  INV_X1 U385 ( .A(n7521), .ZN(n10464) );
  INV_X1 U386 ( .A(n7538), .ZN(n10447) );
  INV_X1 U387 ( .A(n7555), .ZN(n10430) );
  INV_X1 U388 ( .A(n7572), .ZN(n10413) );
  INV_X1 U389 ( .A(n7589), .ZN(n10396) );
  INV_X1 U390 ( .A(n7606), .ZN(n10379) );
  INV_X1 U391 ( .A(n7623), .ZN(n10362) );
  INV_X1 U392 ( .A(n7640), .ZN(n10345) );
  INV_X1 U393 ( .A(n7657), .ZN(n10328) );
  INV_X1 U394 ( .A(n7675), .ZN(n10311) );
  INV_X1 U395 ( .A(n7692), .ZN(n10294) );
  INV_X1 U396 ( .A(n7709), .ZN(n10277) );
  INV_X1 U397 ( .A(n7726), .ZN(n10260) );
  INV_X1 U398 ( .A(n7743), .ZN(n10243) );
  INV_X1 U399 ( .A(n7760), .ZN(n10226) );
  INV_X1 U400 ( .A(n7777), .ZN(n10209) );
  INV_X1 U401 ( .A(n7794), .ZN(n10192) );
  INV_X1 U402 ( .A(n7811), .ZN(n10175) );
  INV_X1 U403 ( .A(n7828), .ZN(n10158) );
  INV_X1 U404 ( .A(n7845), .ZN(n10141) );
  INV_X1 U405 ( .A(n7862), .ZN(n10124) );
  INV_X1 U406 ( .A(n7879), .ZN(n10107) );
  INV_X1 U407 ( .A(n7896), .ZN(n10090) );
  INV_X1 U408 ( .A(n7913), .ZN(n10073) );
  INV_X1 U409 ( .A(n7931), .ZN(n10056) );
  INV_X1 U410 ( .A(n7949), .ZN(n10039) );
  INV_X1 U411 ( .A(n7966), .ZN(n10022) );
  INV_X1 U412 ( .A(n7983), .ZN(n10005) );
  INV_X1 U413 ( .A(n8000), .ZN(n9988) );
  INV_X1 U414 ( .A(n8017), .ZN(n9971) );
  INV_X1 U415 ( .A(n8034), .ZN(n9954) );
  INV_X1 U416 ( .A(n8051), .ZN(n9937) );
  INV_X1 U417 ( .A(n8068), .ZN(n9920) );
  INV_X1 U418 ( .A(n8085), .ZN(n9903) );
  INV_X1 U419 ( .A(n8102), .ZN(n9886) );
  INV_X1 U420 ( .A(n8119), .ZN(n9869) );
  INV_X1 U421 ( .A(n8136), .ZN(n9852) );
  INV_X1 U422 ( .A(n8153), .ZN(n9835) );
  INV_X1 U423 ( .A(n8170), .ZN(n9818) );
  INV_X1 U424 ( .A(n8187), .ZN(n9801) );
  INV_X1 U425 ( .A(n8204), .ZN(n9784) );
  INV_X1 U426 ( .A(n8222), .ZN(n9767) );
  INV_X1 U427 ( .A(n8239), .ZN(n9750) );
  INV_X1 U428 ( .A(n8256), .ZN(n9733) );
  INV_X1 U429 ( .A(n8273), .ZN(n9716) );
  INV_X1 U430 ( .A(n8290), .ZN(n9699) );
  INV_X1 U431 ( .A(n8307), .ZN(n9682) );
  INV_X1 U432 ( .A(n8324), .ZN(n9665) );
  INV_X1 U433 ( .A(n8341), .ZN(n9648) );
  INV_X1 U434 ( .A(n8358), .ZN(n9631) );
  INV_X1 U435 ( .A(n8375), .ZN(n9614) );
  INV_X1 U436 ( .A(n8392), .ZN(n9597) );
  INV_X1 U437 ( .A(n8409), .ZN(n9580) );
  INV_X1 U438 ( .A(n8426), .ZN(n9563) );
  INV_X1 U439 ( .A(n8443), .ZN(n9546) );
  INV_X1 U440 ( .A(n8460), .ZN(n9529) );
  INV_X1 U441 ( .A(n8477), .ZN(n9512) );
  INV_X1 U442 ( .A(n8497), .ZN(n9495) );
  INV_X1 U443 ( .A(n8515), .ZN(n9478) );
  INV_X1 U444 ( .A(n8533), .ZN(n9461) );
  INV_X1 U445 ( .A(n8551), .ZN(n9444) );
  INV_X1 U446 ( .A(n8569), .ZN(n9427) );
  INV_X1 U447 ( .A(n8586), .ZN(n9410) );
  INV_X1 U448 ( .A(n8603), .ZN(n9393) );
  INV_X1 U449 ( .A(n8620), .ZN(n9376) );
  INV_X1 U450 ( .A(n8638), .ZN(n9359) );
  INV_X1 U451 ( .A(n8655), .ZN(n9342) );
  INV_X1 U452 ( .A(n8672), .ZN(n9325) );
  INV_X1 U453 ( .A(n8689), .ZN(n9308) );
  INV_X1 U454 ( .A(n8707), .ZN(n9291) );
  INV_X1 U455 ( .A(n8724), .ZN(n9274) );
  INV_X1 U456 ( .A(n8741), .ZN(n9257) );
  INV_X1 U457 ( .A(n4377), .ZN(n13575) );
  INV_X1 U458 ( .A(n4395), .ZN(n13558) );
  INV_X1 U459 ( .A(n4413), .ZN(n13541) );
  INV_X1 U460 ( .A(n4431), .ZN(n13524) );
  INV_X1 U461 ( .A(n4449), .ZN(n13507) );
  INV_X1 U462 ( .A(n4467), .ZN(n13490) );
  INV_X1 U463 ( .A(n4485), .ZN(n13473) );
  INV_X1 U464 ( .A(n4503), .ZN(n13456) );
  INV_X1 U465 ( .A(n4521), .ZN(n13439) );
  INV_X1 U466 ( .A(n4539), .ZN(n13422) );
  INV_X1 U467 ( .A(n4557), .ZN(n13405) );
  INV_X1 U468 ( .A(n4575), .ZN(n13388) );
  INV_X1 U469 ( .A(n4593), .ZN(n13371) );
  INV_X1 U470 ( .A(n4611), .ZN(n13354) );
  INV_X1 U471 ( .A(n4629), .ZN(n13337) );
  NOR2_X1 U472 ( .A1(mem_access_addr[2]), .A2(mem_access_addr[3]), .ZN(n8495)
         );
  NOR2_X1 U473 ( .A1(n9236), .A2(mem_access_addr[3]), .ZN(n8513) );
  NOR2_X1 U474 ( .A1(mem_access_addr[4]), .A2(mem_access_addr[5]), .ZN(n8494)
         );
  NOR2_X1 U475 ( .A1(n9237), .A2(mem_access_addr[5]), .ZN(n8567) );
  BUF_X1 U476 ( .A(n8853), .Z(n8874) );
  BUF_X1 U477 ( .A(n8877), .Z(n8898) );
  BUF_X1 U478 ( .A(n8901), .Z(n8922) );
  BUF_X1 U479 ( .A(n8925), .Z(n8946) );
  BUF_X1 U480 ( .A(n8949), .Z(n8970) );
  BUF_X1 U481 ( .A(n8973), .Z(n8994) );
  BUF_X1 U482 ( .A(n8997), .Z(n9018) );
  BUF_X1 U483 ( .A(n8853), .Z(n8873) );
  BUF_X1 U484 ( .A(n8877), .Z(n8897) );
  BUF_X1 U485 ( .A(n8901), .Z(n8921) );
  BUF_X1 U486 ( .A(n8925), .Z(n8945) );
  BUF_X1 U487 ( .A(n8949), .Z(n8969) );
  BUF_X1 U488 ( .A(n8973), .Z(n8993) );
  BUF_X1 U489 ( .A(n8997), .Z(n9017) );
  BUF_X1 U490 ( .A(n8853), .Z(n8872) );
  BUF_X1 U491 ( .A(n8877), .Z(n8896) );
  BUF_X1 U492 ( .A(n8901), .Z(n8920) );
  BUF_X1 U493 ( .A(n8925), .Z(n8944) );
  BUF_X1 U494 ( .A(n8949), .Z(n8968) );
  BUF_X1 U495 ( .A(n8973), .Z(n8992) );
  BUF_X1 U496 ( .A(n8997), .Z(n9016) );
  BUF_X1 U497 ( .A(n8853), .Z(n8871) );
  BUF_X1 U498 ( .A(n8877), .Z(n8895) );
  BUF_X1 U499 ( .A(n8901), .Z(n8919) );
  BUF_X1 U500 ( .A(n8925), .Z(n8943) );
  BUF_X1 U501 ( .A(n8949), .Z(n8967) );
  BUF_X1 U502 ( .A(n8973), .Z(n8991) );
  BUF_X1 U503 ( .A(n8997), .Z(n9015) );
  BUF_X1 U504 ( .A(n8852), .Z(n8864) );
  BUF_X1 U505 ( .A(n8876), .Z(n8888) );
  BUF_X1 U506 ( .A(n8900), .Z(n8912) );
  BUF_X1 U507 ( .A(n8924), .Z(n8936) );
  BUF_X1 U508 ( .A(n8948), .Z(n8960) );
  BUF_X1 U509 ( .A(n8972), .Z(n8984) );
  BUF_X1 U510 ( .A(n8996), .Z(n9008) );
  BUF_X1 U511 ( .A(n8852), .Z(n8863) );
  BUF_X1 U512 ( .A(n8876), .Z(n8887) );
  BUF_X1 U513 ( .A(n8900), .Z(n8911) );
  BUF_X1 U514 ( .A(n8924), .Z(n8935) );
  BUF_X1 U515 ( .A(n8948), .Z(n8959) );
  BUF_X1 U516 ( .A(n8972), .Z(n8983) );
  BUF_X1 U517 ( .A(n8996), .Z(n9007) );
  BUF_X1 U518 ( .A(n8852), .Z(n8862) );
  BUF_X1 U519 ( .A(n8876), .Z(n8886) );
  BUF_X1 U520 ( .A(n8900), .Z(n8910) );
  BUF_X1 U521 ( .A(n8924), .Z(n8934) );
  BUF_X1 U522 ( .A(n8948), .Z(n8958) );
  BUF_X1 U523 ( .A(n8972), .Z(n8982) );
  BUF_X1 U524 ( .A(n8996), .Z(n9006) );
  BUF_X1 U525 ( .A(n8852), .Z(n8861) );
  BUF_X1 U526 ( .A(n8876), .Z(n8885) );
  BUF_X1 U527 ( .A(n8900), .Z(n8909) );
  BUF_X1 U528 ( .A(n8924), .Z(n8933) );
  BUF_X1 U529 ( .A(n8948), .Z(n8957) );
  BUF_X1 U530 ( .A(n8972), .Z(n8981) );
  BUF_X1 U531 ( .A(n8996), .Z(n9005) );
  NOR2_X1 U532 ( .A1(n9240), .A2(mem_access_addr[9]), .ZN(n5743) );
  NOR2_X1 U533 ( .A1(mem_access_addr[8]), .A2(mem_access_addr[9]), .ZN(n4646)
         );
  NOR2_X1 U534 ( .A1(n9238), .A2(mem_access_addr[7]), .ZN(n4647) );
  NOR2_X1 U535 ( .A1(n9239), .A2(mem_access_addr[7]), .ZN(n4921) );
  AND2_X1 U536 ( .A1(mem_access_addr[3]), .A2(mem_access_addr[2]), .ZN(n8549)
         );
  AND2_X1 U537 ( .A1(mem_access_addr[3]), .A2(n9236), .ZN(n8531) );
  AND2_X1 U538 ( .A1(mem_access_addr[5]), .A2(n9237), .ZN(n8636) );
  AND2_X1 U539 ( .A1(mem_access_addr[5]), .A2(mem_access_addr[4]), .ZN(n8705)
         );
  AND2_X1 U540 ( .A1(mem_access_addr[9]), .A2(n9240), .ZN(n6836) );
  AND2_X1 U541 ( .A1(mem_access_addr[9]), .A2(mem_access_addr[8]), .ZN(n7929)
         );
  AND2_X1 U542 ( .A1(mem_access_addr[7]), .A2(n9238), .ZN(n5469) );
  AND2_X1 U543 ( .A1(mem_access_addr[7]), .A2(n9239), .ZN(n5195) );
  BUF_X1 U544 ( .A(mem_access_addr[5]), .Z(n4109) );
  BUF_X1 U545 ( .A(mem_access_addr[5]), .Z(n4110) );
  INV_X1 U546 ( .A(mem_access_addr[2]), .ZN(n9236) );
  BUF_X1 U547 ( .A(mem_access_addr[3]), .Z(n4262) );
  BUF_X1 U548 ( .A(mem_access_addr[3]), .Z(n4261) );
  BUF_X1 U549 ( .A(mem_access_addr[3]), .Z(n4260) );
  NAND2_X1 U550 ( .A1(n4665), .A2(n4374), .ZN(n4649) );
  NAND2_X1 U551 ( .A1(n4665), .A2(n4393), .ZN(n4667) );
  NAND2_X1 U552 ( .A1(n4665), .A2(n4411), .ZN(n4684) );
  NAND2_X1 U553 ( .A1(n4665), .A2(n4429), .ZN(n4701) );
  NAND2_X1 U554 ( .A1(n4665), .A2(n4447), .ZN(n4718) );
  NAND2_X1 U555 ( .A1(n4665), .A2(n4465), .ZN(n4735) );
  NAND2_X1 U556 ( .A1(n4665), .A2(n4483), .ZN(n4752) );
  NAND2_X1 U557 ( .A1(n4665), .A2(n4501), .ZN(n4769) );
  NAND2_X1 U558 ( .A1(n4665), .A2(n4519), .ZN(n4786) );
  NAND2_X1 U559 ( .A1(n4665), .A2(n4537), .ZN(n4803) );
  NAND2_X1 U560 ( .A1(n4665), .A2(n4555), .ZN(n4820) );
  NAND2_X1 U561 ( .A1(n4665), .A2(n4573), .ZN(n4837) );
  NAND2_X1 U562 ( .A1(n4665), .A2(n4591), .ZN(n4854) );
  NAND2_X1 U563 ( .A1(n4665), .A2(n4609), .ZN(n4871) );
  NAND2_X1 U564 ( .A1(n4665), .A2(n4627), .ZN(n4888) );
  NAND2_X1 U565 ( .A1(n4665), .A2(n4645), .ZN(n4905) );
  NAND2_X1 U566 ( .A1(n4939), .A2(n4374), .ZN(n4923) );
  NAND2_X1 U567 ( .A1(n4939), .A2(n4393), .ZN(n4941) );
  NAND2_X1 U568 ( .A1(n4939), .A2(n4411), .ZN(n4958) );
  NAND2_X1 U569 ( .A1(n4939), .A2(n4429), .ZN(n4975) );
  NAND2_X1 U570 ( .A1(n4939), .A2(n4447), .ZN(n4992) );
  NAND2_X1 U571 ( .A1(n4939), .A2(n4465), .ZN(n5009) );
  NAND2_X1 U572 ( .A1(n4939), .A2(n4483), .ZN(n5026) );
  NAND2_X1 U573 ( .A1(n4939), .A2(n4501), .ZN(n5043) );
  NAND2_X1 U574 ( .A1(n4939), .A2(n4519), .ZN(n5060) );
  NAND2_X1 U575 ( .A1(n4939), .A2(n4537), .ZN(n5077) );
  NAND2_X1 U576 ( .A1(n4939), .A2(n4555), .ZN(n5094) );
  NAND2_X1 U577 ( .A1(n4939), .A2(n4573), .ZN(n5111) );
  NAND2_X1 U578 ( .A1(n4939), .A2(n4591), .ZN(n5128) );
  NAND2_X1 U579 ( .A1(n4939), .A2(n4609), .ZN(n5145) );
  NAND2_X1 U580 ( .A1(n4939), .A2(n4627), .ZN(n5162) );
  NAND2_X1 U581 ( .A1(n4939), .A2(n4645), .ZN(n5179) );
  NAND2_X1 U582 ( .A1(n5213), .A2(n4374), .ZN(n5197) );
  NAND2_X1 U583 ( .A1(n5213), .A2(n4393), .ZN(n5215) );
  NAND2_X1 U584 ( .A1(n5213), .A2(n4411), .ZN(n5232) );
  NAND2_X1 U585 ( .A1(n5213), .A2(n4429), .ZN(n5249) );
  NAND2_X1 U586 ( .A1(n5213), .A2(n4447), .ZN(n5266) );
  NAND2_X1 U587 ( .A1(n5213), .A2(n4465), .ZN(n5283) );
  NAND2_X1 U588 ( .A1(n5213), .A2(n4483), .ZN(n5300) );
  NAND2_X1 U589 ( .A1(n5213), .A2(n4501), .ZN(n5317) );
  NAND2_X1 U590 ( .A1(n5213), .A2(n4519), .ZN(n5334) );
  NAND2_X1 U591 ( .A1(n5213), .A2(n4537), .ZN(n5351) );
  NAND2_X1 U592 ( .A1(n5213), .A2(n4555), .ZN(n5368) );
  NAND2_X1 U593 ( .A1(n5213), .A2(n4573), .ZN(n5385) );
  NAND2_X1 U594 ( .A1(n5213), .A2(n4591), .ZN(n5402) );
  NAND2_X1 U595 ( .A1(n5213), .A2(n4609), .ZN(n5419) );
  NAND2_X1 U596 ( .A1(n5213), .A2(n4627), .ZN(n5436) );
  NAND2_X1 U597 ( .A1(n5213), .A2(n4645), .ZN(n5453) );
  NAND2_X1 U598 ( .A1(n5487), .A2(n4374), .ZN(n5471) );
  NAND2_X1 U599 ( .A1(n5487), .A2(n4393), .ZN(n5489) );
  NAND2_X1 U600 ( .A1(n5487), .A2(n4411), .ZN(n5506) );
  NAND2_X1 U601 ( .A1(n5487), .A2(n4429), .ZN(n5523) );
  NAND2_X1 U602 ( .A1(n5487), .A2(n4447), .ZN(n5540) );
  NAND2_X1 U603 ( .A1(n5487), .A2(n4465), .ZN(n5557) );
  NAND2_X1 U604 ( .A1(n5487), .A2(n4483), .ZN(n5574) );
  NAND2_X1 U605 ( .A1(n5487), .A2(n4501), .ZN(n5591) );
  NAND2_X1 U606 ( .A1(n5487), .A2(n4519), .ZN(n5608) );
  NAND2_X1 U607 ( .A1(n5487), .A2(n4537), .ZN(n5625) );
  NAND2_X1 U608 ( .A1(n5487), .A2(n4555), .ZN(n5642) );
  NAND2_X1 U609 ( .A1(n5487), .A2(n4573), .ZN(n5659) );
  NAND2_X1 U610 ( .A1(n5487), .A2(n4591), .ZN(n5676) );
  NAND2_X1 U611 ( .A1(n5487), .A2(n4609), .ZN(n5693) );
  NAND2_X1 U612 ( .A1(n5487), .A2(n4627), .ZN(n5710) );
  NAND2_X1 U613 ( .A1(n5487), .A2(n4645), .ZN(n5727) );
  NAND2_X1 U614 ( .A1(n6580), .A2(n4374), .ZN(n6564) );
  NAND2_X1 U615 ( .A1(n6580), .A2(n4393), .ZN(n6582) );
  NAND2_X1 U616 ( .A1(n6580), .A2(n4411), .ZN(n6599) );
  NAND2_X1 U617 ( .A1(n6580), .A2(n4429), .ZN(n6616) );
  NAND2_X1 U618 ( .A1(n6580), .A2(n4447), .ZN(n6633) );
  NAND2_X1 U619 ( .A1(n6580), .A2(n4465), .ZN(n6650) );
  NAND2_X1 U620 ( .A1(n6580), .A2(n4483), .ZN(n6667) );
  NAND2_X1 U621 ( .A1(n6580), .A2(n4501), .ZN(n6684) );
  NAND2_X1 U622 ( .A1(n6580), .A2(n4519), .ZN(n6701) );
  NAND2_X1 U623 ( .A1(n6580), .A2(n4537), .ZN(n6718) );
  NAND2_X1 U624 ( .A1(n6580), .A2(n4555), .ZN(n6735) );
  NAND2_X1 U625 ( .A1(n6580), .A2(n4573), .ZN(n6752) );
  NAND2_X1 U626 ( .A1(n6580), .A2(n4591), .ZN(n6769) );
  NAND2_X1 U627 ( .A1(n6580), .A2(n4609), .ZN(n6786) );
  NAND2_X1 U628 ( .A1(n6580), .A2(n4627), .ZN(n6803) );
  NAND2_X1 U629 ( .A1(n6580), .A2(n4645), .ZN(n6820) );
  NAND2_X1 U630 ( .A1(n7673), .A2(n4374), .ZN(n7657) );
  NAND2_X1 U631 ( .A1(n7673), .A2(n4393), .ZN(n7675) );
  NAND2_X1 U632 ( .A1(n7673), .A2(n4411), .ZN(n7692) );
  NAND2_X1 U633 ( .A1(n7673), .A2(n4429), .ZN(n7709) );
  NAND2_X1 U634 ( .A1(n7673), .A2(n4447), .ZN(n7726) );
  NAND2_X1 U635 ( .A1(n7673), .A2(n4465), .ZN(n7743) );
  NAND2_X1 U636 ( .A1(n7673), .A2(n4483), .ZN(n7760) );
  NAND2_X1 U637 ( .A1(n7673), .A2(n4501), .ZN(n7777) );
  NAND2_X1 U638 ( .A1(n7673), .A2(n4519), .ZN(n7794) );
  NAND2_X1 U639 ( .A1(n7673), .A2(n4537), .ZN(n7811) );
  NAND2_X1 U640 ( .A1(n7673), .A2(n4555), .ZN(n7828) );
  NAND2_X1 U641 ( .A1(n7673), .A2(n4573), .ZN(n7845) );
  NAND2_X1 U642 ( .A1(n7673), .A2(n4591), .ZN(n7862) );
  NAND2_X1 U643 ( .A1(n7673), .A2(n4609), .ZN(n7879) );
  NAND2_X1 U644 ( .A1(n7673), .A2(n4627), .ZN(n7896) );
  NAND2_X1 U645 ( .A1(n7673), .A2(n4645), .ZN(n7913) );
  NAND2_X1 U646 ( .A1(n5761), .A2(n4374), .ZN(n5745) );
  NAND2_X1 U647 ( .A1(n5761), .A2(n4393), .ZN(n5763) );
  NAND2_X1 U648 ( .A1(n5761), .A2(n4411), .ZN(n5780) );
  NAND2_X1 U649 ( .A1(n5761), .A2(n4429), .ZN(n5797) );
  NAND2_X1 U650 ( .A1(n5761), .A2(n4447), .ZN(n5814) );
  NAND2_X1 U651 ( .A1(n5761), .A2(n4465), .ZN(n5831) );
  NAND2_X1 U652 ( .A1(n5761), .A2(n4483), .ZN(n5848) );
  NAND2_X1 U653 ( .A1(n5761), .A2(n4501), .ZN(n5865) );
  NAND2_X1 U654 ( .A1(n5761), .A2(n4519), .ZN(n5882) );
  NAND2_X1 U655 ( .A1(n5761), .A2(n4537), .ZN(n5899) );
  NAND2_X1 U656 ( .A1(n5761), .A2(n4555), .ZN(n5916) );
  NAND2_X1 U657 ( .A1(n5761), .A2(n4573), .ZN(n5933) );
  NAND2_X1 U658 ( .A1(n5761), .A2(n4591), .ZN(n5950) );
  NAND2_X1 U659 ( .A1(n5761), .A2(n4609), .ZN(n5967) );
  NAND2_X1 U660 ( .A1(n5761), .A2(n4627), .ZN(n5984) );
  NAND2_X1 U661 ( .A1(n5761), .A2(n4645), .ZN(n6001) );
  NAND2_X1 U662 ( .A1(n6034), .A2(n4374), .ZN(n6018) );
  NAND2_X1 U663 ( .A1(n6034), .A2(n4393), .ZN(n6036) );
  NAND2_X1 U664 ( .A1(n6034), .A2(n4411), .ZN(n6053) );
  NAND2_X1 U665 ( .A1(n6034), .A2(n4429), .ZN(n6070) );
  NAND2_X1 U666 ( .A1(n6034), .A2(n4447), .ZN(n6087) );
  NAND2_X1 U667 ( .A1(n6034), .A2(n4465), .ZN(n6104) );
  NAND2_X1 U668 ( .A1(n6034), .A2(n4483), .ZN(n6121) );
  NAND2_X1 U669 ( .A1(n6034), .A2(n4501), .ZN(n6138) );
  NAND2_X1 U670 ( .A1(n6034), .A2(n4519), .ZN(n6155) );
  NAND2_X1 U671 ( .A1(n6034), .A2(n4537), .ZN(n6172) );
  NAND2_X1 U672 ( .A1(n6034), .A2(n4555), .ZN(n6189) );
  NAND2_X1 U673 ( .A1(n6034), .A2(n4573), .ZN(n6206) );
  NAND2_X1 U674 ( .A1(n6034), .A2(n4591), .ZN(n6223) );
  NAND2_X1 U675 ( .A1(n6034), .A2(n4609), .ZN(n6240) );
  NAND2_X1 U676 ( .A1(n6034), .A2(n4627), .ZN(n6257) );
  NAND2_X1 U677 ( .A1(n6034), .A2(n4645), .ZN(n6274) );
  NAND2_X1 U678 ( .A1(n6307), .A2(n4374), .ZN(n6291) );
  NAND2_X1 U679 ( .A1(n6307), .A2(n4393), .ZN(n6309) );
  NAND2_X1 U680 ( .A1(n6307), .A2(n4411), .ZN(n6326) );
  NAND2_X1 U681 ( .A1(n6307), .A2(n4429), .ZN(n6343) );
  NAND2_X1 U682 ( .A1(n6307), .A2(n4447), .ZN(n6360) );
  NAND2_X1 U683 ( .A1(n6307), .A2(n4465), .ZN(n6377) );
  NAND2_X1 U684 ( .A1(n6307), .A2(n4483), .ZN(n6394) );
  NAND2_X1 U685 ( .A1(n6307), .A2(n4501), .ZN(n6411) );
  NAND2_X1 U686 ( .A1(n6307), .A2(n4519), .ZN(n6428) );
  NAND2_X1 U687 ( .A1(n6307), .A2(n4537), .ZN(n6445) );
  NAND2_X1 U688 ( .A1(n6307), .A2(n4555), .ZN(n6462) );
  NAND2_X1 U689 ( .A1(n6307), .A2(n4573), .ZN(n6479) );
  NAND2_X1 U690 ( .A1(n6307), .A2(n4591), .ZN(n6496) );
  NAND2_X1 U691 ( .A1(n6307), .A2(n4609), .ZN(n6513) );
  NAND2_X1 U692 ( .A1(n6307), .A2(n4627), .ZN(n6530) );
  NAND2_X1 U693 ( .A1(n6307), .A2(n4645), .ZN(n6547) );
  NAND2_X1 U694 ( .A1(n6854), .A2(n4374), .ZN(n6838) );
  NAND2_X1 U695 ( .A1(n6854), .A2(n4393), .ZN(n6856) );
  NAND2_X1 U696 ( .A1(n6854), .A2(n4411), .ZN(n6873) );
  NAND2_X1 U697 ( .A1(n6854), .A2(n4429), .ZN(n6890) );
  NAND2_X1 U698 ( .A1(n6854), .A2(n4447), .ZN(n6907) );
  NAND2_X1 U699 ( .A1(n6854), .A2(n4465), .ZN(n6924) );
  NAND2_X1 U700 ( .A1(n6854), .A2(n4483), .ZN(n6941) );
  NAND2_X1 U701 ( .A1(n6854), .A2(n4501), .ZN(n6958) );
  NAND2_X1 U702 ( .A1(n6854), .A2(n4519), .ZN(n6975) );
  NAND2_X1 U703 ( .A1(n6854), .A2(n4537), .ZN(n6992) );
  NAND2_X1 U704 ( .A1(n6854), .A2(n4555), .ZN(n7009) );
  NAND2_X1 U705 ( .A1(n6854), .A2(n4573), .ZN(n7026) );
  NAND2_X1 U706 ( .A1(n6854), .A2(n4591), .ZN(n7043) );
  NAND2_X1 U707 ( .A1(n6854), .A2(n4609), .ZN(n7060) );
  NAND2_X1 U708 ( .A1(n6854), .A2(n4627), .ZN(n7077) );
  NAND2_X1 U709 ( .A1(n6854), .A2(n4645), .ZN(n7094) );
  NAND2_X1 U710 ( .A1(n7127), .A2(n4374), .ZN(n7111) );
  NAND2_X1 U711 ( .A1(n7127), .A2(n4393), .ZN(n7129) );
  NAND2_X1 U712 ( .A1(n7127), .A2(n4411), .ZN(n7146) );
  NAND2_X1 U713 ( .A1(n7127), .A2(n4429), .ZN(n7163) );
  NAND2_X1 U714 ( .A1(n7127), .A2(n4447), .ZN(n7180) );
  NAND2_X1 U715 ( .A1(n7127), .A2(n4465), .ZN(n7197) );
  NAND2_X1 U716 ( .A1(n7127), .A2(n4483), .ZN(n7214) );
  NAND2_X1 U717 ( .A1(n7127), .A2(n4501), .ZN(n7231) );
  NAND2_X1 U718 ( .A1(n7127), .A2(n4519), .ZN(n7248) );
  NAND2_X1 U719 ( .A1(n7127), .A2(n4537), .ZN(n7265) );
  NAND2_X1 U720 ( .A1(n7127), .A2(n4555), .ZN(n7282) );
  NAND2_X1 U721 ( .A1(n7127), .A2(n4573), .ZN(n7299) );
  NAND2_X1 U722 ( .A1(n7127), .A2(n4591), .ZN(n7316) );
  NAND2_X1 U723 ( .A1(n7127), .A2(n4609), .ZN(n7333) );
  NAND2_X1 U724 ( .A1(n7127), .A2(n4627), .ZN(n7350) );
  NAND2_X1 U725 ( .A1(n7127), .A2(n4645), .ZN(n7367) );
  NAND2_X1 U726 ( .A1(n7400), .A2(n4374), .ZN(n7384) );
  NAND2_X1 U727 ( .A1(n7400), .A2(n4393), .ZN(n7402) );
  NAND2_X1 U728 ( .A1(n7400), .A2(n4411), .ZN(n7419) );
  NAND2_X1 U729 ( .A1(n7400), .A2(n4429), .ZN(n7436) );
  NAND2_X1 U730 ( .A1(n7400), .A2(n4447), .ZN(n7453) );
  NAND2_X1 U731 ( .A1(n7400), .A2(n4465), .ZN(n7470) );
  NAND2_X1 U732 ( .A1(n7400), .A2(n4483), .ZN(n7487) );
  NAND2_X1 U733 ( .A1(n7400), .A2(n4501), .ZN(n7504) );
  NAND2_X1 U734 ( .A1(n7400), .A2(n4519), .ZN(n7521) );
  NAND2_X1 U735 ( .A1(n7400), .A2(n4537), .ZN(n7538) );
  NAND2_X1 U736 ( .A1(n7400), .A2(n4555), .ZN(n7555) );
  NAND2_X1 U737 ( .A1(n7400), .A2(n4573), .ZN(n7572) );
  NAND2_X1 U738 ( .A1(n7400), .A2(n4591), .ZN(n7589) );
  NAND2_X1 U739 ( .A1(n7400), .A2(n4609), .ZN(n7606) );
  NAND2_X1 U740 ( .A1(n7400), .A2(n4627), .ZN(n7623) );
  NAND2_X1 U741 ( .A1(n7400), .A2(n4645), .ZN(n7640) );
  NAND2_X1 U742 ( .A1(n7947), .A2(n4374), .ZN(n7931) );
  NAND2_X1 U743 ( .A1(n7947), .A2(n4393), .ZN(n7949) );
  NAND2_X1 U744 ( .A1(n7947), .A2(n4411), .ZN(n7966) );
  NAND2_X1 U745 ( .A1(n7947), .A2(n4429), .ZN(n7983) );
  NAND2_X1 U746 ( .A1(n7947), .A2(n4447), .ZN(n8000) );
  NAND2_X1 U747 ( .A1(n7947), .A2(n4465), .ZN(n8017) );
  NAND2_X1 U748 ( .A1(n7947), .A2(n4483), .ZN(n8034) );
  NAND2_X1 U749 ( .A1(n7947), .A2(n4501), .ZN(n8051) );
  NAND2_X1 U750 ( .A1(n7947), .A2(n4519), .ZN(n8068) );
  NAND2_X1 U751 ( .A1(n7947), .A2(n4537), .ZN(n8085) );
  NAND2_X1 U752 ( .A1(n7947), .A2(n4555), .ZN(n8102) );
  NAND2_X1 U753 ( .A1(n7947), .A2(n4573), .ZN(n8119) );
  NAND2_X1 U754 ( .A1(n7947), .A2(n4591), .ZN(n8136) );
  NAND2_X1 U755 ( .A1(n7947), .A2(n4609), .ZN(n8153) );
  NAND2_X1 U756 ( .A1(n7947), .A2(n4627), .ZN(n8170) );
  NAND2_X1 U757 ( .A1(n7947), .A2(n4645), .ZN(n8187) );
  NAND2_X1 U758 ( .A1(n8220), .A2(n4374), .ZN(n8204) );
  NAND2_X1 U759 ( .A1(n8220), .A2(n4393), .ZN(n8222) );
  NAND2_X1 U760 ( .A1(n8220), .A2(n4411), .ZN(n8239) );
  NAND2_X1 U761 ( .A1(n8220), .A2(n4429), .ZN(n8256) );
  NAND2_X1 U762 ( .A1(n8220), .A2(n4447), .ZN(n8273) );
  NAND2_X1 U763 ( .A1(n8220), .A2(n4465), .ZN(n8290) );
  NAND2_X1 U764 ( .A1(n8220), .A2(n4483), .ZN(n8307) );
  NAND2_X1 U765 ( .A1(n8220), .A2(n4501), .ZN(n8324) );
  NAND2_X1 U766 ( .A1(n8220), .A2(n4519), .ZN(n8341) );
  NAND2_X1 U767 ( .A1(n8220), .A2(n4537), .ZN(n8358) );
  NAND2_X1 U768 ( .A1(n8220), .A2(n4555), .ZN(n8375) );
  NAND2_X1 U769 ( .A1(n8220), .A2(n4573), .ZN(n8392) );
  NAND2_X1 U770 ( .A1(n8220), .A2(n4591), .ZN(n8409) );
  NAND2_X1 U771 ( .A1(n8220), .A2(n4609), .ZN(n8426) );
  NAND2_X1 U772 ( .A1(n8220), .A2(n4627), .ZN(n8443) );
  NAND2_X1 U773 ( .A1(n8220), .A2(n4645), .ZN(n8460) );
  NAND2_X1 U774 ( .A1(n8493), .A2(n4374), .ZN(n8477) );
  NAND2_X1 U775 ( .A1(n8493), .A2(n4393), .ZN(n8497) );
  NAND2_X1 U776 ( .A1(n8493), .A2(n4411), .ZN(n8515) );
  NAND2_X1 U777 ( .A1(n8493), .A2(n4429), .ZN(n8533) );
  NAND2_X1 U778 ( .A1(n8493), .A2(n4447), .ZN(n8551) );
  NAND2_X1 U779 ( .A1(n8493), .A2(n4465), .ZN(n8569) );
  NAND2_X1 U780 ( .A1(n8493), .A2(n4483), .ZN(n8586) );
  NAND2_X1 U781 ( .A1(n8493), .A2(n4501), .ZN(n8603) );
  NAND2_X1 U782 ( .A1(n8493), .A2(n4519), .ZN(n8620) );
  NAND2_X1 U783 ( .A1(n8493), .A2(n4537), .ZN(n8638) );
  NAND2_X1 U784 ( .A1(n8493), .A2(n4555), .ZN(n8655) );
  NAND2_X1 U785 ( .A1(n8493), .A2(n4573), .ZN(n8672) );
  NAND2_X1 U786 ( .A1(n8493), .A2(n4591), .ZN(n8689) );
  NAND2_X1 U787 ( .A1(n8493), .A2(n4609), .ZN(n8707) );
  NAND2_X1 U788 ( .A1(n8493), .A2(n4627), .ZN(n8724) );
  NAND2_X1 U789 ( .A1(n8493), .A2(n4645), .ZN(n8741) );
  NAND2_X1 U790 ( .A1(n4374), .A2(n4375), .ZN(n4358) );
  NAND2_X1 U791 ( .A1(n4393), .A2(n4375), .ZN(n4377) );
  NAND2_X1 U792 ( .A1(n4411), .A2(n4375), .ZN(n4395) );
  NAND2_X1 U793 ( .A1(n4429), .A2(n4375), .ZN(n4413) );
  NAND2_X1 U794 ( .A1(n4447), .A2(n4375), .ZN(n4431) );
  NAND2_X1 U795 ( .A1(n4465), .A2(n4375), .ZN(n4449) );
  NAND2_X1 U796 ( .A1(n4483), .A2(n4375), .ZN(n4467) );
  NAND2_X1 U797 ( .A1(n4501), .A2(n4375), .ZN(n4485) );
  NAND2_X1 U798 ( .A1(n4519), .A2(n4375), .ZN(n4503) );
  NAND2_X1 U799 ( .A1(n4537), .A2(n4375), .ZN(n4521) );
  NAND2_X1 U800 ( .A1(n4555), .A2(n4375), .ZN(n4539) );
  NAND2_X1 U801 ( .A1(n4573), .A2(n4375), .ZN(n4557) );
  NAND2_X1 U802 ( .A1(n4591), .A2(n4375), .ZN(n4575) );
  NAND2_X1 U803 ( .A1(n4609), .A2(n4375), .ZN(n4593) );
  NAND2_X1 U804 ( .A1(n4627), .A2(n4375), .ZN(n4611) );
  NAND2_X1 U805 ( .A1(n4645), .A2(n4375), .ZN(n4629) );
  AND2_X1 U806 ( .A1(N286), .A2(mem_read), .ZN(mem_read_data[15]) );
  BUF_X1 U807 ( .A(n9021), .Z(n9042) );
  BUF_X1 U808 ( .A(n9045), .Z(n9066) );
  BUF_X1 U809 ( .A(n9069), .Z(n9090) );
  BUF_X1 U810 ( .A(n9093), .Z(n9114) );
  BUF_X1 U811 ( .A(n9117), .Z(n9138) );
  BUF_X1 U812 ( .A(n9141), .Z(n9162) );
  BUF_X1 U813 ( .A(n9165), .Z(n9186) );
  BUF_X1 U814 ( .A(n9189), .Z(n9210) );
  BUF_X1 U815 ( .A(n9213), .Z(n9234) );
  BUF_X1 U816 ( .A(n9021), .Z(n9041) );
  BUF_X1 U817 ( .A(n9045), .Z(n9065) );
  BUF_X1 U818 ( .A(n9069), .Z(n9089) );
  BUF_X1 U819 ( .A(n9093), .Z(n9113) );
  BUF_X1 U820 ( .A(n9117), .Z(n9137) );
  BUF_X1 U821 ( .A(n9141), .Z(n9161) );
  BUF_X1 U822 ( .A(n9165), .Z(n9185) );
  BUF_X1 U823 ( .A(n9189), .Z(n9209) );
  BUF_X1 U824 ( .A(n9213), .Z(n9233) );
  BUF_X1 U825 ( .A(n9021), .Z(n9040) );
  BUF_X1 U826 ( .A(n9045), .Z(n9064) );
  BUF_X1 U827 ( .A(n9069), .Z(n9088) );
  BUF_X1 U828 ( .A(n9093), .Z(n9112) );
  BUF_X1 U829 ( .A(n9117), .Z(n9136) );
  BUF_X1 U830 ( .A(n9141), .Z(n9160) );
  BUF_X1 U831 ( .A(n9165), .Z(n9184) );
  BUF_X1 U832 ( .A(n9189), .Z(n9208) );
  BUF_X1 U833 ( .A(n9213), .Z(n9232) );
  BUF_X1 U834 ( .A(n9021), .Z(n9039) );
  BUF_X1 U835 ( .A(n9045), .Z(n9063) );
  BUF_X1 U836 ( .A(n9069), .Z(n9087) );
  BUF_X1 U837 ( .A(n9093), .Z(n9111) );
  BUF_X1 U838 ( .A(n9117), .Z(n9135) );
  BUF_X1 U839 ( .A(n9141), .Z(n9159) );
  BUF_X1 U840 ( .A(n9165), .Z(n9183) );
  BUF_X1 U841 ( .A(n9189), .Z(n9207) );
  BUF_X1 U842 ( .A(n9213), .Z(n9231) );
  BUF_X1 U843 ( .A(n9020), .Z(n9032) );
  BUF_X1 U844 ( .A(n9044), .Z(n9056) );
  BUF_X1 U845 ( .A(n9068), .Z(n9080) );
  BUF_X1 U846 ( .A(n9092), .Z(n9104) );
  BUF_X1 U847 ( .A(n9116), .Z(n9128) );
  BUF_X1 U848 ( .A(n9140), .Z(n9152) );
  BUF_X1 U849 ( .A(n9164), .Z(n9176) );
  BUF_X1 U850 ( .A(n9188), .Z(n9200) );
  BUF_X1 U851 ( .A(n9212), .Z(n9224) );
  BUF_X1 U852 ( .A(n9020), .Z(n9031) );
  BUF_X1 U853 ( .A(n9044), .Z(n9055) );
  BUF_X1 U854 ( .A(n9068), .Z(n9079) );
  BUF_X1 U855 ( .A(n9092), .Z(n9103) );
  BUF_X1 U856 ( .A(n9116), .Z(n9127) );
  BUF_X1 U857 ( .A(n9140), .Z(n9151) );
  BUF_X1 U858 ( .A(n9164), .Z(n9175) );
  BUF_X1 U859 ( .A(n9188), .Z(n9199) );
  BUF_X1 U860 ( .A(n9212), .Z(n9223) );
  BUF_X1 U861 ( .A(n9020), .Z(n9030) );
  BUF_X1 U862 ( .A(n9044), .Z(n9054) );
  BUF_X1 U863 ( .A(n9068), .Z(n9078) );
  BUF_X1 U864 ( .A(n9092), .Z(n9102) );
  BUF_X1 U865 ( .A(n9116), .Z(n9126) );
  BUF_X1 U866 ( .A(n9140), .Z(n9150) );
  BUF_X1 U867 ( .A(n9164), .Z(n9174) );
  BUF_X1 U868 ( .A(n9188), .Z(n9198) );
  BUF_X1 U869 ( .A(n9212), .Z(n9222) );
  BUF_X1 U870 ( .A(n9020), .Z(n9029) );
  BUF_X1 U871 ( .A(n9044), .Z(n9053) );
  BUF_X1 U872 ( .A(n9068), .Z(n9077) );
  BUF_X1 U873 ( .A(n9092), .Z(n9101) );
  BUF_X1 U874 ( .A(n9116), .Z(n9125) );
  BUF_X1 U875 ( .A(n9140), .Z(n9149) );
  BUF_X1 U876 ( .A(n9164), .Z(n9173) );
  BUF_X1 U877 ( .A(n9188), .Z(n9197) );
  BUF_X1 U878 ( .A(n9212), .Z(n9221) );
  BUF_X1 U879 ( .A(mem_write_data[0]), .Z(n8853) );
  BUF_X1 U880 ( .A(mem_write_data[1]), .Z(n8877) );
  BUF_X1 U881 ( .A(mem_write_data[2]), .Z(n8901) );
  BUF_X1 U882 ( .A(mem_write_data[3]), .Z(n8925) );
  BUF_X1 U883 ( .A(mem_write_data[4]), .Z(n8949) );
  BUF_X1 U884 ( .A(mem_write_data[5]), .Z(n8973) );
  BUF_X1 U885 ( .A(mem_write_data[6]), .Z(n8997) );
  BUF_X1 U886 ( .A(mem_write_data[0]), .Z(n8852) );
  BUF_X1 U887 ( .A(mem_write_data[1]), .Z(n8876) );
  BUF_X1 U888 ( .A(mem_write_data[2]), .Z(n8900) );
  BUF_X1 U889 ( .A(mem_write_data[3]), .Z(n8924) );
  BUF_X1 U890 ( .A(mem_write_data[4]), .Z(n8948) );
  BUF_X1 U891 ( .A(mem_write_data[5]), .Z(n8972) );
  BUF_X1 U892 ( .A(mem_write_data[6]), .Z(n8996) );
  AND2_X1 U893 ( .A1(mem_read), .A2(N292), .ZN(mem_read_data[9]) );
  AND2_X1 U894 ( .A1(N301), .A2(mem_read), .ZN(mem_read_data[0]) );
  AND2_X1 U895 ( .A1(N299), .A2(mem_read), .ZN(mem_read_data[2]) );
  AND2_X1 U896 ( .A1(N298), .A2(mem_read), .ZN(mem_read_data[3]) );
  AND2_X1 U897 ( .A1(N297), .A2(mem_read), .ZN(mem_read_data[4]) );
  AND2_X1 U898 ( .A1(N296), .A2(mem_read), .ZN(mem_read_data[5]) );
  AND2_X1 U899 ( .A1(N295), .A2(mem_read), .ZN(mem_read_data[6]) );
  AND2_X1 U900 ( .A1(N294), .A2(mem_read), .ZN(mem_read_data[7]) );
  AND2_X1 U901 ( .A1(N293), .A2(mem_read), .ZN(mem_read_data[8]) );
  AND2_X1 U902 ( .A1(N291), .A2(mem_read), .ZN(mem_read_data[10]) );
  AND2_X1 U903 ( .A1(N290), .A2(mem_read), .ZN(mem_read_data[11]) );
  AND2_X1 U904 ( .A1(N289), .A2(mem_read), .ZN(mem_read_data[12]) );
  AND2_X1 U905 ( .A1(N288), .A2(mem_read), .ZN(mem_read_data[13]) );
  AND2_X1 U906 ( .A1(N287), .A2(mem_read), .ZN(mem_read_data[14]) );
  AND3_X1 U907 ( .A1(n4646), .A2(n4647), .A3(mem_write_en), .ZN(n4375) );
  AND3_X1 U908 ( .A1(mem_write_en), .A2(n4646), .A3(n4921), .ZN(n4665) );
  AND3_X1 U909 ( .A1(mem_write_en), .A2(n4646), .A3(n5195), .ZN(n4939) );
  AND3_X1 U910 ( .A1(mem_write_en), .A2(n4646), .A3(n5469), .ZN(n5213) );
  AND3_X1 U911 ( .A1(mem_write_en), .A2(n4647), .A3(n5743), .ZN(n5487) );
  AND3_X1 U912 ( .A1(mem_write_en), .A2(n4647), .A3(n6836), .ZN(n6580) );
  AND3_X1 U913 ( .A1(mem_write_en), .A2(n4647), .A3(n7929), .ZN(n7673) );
  AND3_X1 U914 ( .A1(n4921), .A2(mem_write_en), .A3(n5743), .ZN(n5761) );
  AND3_X1 U915 ( .A1(n5195), .A2(mem_write_en), .A3(n5743), .ZN(n6034) );
  AND3_X1 U916 ( .A1(n5469), .A2(mem_write_en), .A3(n5743), .ZN(n6307) );
  AND3_X1 U917 ( .A1(n4921), .A2(mem_write_en), .A3(n6836), .ZN(n6854) );
  AND3_X1 U918 ( .A1(n5195), .A2(mem_write_en), .A3(n6836), .ZN(n7127) );
  AND3_X1 U919 ( .A1(n5469), .A2(mem_write_en), .A3(n6836), .ZN(n7400) );
  AND3_X1 U920 ( .A1(n4921), .A2(mem_write_en), .A3(n7929), .ZN(n7947) );
  AND3_X1 U921 ( .A1(n5195), .A2(mem_write_en), .A3(n7929), .ZN(n8220) );
  AND3_X1 U922 ( .A1(n5469), .A2(mem_write_en), .A3(n7929), .ZN(n8493) );
  BUF_X1 U923 ( .A(mem_write_data[7]), .Z(n9021) );
  BUF_X1 U924 ( .A(mem_write_data[8]), .Z(n9045) );
  BUF_X1 U925 ( .A(mem_write_data[9]), .Z(n9069) );
  BUF_X1 U926 ( .A(mem_write_data[10]), .Z(n9093) );
  BUF_X1 U927 ( .A(mem_write_data[11]), .Z(n9117) );
  BUF_X1 U928 ( .A(mem_write_data[12]), .Z(n9141) );
  BUF_X1 U929 ( .A(mem_write_data[13]), .Z(n9165) );
  BUF_X1 U930 ( .A(mem_write_data[14]), .Z(n9189) );
  BUF_X1 U931 ( .A(mem_write_data[15]), .Z(n9213) );
  BUF_X1 U932 ( .A(mem_write_data[7]), .Z(n9020) );
  BUF_X1 U933 ( .A(mem_write_data[8]), .Z(n9044) );
  BUF_X1 U934 ( .A(mem_write_data[9]), .Z(n9068) );
  BUF_X1 U935 ( .A(mem_write_data[10]), .Z(n9092) );
  BUF_X1 U936 ( .A(mem_write_data[11]), .Z(n9116) );
  BUF_X1 U937 ( .A(mem_write_data[12]), .Z(n9140) );
  BUF_X1 U938 ( .A(mem_write_data[13]), .Z(n9164) );
  BUF_X1 U939 ( .A(mem_write_data[14]), .Z(n9188) );
  BUF_X1 U940 ( .A(mem_write_data[15]), .Z(n9212) );
  INV_X1 U941 ( .A(n4357), .ZN(n13576) );
  AOI22_X1 U942 ( .A1(ram[0]), .A2(n4358), .B1(n8875), .B2(n13592), .ZN(n4357)
         );
  INV_X1 U943 ( .A(n4359), .ZN(n13577) );
  AOI22_X1 U944 ( .A1(ram[1]), .A2(n4358), .B1(n8899), .B2(n13592), .ZN(n4359)
         );
  INV_X1 U945 ( .A(n4360), .ZN(n13578) );
  AOI22_X1 U946 ( .A1(ram[2]), .A2(n4358), .B1(n8923), .B2(n13592), .ZN(n4360)
         );
  INV_X1 U947 ( .A(n4361), .ZN(n13579) );
  AOI22_X1 U948 ( .A1(ram[3]), .A2(n4358), .B1(n8947), .B2(n13592), .ZN(n4361)
         );
  INV_X1 U949 ( .A(n4362), .ZN(n13580) );
  AOI22_X1 U950 ( .A1(ram[4]), .A2(n4358), .B1(n8971), .B2(n13592), .ZN(n4362)
         );
  INV_X1 U951 ( .A(n4363), .ZN(n13581) );
  AOI22_X1 U952 ( .A1(ram[5]), .A2(n4358), .B1(n8995), .B2(n13592), .ZN(n4363)
         );
  INV_X1 U953 ( .A(n4364), .ZN(n13582) );
  AOI22_X1 U954 ( .A1(ram[6]), .A2(n4358), .B1(n9019), .B2(n13592), .ZN(n4364)
         );
  INV_X1 U955 ( .A(n4365), .ZN(n13583) );
  AOI22_X1 U956 ( .A1(ram[7]), .A2(n4358), .B1(n9043), .B2(n13592), .ZN(n4365)
         );
  INV_X1 U957 ( .A(n4366), .ZN(n13584) );
  AOI22_X1 U958 ( .A1(ram[8]), .A2(n4358), .B1(n9067), .B2(n13592), .ZN(n4366)
         );
  INV_X1 U959 ( .A(n4367), .ZN(n13585) );
  AOI22_X1 U960 ( .A1(ram[9]), .A2(n4358), .B1(n9091), .B2(n13592), .ZN(n4367)
         );
  INV_X1 U961 ( .A(n4368), .ZN(n13586) );
  AOI22_X1 U962 ( .A1(ram[10]), .A2(n4358), .B1(n9115), .B2(n13592), .ZN(n4368) );
  INV_X1 U963 ( .A(n4369), .ZN(n13587) );
  AOI22_X1 U964 ( .A1(ram[11]), .A2(n4358), .B1(n9139), .B2(n13592), .ZN(n4369) );
  INV_X1 U965 ( .A(n4370), .ZN(n13588) );
  AOI22_X1 U966 ( .A1(ram[12]), .A2(n4358), .B1(n9163), .B2(n13592), .ZN(n4370) );
  INV_X1 U967 ( .A(n4371), .ZN(n13589) );
  AOI22_X1 U968 ( .A1(ram[13]), .A2(n4358), .B1(n9187), .B2(n13592), .ZN(n4371) );
  INV_X1 U969 ( .A(n4372), .ZN(n13590) );
  AOI22_X1 U970 ( .A1(ram[14]), .A2(n4358), .B1(n9211), .B2(n13592), .ZN(n4372) );
  INV_X1 U971 ( .A(n4373), .ZN(n13591) );
  AOI22_X1 U972 ( .A1(ram[15]), .A2(n4358), .B1(n9235), .B2(n13592), .ZN(n4373) );
  INV_X1 U973 ( .A(n4394), .ZN(n13542) );
  AOI22_X1 U974 ( .A1(ram[32]), .A2(n4395), .B1(n13558), .B2(n8875), .ZN(n4394) );
  INV_X1 U975 ( .A(n4396), .ZN(n13543) );
  AOI22_X1 U976 ( .A1(ram[33]), .A2(n4395), .B1(n13558), .B2(n8899), .ZN(n4396) );
  INV_X1 U977 ( .A(n4397), .ZN(n13544) );
  AOI22_X1 U978 ( .A1(ram[34]), .A2(n4395), .B1(n13558), .B2(n8923), .ZN(n4397) );
  INV_X1 U979 ( .A(n4398), .ZN(n13545) );
  AOI22_X1 U980 ( .A1(ram[35]), .A2(n4395), .B1(n13558), .B2(n8947), .ZN(n4398) );
  INV_X1 U981 ( .A(n4399), .ZN(n13546) );
  AOI22_X1 U982 ( .A1(ram[36]), .A2(n4395), .B1(n13558), .B2(n8971), .ZN(n4399) );
  INV_X1 U983 ( .A(n4400), .ZN(n13547) );
  AOI22_X1 U984 ( .A1(ram[37]), .A2(n4395), .B1(n13558), .B2(n8995), .ZN(n4400) );
  INV_X1 U985 ( .A(n4401), .ZN(n13548) );
  AOI22_X1 U986 ( .A1(ram[38]), .A2(n4395), .B1(n13558), .B2(n9019), .ZN(n4401) );
  INV_X1 U987 ( .A(n4402), .ZN(n13549) );
  AOI22_X1 U988 ( .A1(ram[39]), .A2(n4395), .B1(n13558), .B2(n9043), .ZN(n4402) );
  INV_X1 U989 ( .A(n4403), .ZN(n13550) );
  AOI22_X1 U990 ( .A1(ram[40]), .A2(n4395), .B1(n13558), .B2(n9067), .ZN(n4403) );
  INV_X1 U991 ( .A(n4404), .ZN(n13551) );
  AOI22_X1 U992 ( .A1(ram[41]), .A2(n4395), .B1(n13558), .B2(n9091), .ZN(n4404) );
  INV_X1 U993 ( .A(n4405), .ZN(n13552) );
  AOI22_X1 U994 ( .A1(ram[42]), .A2(n4395), .B1(n13558), .B2(n9115), .ZN(n4405) );
  INV_X1 U995 ( .A(n4406), .ZN(n13553) );
  AOI22_X1 U996 ( .A1(ram[43]), .A2(n4395), .B1(n13558), .B2(n9139), .ZN(n4406) );
  INV_X1 U997 ( .A(n4407), .ZN(n13554) );
  AOI22_X1 U998 ( .A1(ram[44]), .A2(n4395), .B1(n13558), .B2(n9163), .ZN(n4407) );
  INV_X1 U999 ( .A(n4408), .ZN(n13555) );
  AOI22_X1 U1000 ( .A1(ram[45]), .A2(n4395), .B1(n13558), .B2(n9187), .ZN(
        n4408) );
  INV_X1 U1001 ( .A(n4409), .ZN(n13556) );
  AOI22_X1 U1002 ( .A1(ram[46]), .A2(n4395), .B1(n13558), .B2(n9211), .ZN(
        n4409) );
  INV_X1 U1003 ( .A(n4410), .ZN(n13557) );
  AOI22_X1 U1004 ( .A1(ram[47]), .A2(n4395), .B1(n13558), .B2(n9235), .ZN(
        n4410) );
  INV_X1 U1005 ( .A(n4430), .ZN(n13508) );
  AOI22_X1 U1006 ( .A1(ram[64]), .A2(n4431), .B1(n13524), .B2(n8874), .ZN(
        n4430) );
  INV_X1 U1007 ( .A(n4432), .ZN(n13509) );
  AOI22_X1 U1008 ( .A1(ram[65]), .A2(n4431), .B1(n13524), .B2(n8898), .ZN(
        n4432) );
  INV_X1 U1009 ( .A(n4433), .ZN(n13510) );
  AOI22_X1 U1010 ( .A1(ram[66]), .A2(n4431), .B1(n13524), .B2(n8922), .ZN(
        n4433) );
  INV_X1 U1011 ( .A(n4434), .ZN(n13511) );
  AOI22_X1 U1012 ( .A1(ram[67]), .A2(n4431), .B1(n13524), .B2(n8946), .ZN(
        n4434) );
  INV_X1 U1013 ( .A(n4435), .ZN(n13512) );
  AOI22_X1 U1014 ( .A1(ram[68]), .A2(n4431), .B1(n13524), .B2(n8970), .ZN(
        n4435) );
  INV_X1 U1015 ( .A(n4436), .ZN(n13513) );
  AOI22_X1 U1016 ( .A1(ram[69]), .A2(n4431), .B1(n13524), .B2(n8994), .ZN(
        n4436) );
  INV_X1 U1017 ( .A(n4437), .ZN(n13514) );
  AOI22_X1 U1018 ( .A1(ram[70]), .A2(n4431), .B1(n13524), .B2(n9018), .ZN(
        n4437) );
  INV_X1 U1019 ( .A(n4438), .ZN(n13515) );
  AOI22_X1 U1020 ( .A1(ram[71]), .A2(n4431), .B1(n13524), .B2(n9042), .ZN(
        n4438) );
  INV_X1 U1021 ( .A(n4439), .ZN(n13516) );
  AOI22_X1 U1022 ( .A1(ram[72]), .A2(n4431), .B1(n13524), .B2(n9066), .ZN(
        n4439) );
  INV_X1 U1023 ( .A(n4440), .ZN(n13517) );
  AOI22_X1 U1024 ( .A1(ram[73]), .A2(n4431), .B1(n13524), .B2(n9090), .ZN(
        n4440) );
  INV_X1 U1025 ( .A(n4441), .ZN(n13518) );
  AOI22_X1 U1026 ( .A1(ram[74]), .A2(n4431), .B1(n13524), .B2(n9114), .ZN(
        n4441) );
  INV_X1 U1027 ( .A(n4442), .ZN(n13519) );
  AOI22_X1 U1028 ( .A1(ram[75]), .A2(n4431), .B1(n13524), .B2(n9138), .ZN(
        n4442) );
  INV_X1 U1029 ( .A(n4443), .ZN(n13520) );
  AOI22_X1 U1030 ( .A1(ram[76]), .A2(n4431), .B1(n13524), .B2(n9162), .ZN(
        n4443) );
  INV_X1 U1031 ( .A(n4444), .ZN(n13521) );
  AOI22_X1 U1032 ( .A1(ram[77]), .A2(n4431), .B1(n13524), .B2(n9186), .ZN(
        n4444) );
  INV_X1 U1033 ( .A(n4445), .ZN(n13522) );
  AOI22_X1 U1034 ( .A1(ram[78]), .A2(n4431), .B1(n13524), .B2(n9210), .ZN(
        n4445) );
  INV_X1 U1035 ( .A(n4446), .ZN(n13523) );
  AOI22_X1 U1036 ( .A1(ram[79]), .A2(n4431), .B1(n13524), .B2(n9234), .ZN(
        n4446) );
  INV_X1 U1037 ( .A(n4466), .ZN(n13474) );
  AOI22_X1 U1038 ( .A1(ram[96]), .A2(n4467), .B1(n13490), .B2(n8874), .ZN(
        n4466) );
  INV_X1 U1039 ( .A(n4468), .ZN(n13475) );
  AOI22_X1 U1040 ( .A1(ram[97]), .A2(n4467), .B1(n13490), .B2(n8898), .ZN(
        n4468) );
  INV_X1 U1041 ( .A(n4469), .ZN(n13476) );
  AOI22_X1 U1042 ( .A1(ram[98]), .A2(n4467), .B1(n13490), .B2(n8922), .ZN(
        n4469) );
  INV_X1 U1043 ( .A(n4470), .ZN(n13477) );
  AOI22_X1 U1044 ( .A1(ram[99]), .A2(n4467), .B1(n13490), .B2(n8946), .ZN(
        n4470) );
  INV_X1 U1045 ( .A(n4471), .ZN(n13478) );
  AOI22_X1 U1046 ( .A1(ram[100]), .A2(n4467), .B1(n13490), .B2(n8970), .ZN(
        n4471) );
  INV_X1 U1047 ( .A(n4472), .ZN(n13479) );
  AOI22_X1 U1048 ( .A1(ram[101]), .A2(n4467), .B1(n13490), .B2(n8994), .ZN(
        n4472) );
  INV_X1 U1049 ( .A(n4473), .ZN(n13480) );
  AOI22_X1 U1050 ( .A1(ram[102]), .A2(n4467), .B1(n13490), .B2(n9018), .ZN(
        n4473) );
  INV_X1 U1051 ( .A(n4474), .ZN(n13481) );
  AOI22_X1 U1052 ( .A1(ram[103]), .A2(n4467), .B1(n13490), .B2(n9042), .ZN(
        n4474) );
  INV_X1 U1053 ( .A(n4475), .ZN(n13482) );
  AOI22_X1 U1054 ( .A1(ram[104]), .A2(n4467), .B1(n13490), .B2(n9066), .ZN(
        n4475) );
  INV_X1 U1055 ( .A(n4476), .ZN(n13483) );
  AOI22_X1 U1056 ( .A1(ram[105]), .A2(n4467), .B1(n13490), .B2(n9090), .ZN(
        n4476) );
  INV_X1 U1057 ( .A(n4477), .ZN(n13484) );
  AOI22_X1 U1058 ( .A1(ram[106]), .A2(n4467), .B1(n13490), .B2(n9114), .ZN(
        n4477) );
  INV_X1 U1059 ( .A(n4478), .ZN(n13485) );
  AOI22_X1 U1060 ( .A1(ram[107]), .A2(n4467), .B1(n13490), .B2(n9138), .ZN(
        n4478) );
  INV_X1 U1061 ( .A(n4479), .ZN(n13486) );
  AOI22_X1 U1062 ( .A1(ram[108]), .A2(n4467), .B1(n13490), .B2(n9162), .ZN(
        n4479) );
  INV_X1 U1063 ( .A(n4480), .ZN(n13487) );
  AOI22_X1 U1064 ( .A1(ram[109]), .A2(n4467), .B1(n13490), .B2(n9186), .ZN(
        n4480) );
  INV_X1 U1065 ( .A(n4481), .ZN(n13488) );
  AOI22_X1 U1066 ( .A1(ram[110]), .A2(n4467), .B1(n13490), .B2(n9210), .ZN(
        n4481) );
  INV_X1 U1067 ( .A(n4482), .ZN(n13489) );
  AOI22_X1 U1068 ( .A1(ram[111]), .A2(n4467), .B1(n13490), .B2(n9234), .ZN(
        n4482) );
  INV_X1 U1069 ( .A(n4502), .ZN(n13440) );
  AOI22_X1 U1070 ( .A1(ram[128]), .A2(n4503), .B1(n13456), .B2(n8874), .ZN(
        n4502) );
  INV_X1 U1071 ( .A(n4504), .ZN(n13441) );
  AOI22_X1 U1072 ( .A1(ram[129]), .A2(n4503), .B1(n13456), .B2(n8898), .ZN(
        n4504) );
  INV_X1 U1073 ( .A(n4505), .ZN(n13442) );
  AOI22_X1 U1074 ( .A1(ram[130]), .A2(n4503), .B1(n13456), .B2(n8922), .ZN(
        n4505) );
  INV_X1 U1075 ( .A(n4506), .ZN(n13443) );
  AOI22_X1 U1076 ( .A1(ram[131]), .A2(n4503), .B1(n13456), .B2(n8946), .ZN(
        n4506) );
  INV_X1 U1077 ( .A(n4507), .ZN(n13444) );
  AOI22_X1 U1078 ( .A1(ram[132]), .A2(n4503), .B1(n13456), .B2(n8970), .ZN(
        n4507) );
  INV_X1 U1079 ( .A(n4508), .ZN(n13445) );
  AOI22_X1 U1080 ( .A1(ram[133]), .A2(n4503), .B1(n13456), .B2(n8994), .ZN(
        n4508) );
  INV_X1 U1081 ( .A(n4509), .ZN(n13446) );
  AOI22_X1 U1082 ( .A1(ram[134]), .A2(n4503), .B1(n13456), .B2(n9018), .ZN(
        n4509) );
  INV_X1 U1083 ( .A(n4510), .ZN(n13447) );
  AOI22_X1 U1084 ( .A1(ram[135]), .A2(n4503), .B1(n13456), .B2(n9042), .ZN(
        n4510) );
  INV_X1 U1085 ( .A(n4511), .ZN(n13448) );
  AOI22_X1 U1086 ( .A1(ram[136]), .A2(n4503), .B1(n13456), .B2(n9066), .ZN(
        n4511) );
  INV_X1 U1087 ( .A(n4512), .ZN(n13449) );
  AOI22_X1 U1088 ( .A1(ram[137]), .A2(n4503), .B1(n13456), .B2(n9090), .ZN(
        n4512) );
  INV_X1 U1089 ( .A(n4513), .ZN(n13450) );
  AOI22_X1 U1090 ( .A1(ram[138]), .A2(n4503), .B1(n13456), .B2(n9114), .ZN(
        n4513) );
  INV_X1 U1091 ( .A(n4514), .ZN(n13451) );
  AOI22_X1 U1092 ( .A1(ram[139]), .A2(n4503), .B1(n13456), .B2(n9138), .ZN(
        n4514) );
  INV_X1 U1093 ( .A(n4515), .ZN(n13452) );
  AOI22_X1 U1094 ( .A1(ram[140]), .A2(n4503), .B1(n13456), .B2(n9162), .ZN(
        n4515) );
  INV_X1 U1095 ( .A(n4516), .ZN(n13453) );
  AOI22_X1 U1096 ( .A1(ram[141]), .A2(n4503), .B1(n13456), .B2(n9186), .ZN(
        n4516) );
  INV_X1 U1097 ( .A(n4517), .ZN(n13454) );
  AOI22_X1 U1098 ( .A1(ram[142]), .A2(n4503), .B1(n13456), .B2(n9210), .ZN(
        n4517) );
  INV_X1 U1099 ( .A(n4518), .ZN(n13455) );
  AOI22_X1 U1100 ( .A1(ram[143]), .A2(n4503), .B1(n13456), .B2(n9234), .ZN(
        n4518) );
  INV_X1 U1101 ( .A(n4538), .ZN(n13406) );
  AOI22_X1 U1102 ( .A1(ram[160]), .A2(n4539), .B1(n13422), .B2(n8874), .ZN(
        n4538) );
  INV_X1 U1103 ( .A(n4540), .ZN(n13407) );
  AOI22_X1 U1104 ( .A1(ram[161]), .A2(n4539), .B1(n13422), .B2(n8898), .ZN(
        n4540) );
  INV_X1 U1105 ( .A(n4541), .ZN(n13408) );
  AOI22_X1 U1106 ( .A1(ram[162]), .A2(n4539), .B1(n13422), .B2(n8922), .ZN(
        n4541) );
  INV_X1 U1107 ( .A(n4542), .ZN(n13409) );
  AOI22_X1 U1108 ( .A1(ram[163]), .A2(n4539), .B1(n13422), .B2(n8946), .ZN(
        n4542) );
  INV_X1 U1109 ( .A(n4543), .ZN(n13410) );
  AOI22_X1 U1110 ( .A1(ram[164]), .A2(n4539), .B1(n13422), .B2(n8970), .ZN(
        n4543) );
  INV_X1 U1111 ( .A(n4544), .ZN(n13411) );
  AOI22_X1 U1112 ( .A1(ram[165]), .A2(n4539), .B1(n13422), .B2(n8994), .ZN(
        n4544) );
  INV_X1 U1113 ( .A(n4545), .ZN(n13412) );
  AOI22_X1 U1114 ( .A1(ram[166]), .A2(n4539), .B1(n13422), .B2(n9018), .ZN(
        n4545) );
  INV_X1 U1115 ( .A(n4546), .ZN(n13413) );
  AOI22_X1 U1116 ( .A1(ram[167]), .A2(n4539), .B1(n13422), .B2(n9042), .ZN(
        n4546) );
  INV_X1 U1117 ( .A(n4547), .ZN(n13414) );
  AOI22_X1 U1118 ( .A1(ram[168]), .A2(n4539), .B1(n13422), .B2(n9066), .ZN(
        n4547) );
  INV_X1 U1119 ( .A(n4548), .ZN(n13415) );
  AOI22_X1 U1120 ( .A1(ram[169]), .A2(n4539), .B1(n13422), .B2(n9090), .ZN(
        n4548) );
  INV_X1 U1121 ( .A(n4549), .ZN(n13416) );
  AOI22_X1 U1122 ( .A1(ram[170]), .A2(n4539), .B1(n13422), .B2(n9114), .ZN(
        n4549) );
  INV_X1 U1123 ( .A(n4550), .ZN(n13417) );
  AOI22_X1 U1124 ( .A1(ram[171]), .A2(n4539), .B1(n13422), .B2(n9138), .ZN(
        n4550) );
  INV_X1 U1125 ( .A(n4551), .ZN(n13418) );
  AOI22_X1 U1126 ( .A1(ram[172]), .A2(n4539), .B1(n13422), .B2(n9162), .ZN(
        n4551) );
  INV_X1 U1127 ( .A(n4552), .ZN(n13419) );
  AOI22_X1 U1128 ( .A1(ram[173]), .A2(n4539), .B1(n13422), .B2(n9186), .ZN(
        n4552) );
  INV_X1 U1129 ( .A(n4553), .ZN(n13420) );
  AOI22_X1 U1130 ( .A1(ram[174]), .A2(n4539), .B1(n13422), .B2(n9210), .ZN(
        n4553) );
  INV_X1 U1131 ( .A(n4554), .ZN(n13421) );
  AOI22_X1 U1132 ( .A1(ram[175]), .A2(n4539), .B1(n13422), .B2(n9234), .ZN(
        n4554) );
  INV_X1 U1133 ( .A(n4574), .ZN(n13372) );
  AOI22_X1 U1134 ( .A1(ram[192]), .A2(n4575), .B1(n13388), .B2(n8874), .ZN(
        n4574) );
  INV_X1 U1135 ( .A(n4576), .ZN(n13373) );
  AOI22_X1 U1136 ( .A1(ram[193]), .A2(n4575), .B1(n13388), .B2(n8898), .ZN(
        n4576) );
  INV_X1 U1137 ( .A(n4577), .ZN(n13374) );
  AOI22_X1 U1138 ( .A1(ram[194]), .A2(n4575), .B1(n13388), .B2(n8922), .ZN(
        n4577) );
  INV_X1 U1139 ( .A(n4578), .ZN(n13375) );
  AOI22_X1 U1140 ( .A1(ram[195]), .A2(n4575), .B1(n13388), .B2(n8946), .ZN(
        n4578) );
  INV_X1 U1141 ( .A(n4579), .ZN(n13376) );
  AOI22_X1 U1142 ( .A1(ram[196]), .A2(n4575), .B1(n13388), .B2(n8970), .ZN(
        n4579) );
  INV_X1 U1143 ( .A(n4580), .ZN(n13377) );
  AOI22_X1 U1144 ( .A1(ram[197]), .A2(n4575), .B1(n13388), .B2(n8994), .ZN(
        n4580) );
  INV_X1 U1145 ( .A(n4581), .ZN(n13378) );
  AOI22_X1 U1146 ( .A1(ram[198]), .A2(n4575), .B1(n13388), .B2(n9018), .ZN(
        n4581) );
  INV_X1 U1147 ( .A(n4582), .ZN(n13379) );
  AOI22_X1 U1148 ( .A1(ram[199]), .A2(n4575), .B1(n13388), .B2(n9042), .ZN(
        n4582) );
  INV_X1 U1149 ( .A(n4583), .ZN(n13380) );
  AOI22_X1 U1150 ( .A1(ram[200]), .A2(n4575), .B1(n13388), .B2(n9066), .ZN(
        n4583) );
  INV_X1 U1151 ( .A(n4584), .ZN(n13381) );
  AOI22_X1 U1152 ( .A1(ram[201]), .A2(n4575), .B1(n13388), .B2(n9090), .ZN(
        n4584) );
  INV_X1 U1153 ( .A(n4585), .ZN(n13382) );
  AOI22_X1 U1154 ( .A1(ram[202]), .A2(n4575), .B1(n13388), .B2(n9114), .ZN(
        n4585) );
  INV_X1 U1155 ( .A(n4586), .ZN(n13383) );
  AOI22_X1 U1156 ( .A1(ram[203]), .A2(n4575), .B1(n13388), .B2(n9138), .ZN(
        n4586) );
  INV_X1 U1157 ( .A(n4587), .ZN(n13384) );
  AOI22_X1 U1158 ( .A1(ram[204]), .A2(n4575), .B1(n13388), .B2(n9162), .ZN(
        n4587) );
  INV_X1 U1159 ( .A(n4588), .ZN(n13385) );
  AOI22_X1 U1160 ( .A1(ram[205]), .A2(n4575), .B1(n13388), .B2(n9186), .ZN(
        n4588) );
  INV_X1 U1161 ( .A(n4589), .ZN(n13386) );
  AOI22_X1 U1162 ( .A1(ram[206]), .A2(n4575), .B1(n13388), .B2(n9210), .ZN(
        n4589) );
  INV_X1 U1163 ( .A(n4590), .ZN(n13387) );
  AOI22_X1 U1164 ( .A1(ram[207]), .A2(n4575), .B1(n13388), .B2(n9234), .ZN(
        n4590) );
  INV_X1 U1165 ( .A(n4610), .ZN(n13338) );
  AOI22_X1 U1166 ( .A1(ram[224]), .A2(n4611), .B1(n13354), .B2(n8874), .ZN(
        n4610) );
  INV_X1 U1167 ( .A(n4612), .ZN(n13339) );
  AOI22_X1 U1168 ( .A1(ram[225]), .A2(n4611), .B1(n13354), .B2(n8898), .ZN(
        n4612) );
  INV_X1 U1169 ( .A(n4613), .ZN(n13340) );
  AOI22_X1 U1170 ( .A1(ram[226]), .A2(n4611), .B1(n13354), .B2(n8922), .ZN(
        n4613) );
  INV_X1 U1171 ( .A(n4614), .ZN(n13341) );
  AOI22_X1 U1172 ( .A1(ram[227]), .A2(n4611), .B1(n13354), .B2(n8946), .ZN(
        n4614) );
  INV_X1 U1173 ( .A(n4615), .ZN(n13342) );
  AOI22_X1 U1174 ( .A1(ram[228]), .A2(n4611), .B1(n13354), .B2(n8970), .ZN(
        n4615) );
  INV_X1 U1175 ( .A(n4616), .ZN(n13343) );
  AOI22_X1 U1176 ( .A1(ram[229]), .A2(n4611), .B1(n13354), .B2(n8994), .ZN(
        n4616) );
  INV_X1 U1177 ( .A(n4617), .ZN(n13344) );
  AOI22_X1 U1178 ( .A1(ram[230]), .A2(n4611), .B1(n13354), .B2(n9018), .ZN(
        n4617) );
  INV_X1 U1179 ( .A(n4618), .ZN(n13345) );
  AOI22_X1 U1180 ( .A1(ram[231]), .A2(n4611), .B1(n13354), .B2(n9042), .ZN(
        n4618) );
  INV_X1 U1181 ( .A(n4619), .ZN(n13346) );
  AOI22_X1 U1182 ( .A1(ram[232]), .A2(n4611), .B1(n13354), .B2(n9066), .ZN(
        n4619) );
  INV_X1 U1183 ( .A(n4620), .ZN(n13347) );
  AOI22_X1 U1184 ( .A1(ram[233]), .A2(n4611), .B1(n13354), .B2(n9090), .ZN(
        n4620) );
  INV_X1 U1185 ( .A(n4621), .ZN(n13348) );
  AOI22_X1 U1186 ( .A1(ram[234]), .A2(n4611), .B1(n13354), .B2(n9114), .ZN(
        n4621) );
  INV_X1 U1187 ( .A(n4622), .ZN(n13349) );
  AOI22_X1 U1188 ( .A1(ram[235]), .A2(n4611), .B1(n13354), .B2(n9138), .ZN(
        n4622) );
  INV_X1 U1189 ( .A(n4623), .ZN(n13350) );
  AOI22_X1 U1190 ( .A1(ram[236]), .A2(n4611), .B1(n13354), .B2(n9162), .ZN(
        n4623) );
  INV_X1 U1191 ( .A(n4624), .ZN(n13351) );
  AOI22_X1 U1192 ( .A1(ram[237]), .A2(n4611), .B1(n13354), .B2(n9186), .ZN(
        n4624) );
  INV_X1 U1193 ( .A(n4625), .ZN(n13352) );
  AOI22_X1 U1194 ( .A1(ram[238]), .A2(n4611), .B1(n13354), .B2(n9210), .ZN(
        n4625) );
  INV_X1 U1195 ( .A(n4626), .ZN(n13353) );
  AOI22_X1 U1196 ( .A1(ram[239]), .A2(n4611), .B1(n13354), .B2(n9234), .ZN(
        n4626) );
  INV_X1 U1197 ( .A(n4648), .ZN(n13304) );
  AOI22_X1 U1198 ( .A1(ram[256]), .A2(n4649), .B1(n13320), .B2(n8873), .ZN(
        n4648) );
  INV_X1 U1199 ( .A(n4650), .ZN(n13305) );
  AOI22_X1 U1200 ( .A1(ram[257]), .A2(n4649), .B1(n13320), .B2(n8897), .ZN(
        n4650) );
  INV_X1 U1201 ( .A(n4651), .ZN(n13306) );
  AOI22_X1 U1202 ( .A1(ram[258]), .A2(n4649), .B1(n13320), .B2(n8921), .ZN(
        n4651) );
  INV_X1 U1203 ( .A(n4652), .ZN(n13307) );
  AOI22_X1 U1204 ( .A1(ram[259]), .A2(n4649), .B1(n13320), .B2(n8945), .ZN(
        n4652) );
  INV_X1 U1205 ( .A(n4653), .ZN(n13308) );
  AOI22_X1 U1206 ( .A1(ram[260]), .A2(n4649), .B1(n13320), .B2(n8969), .ZN(
        n4653) );
  INV_X1 U1207 ( .A(n4654), .ZN(n13309) );
  AOI22_X1 U1208 ( .A1(ram[261]), .A2(n4649), .B1(n13320), .B2(n8993), .ZN(
        n4654) );
  INV_X1 U1209 ( .A(n4655), .ZN(n13310) );
  AOI22_X1 U1210 ( .A1(ram[262]), .A2(n4649), .B1(n13320), .B2(n9017), .ZN(
        n4655) );
  INV_X1 U1211 ( .A(n4656), .ZN(n13311) );
  AOI22_X1 U1212 ( .A1(ram[263]), .A2(n4649), .B1(n13320), .B2(n9041), .ZN(
        n4656) );
  INV_X1 U1213 ( .A(n4657), .ZN(n13312) );
  AOI22_X1 U1214 ( .A1(ram[264]), .A2(n4649), .B1(n13320), .B2(n9065), .ZN(
        n4657) );
  INV_X1 U1215 ( .A(n4658), .ZN(n13313) );
  AOI22_X1 U1216 ( .A1(ram[265]), .A2(n4649), .B1(n13320), .B2(n9089), .ZN(
        n4658) );
  INV_X1 U1217 ( .A(n4659), .ZN(n13314) );
  AOI22_X1 U1218 ( .A1(ram[266]), .A2(n4649), .B1(n13320), .B2(n9113), .ZN(
        n4659) );
  INV_X1 U1219 ( .A(n4660), .ZN(n13315) );
  AOI22_X1 U1220 ( .A1(ram[267]), .A2(n4649), .B1(n13320), .B2(n9137), .ZN(
        n4660) );
  INV_X1 U1221 ( .A(n4661), .ZN(n13316) );
  AOI22_X1 U1222 ( .A1(ram[268]), .A2(n4649), .B1(n13320), .B2(n9161), .ZN(
        n4661) );
  INV_X1 U1223 ( .A(n4662), .ZN(n13317) );
  AOI22_X1 U1224 ( .A1(ram[269]), .A2(n4649), .B1(n13320), .B2(n9185), .ZN(
        n4662) );
  INV_X1 U1225 ( .A(n4663), .ZN(n13318) );
  AOI22_X1 U1226 ( .A1(ram[270]), .A2(n4649), .B1(n13320), .B2(n9209), .ZN(
        n4663) );
  INV_X1 U1227 ( .A(n4664), .ZN(n13319) );
  AOI22_X1 U1228 ( .A1(ram[271]), .A2(n4649), .B1(n13320), .B2(n9233), .ZN(
        n4664) );
  INV_X1 U1229 ( .A(n4683), .ZN(n13270) );
  AOI22_X1 U1230 ( .A1(ram[288]), .A2(n4684), .B1(n13286), .B2(n8873), .ZN(
        n4683) );
  INV_X1 U1231 ( .A(n4685), .ZN(n13271) );
  AOI22_X1 U1232 ( .A1(ram[289]), .A2(n4684), .B1(n13286), .B2(n8897), .ZN(
        n4685) );
  INV_X1 U1233 ( .A(n4686), .ZN(n13272) );
  AOI22_X1 U1234 ( .A1(ram[290]), .A2(n4684), .B1(n13286), .B2(n8921), .ZN(
        n4686) );
  INV_X1 U1235 ( .A(n4687), .ZN(n13273) );
  AOI22_X1 U1236 ( .A1(ram[291]), .A2(n4684), .B1(n13286), .B2(n8945), .ZN(
        n4687) );
  INV_X1 U1237 ( .A(n4688), .ZN(n13274) );
  AOI22_X1 U1238 ( .A1(ram[292]), .A2(n4684), .B1(n13286), .B2(n8969), .ZN(
        n4688) );
  INV_X1 U1239 ( .A(n4689), .ZN(n13275) );
  AOI22_X1 U1240 ( .A1(ram[293]), .A2(n4684), .B1(n13286), .B2(n8993), .ZN(
        n4689) );
  INV_X1 U1241 ( .A(n4690), .ZN(n13276) );
  AOI22_X1 U1242 ( .A1(ram[294]), .A2(n4684), .B1(n13286), .B2(n9017), .ZN(
        n4690) );
  INV_X1 U1243 ( .A(n4691), .ZN(n13277) );
  AOI22_X1 U1244 ( .A1(ram[295]), .A2(n4684), .B1(n13286), .B2(n9041), .ZN(
        n4691) );
  INV_X1 U1245 ( .A(n4692), .ZN(n13278) );
  AOI22_X1 U1246 ( .A1(ram[296]), .A2(n4684), .B1(n13286), .B2(n9065), .ZN(
        n4692) );
  INV_X1 U1247 ( .A(n4693), .ZN(n13279) );
  AOI22_X1 U1248 ( .A1(ram[297]), .A2(n4684), .B1(n13286), .B2(n9089), .ZN(
        n4693) );
  INV_X1 U1249 ( .A(n4694), .ZN(n13280) );
  AOI22_X1 U1250 ( .A1(ram[298]), .A2(n4684), .B1(n13286), .B2(n9113), .ZN(
        n4694) );
  INV_X1 U1251 ( .A(n4695), .ZN(n13281) );
  AOI22_X1 U1252 ( .A1(ram[299]), .A2(n4684), .B1(n13286), .B2(n9137), .ZN(
        n4695) );
  INV_X1 U1253 ( .A(n4696), .ZN(n13282) );
  AOI22_X1 U1254 ( .A1(ram[300]), .A2(n4684), .B1(n13286), .B2(n9161), .ZN(
        n4696) );
  INV_X1 U1255 ( .A(n4697), .ZN(n13283) );
  AOI22_X1 U1256 ( .A1(ram[301]), .A2(n4684), .B1(n13286), .B2(n9185), .ZN(
        n4697) );
  INV_X1 U1257 ( .A(n4698), .ZN(n13284) );
  AOI22_X1 U1258 ( .A1(ram[302]), .A2(n4684), .B1(n13286), .B2(n9209), .ZN(
        n4698) );
  INV_X1 U1259 ( .A(n4699), .ZN(n13285) );
  AOI22_X1 U1260 ( .A1(ram[303]), .A2(n4684), .B1(n13286), .B2(n9233), .ZN(
        n4699) );
  INV_X1 U1261 ( .A(n4717), .ZN(n13236) );
  AOI22_X1 U1262 ( .A1(ram[320]), .A2(n4718), .B1(n13252), .B2(n8873), .ZN(
        n4717) );
  INV_X1 U1263 ( .A(n4719), .ZN(n13237) );
  AOI22_X1 U1264 ( .A1(ram[321]), .A2(n4718), .B1(n13252), .B2(n8897), .ZN(
        n4719) );
  INV_X1 U1265 ( .A(n4720), .ZN(n13238) );
  AOI22_X1 U1266 ( .A1(ram[322]), .A2(n4718), .B1(n13252), .B2(n8921), .ZN(
        n4720) );
  INV_X1 U1267 ( .A(n4721), .ZN(n13239) );
  AOI22_X1 U1268 ( .A1(ram[323]), .A2(n4718), .B1(n13252), .B2(n8945), .ZN(
        n4721) );
  INV_X1 U1269 ( .A(n4722), .ZN(n13240) );
  AOI22_X1 U1270 ( .A1(ram[324]), .A2(n4718), .B1(n13252), .B2(n8969), .ZN(
        n4722) );
  INV_X1 U1271 ( .A(n4723), .ZN(n13241) );
  AOI22_X1 U1272 ( .A1(ram[325]), .A2(n4718), .B1(n13252), .B2(n8993), .ZN(
        n4723) );
  INV_X1 U1273 ( .A(n4724), .ZN(n13242) );
  AOI22_X1 U1274 ( .A1(ram[326]), .A2(n4718), .B1(n13252), .B2(n9017), .ZN(
        n4724) );
  INV_X1 U1275 ( .A(n4725), .ZN(n13243) );
  AOI22_X1 U1276 ( .A1(ram[327]), .A2(n4718), .B1(n13252), .B2(n9041), .ZN(
        n4725) );
  INV_X1 U1277 ( .A(n4726), .ZN(n13244) );
  AOI22_X1 U1278 ( .A1(ram[328]), .A2(n4718), .B1(n13252), .B2(n9065), .ZN(
        n4726) );
  INV_X1 U1279 ( .A(n4727), .ZN(n13245) );
  AOI22_X1 U1280 ( .A1(ram[329]), .A2(n4718), .B1(n13252), .B2(n9089), .ZN(
        n4727) );
  INV_X1 U1281 ( .A(n4728), .ZN(n13246) );
  AOI22_X1 U1282 ( .A1(ram[330]), .A2(n4718), .B1(n13252), .B2(n9113), .ZN(
        n4728) );
  INV_X1 U1283 ( .A(n4729), .ZN(n13247) );
  AOI22_X1 U1284 ( .A1(ram[331]), .A2(n4718), .B1(n13252), .B2(n9137), .ZN(
        n4729) );
  INV_X1 U1285 ( .A(n4730), .ZN(n13248) );
  AOI22_X1 U1286 ( .A1(ram[332]), .A2(n4718), .B1(n13252), .B2(n9161), .ZN(
        n4730) );
  INV_X1 U1287 ( .A(n4731), .ZN(n13249) );
  AOI22_X1 U1288 ( .A1(ram[333]), .A2(n4718), .B1(n13252), .B2(n9185), .ZN(
        n4731) );
  INV_X1 U1289 ( .A(n4732), .ZN(n13250) );
  AOI22_X1 U1290 ( .A1(ram[334]), .A2(n4718), .B1(n13252), .B2(n9209), .ZN(
        n4732) );
  INV_X1 U1291 ( .A(n4733), .ZN(n13251) );
  AOI22_X1 U1292 ( .A1(ram[335]), .A2(n4718), .B1(n13252), .B2(n9233), .ZN(
        n4733) );
  INV_X1 U1293 ( .A(n4751), .ZN(n13202) );
  AOI22_X1 U1294 ( .A1(ram[352]), .A2(n4752), .B1(n13218), .B2(n8873), .ZN(
        n4751) );
  INV_X1 U1295 ( .A(n4753), .ZN(n13203) );
  AOI22_X1 U1296 ( .A1(ram[353]), .A2(n4752), .B1(n13218), .B2(n8897), .ZN(
        n4753) );
  INV_X1 U1297 ( .A(n4754), .ZN(n13204) );
  AOI22_X1 U1298 ( .A1(ram[354]), .A2(n4752), .B1(n13218), .B2(n8921), .ZN(
        n4754) );
  INV_X1 U1299 ( .A(n4755), .ZN(n13205) );
  AOI22_X1 U1300 ( .A1(ram[355]), .A2(n4752), .B1(n13218), .B2(n8945), .ZN(
        n4755) );
  INV_X1 U1301 ( .A(n4756), .ZN(n13206) );
  AOI22_X1 U1302 ( .A1(ram[356]), .A2(n4752), .B1(n13218), .B2(n8969), .ZN(
        n4756) );
  INV_X1 U1303 ( .A(n4757), .ZN(n13207) );
  AOI22_X1 U1304 ( .A1(ram[357]), .A2(n4752), .B1(n13218), .B2(n8993), .ZN(
        n4757) );
  INV_X1 U1305 ( .A(n4758), .ZN(n13208) );
  AOI22_X1 U1306 ( .A1(ram[358]), .A2(n4752), .B1(n13218), .B2(n9017), .ZN(
        n4758) );
  INV_X1 U1307 ( .A(n4759), .ZN(n13209) );
  AOI22_X1 U1308 ( .A1(ram[359]), .A2(n4752), .B1(n13218), .B2(n9041), .ZN(
        n4759) );
  INV_X1 U1309 ( .A(n4760), .ZN(n13210) );
  AOI22_X1 U1310 ( .A1(ram[360]), .A2(n4752), .B1(n13218), .B2(n9065), .ZN(
        n4760) );
  INV_X1 U1311 ( .A(n4761), .ZN(n13211) );
  AOI22_X1 U1312 ( .A1(ram[361]), .A2(n4752), .B1(n13218), .B2(n9089), .ZN(
        n4761) );
  INV_X1 U1313 ( .A(n4762), .ZN(n13212) );
  AOI22_X1 U1314 ( .A1(ram[362]), .A2(n4752), .B1(n13218), .B2(n9113), .ZN(
        n4762) );
  INV_X1 U1315 ( .A(n4763), .ZN(n13213) );
  AOI22_X1 U1316 ( .A1(ram[363]), .A2(n4752), .B1(n13218), .B2(n9137), .ZN(
        n4763) );
  INV_X1 U1317 ( .A(n4764), .ZN(n13214) );
  AOI22_X1 U1318 ( .A1(ram[364]), .A2(n4752), .B1(n13218), .B2(n9161), .ZN(
        n4764) );
  INV_X1 U1319 ( .A(n4765), .ZN(n13215) );
  AOI22_X1 U1320 ( .A1(ram[365]), .A2(n4752), .B1(n13218), .B2(n9185), .ZN(
        n4765) );
  INV_X1 U1321 ( .A(n4766), .ZN(n13216) );
  AOI22_X1 U1322 ( .A1(ram[366]), .A2(n4752), .B1(n13218), .B2(n9209), .ZN(
        n4766) );
  INV_X1 U1323 ( .A(n4767), .ZN(n13217) );
  AOI22_X1 U1324 ( .A1(ram[367]), .A2(n4752), .B1(n13218), .B2(n9233), .ZN(
        n4767) );
  INV_X1 U1325 ( .A(n4785), .ZN(n13168) );
  AOI22_X1 U1326 ( .A1(ram[384]), .A2(n4786), .B1(n13184), .B2(n8873), .ZN(
        n4785) );
  INV_X1 U1327 ( .A(n4787), .ZN(n13169) );
  AOI22_X1 U1328 ( .A1(ram[385]), .A2(n4786), .B1(n13184), .B2(n8897), .ZN(
        n4787) );
  INV_X1 U1329 ( .A(n4788), .ZN(n13170) );
  AOI22_X1 U1330 ( .A1(ram[386]), .A2(n4786), .B1(n13184), .B2(n8921), .ZN(
        n4788) );
  INV_X1 U1331 ( .A(n4789), .ZN(n13171) );
  AOI22_X1 U1332 ( .A1(ram[387]), .A2(n4786), .B1(n13184), .B2(n8945), .ZN(
        n4789) );
  INV_X1 U1333 ( .A(n4790), .ZN(n13172) );
  AOI22_X1 U1334 ( .A1(ram[388]), .A2(n4786), .B1(n13184), .B2(n8969), .ZN(
        n4790) );
  INV_X1 U1335 ( .A(n4791), .ZN(n13173) );
  AOI22_X1 U1336 ( .A1(ram[389]), .A2(n4786), .B1(n13184), .B2(n8993), .ZN(
        n4791) );
  INV_X1 U1337 ( .A(n4792), .ZN(n13174) );
  AOI22_X1 U1338 ( .A1(ram[390]), .A2(n4786), .B1(n13184), .B2(n9017), .ZN(
        n4792) );
  INV_X1 U1339 ( .A(n4793), .ZN(n13175) );
  AOI22_X1 U1340 ( .A1(ram[391]), .A2(n4786), .B1(n13184), .B2(n9041), .ZN(
        n4793) );
  INV_X1 U1341 ( .A(n4794), .ZN(n13176) );
  AOI22_X1 U1342 ( .A1(ram[392]), .A2(n4786), .B1(n13184), .B2(n9065), .ZN(
        n4794) );
  INV_X1 U1343 ( .A(n4795), .ZN(n13177) );
  AOI22_X1 U1344 ( .A1(ram[393]), .A2(n4786), .B1(n13184), .B2(n9089), .ZN(
        n4795) );
  INV_X1 U1345 ( .A(n4796), .ZN(n13178) );
  AOI22_X1 U1346 ( .A1(ram[394]), .A2(n4786), .B1(n13184), .B2(n9113), .ZN(
        n4796) );
  INV_X1 U1347 ( .A(n4797), .ZN(n13179) );
  AOI22_X1 U1348 ( .A1(ram[395]), .A2(n4786), .B1(n13184), .B2(n9137), .ZN(
        n4797) );
  INV_X1 U1349 ( .A(n4798), .ZN(n13180) );
  AOI22_X1 U1350 ( .A1(ram[396]), .A2(n4786), .B1(n13184), .B2(n9161), .ZN(
        n4798) );
  INV_X1 U1351 ( .A(n4799), .ZN(n13181) );
  AOI22_X1 U1352 ( .A1(ram[397]), .A2(n4786), .B1(n13184), .B2(n9185), .ZN(
        n4799) );
  INV_X1 U1353 ( .A(n4800), .ZN(n13182) );
  AOI22_X1 U1354 ( .A1(ram[398]), .A2(n4786), .B1(n13184), .B2(n9209), .ZN(
        n4800) );
  INV_X1 U1355 ( .A(n4801), .ZN(n13183) );
  AOI22_X1 U1356 ( .A1(ram[399]), .A2(n4786), .B1(n13184), .B2(n9233), .ZN(
        n4801) );
  INV_X1 U1357 ( .A(n4819), .ZN(n13134) );
  AOI22_X1 U1358 ( .A1(ram[416]), .A2(n4820), .B1(n13150), .B2(n8873), .ZN(
        n4819) );
  INV_X1 U1359 ( .A(n4821), .ZN(n13135) );
  AOI22_X1 U1360 ( .A1(ram[417]), .A2(n4820), .B1(n13150), .B2(n8897), .ZN(
        n4821) );
  INV_X1 U1361 ( .A(n4822), .ZN(n13136) );
  AOI22_X1 U1362 ( .A1(ram[418]), .A2(n4820), .B1(n13150), .B2(n8921), .ZN(
        n4822) );
  INV_X1 U1363 ( .A(n4823), .ZN(n13137) );
  AOI22_X1 U1364 ( .A1(ram[419]), .A2(n4820), .B1(n13150), .B2(n8945), .ZN(
        n4823) );
  INV_X1 U1365 ( .A(n4824), .ZN(n13138) );
  AOI22_X1 U1366 ( .A1(ram[420]), .A2(n4820), .B1(n13150), .B2(n8969), .ZN(
        n4824) );
  INV_X1 U1367 ( .A(n4825), .ZN(n13139) );
  AOI22_X1 U1368 ( .A1(ram[421]), .A2(n4820), .B1(n13150), .B2(n8993), .ZN(
        n4825) );
  INV_X1 U1369 ( .A(n4826), .ZN(n13140) );
  AOI22_X1 U1370 ( .A1(ram[422]), .A2(n4820), .B1(n13150), .B2(n9017), .ZN(
        n4826) );
  INV_X1 U1371 ( .A(n4827), .ZN(n13141) );
  AOI22_X1 U1372 ( .A1(ram[423]), .A2(n4820), .B1(n13150), .B2(n9041), .ZN(
        n4827) );
  INV_X1 U1373 ( .A(n4828), .ZN(n13142) );
  AOI22_X1 U1374 ( .A1(ram[424]), .A2(n4820), .B1(n13150), .B2(n9065), .ZN(
        n4828) );
  INV_X1 U1375 ( .A(n4829), .ZN(n13143) );
  AOI22_X1 U1376 ( .A1(ram[425]), .A2(n4820), .B1(n13150), .B2(n9089), .ZN(
        n4829) );
  INV_X1 U1377 ( .A(n4830), .ZN(n13144) );
  AOI22_X1 U1378 ( .A1(ram[426]), .A2(n4820), .B1(n13150), .B2(n9113), .ZN(
        n4830) );
  INV_X1 U1379 ( .A(n4831), .ZN(n13145) );
  AOI22_X1 U1380 ( .A1(ram[427]), .A2(n4820), .B1(n13150), .B2(n9137), .ZN(
        n4831) );
  INV_X1 U1381 ( .A(n4832), .ZN(n13146) );
  AOI22_X1 U1382 ( .A1(ram[428]), .A2(n4820), .B1(n13150), .B2(n9161), .ZN(
        n4832) );
  INV_X1 U1383 ( .A(n4833), .ZN(n13147) );
  AOI22_X1 U1384 ( .A1(ram[429]), .A2(n4820), .B1(n13150), .B2(n9185), .ZN(
        n4833) );
  INV_X1 U1385 ( .A(n4834), .ZN(n13148) );
  AOI22_X1 U1386 ( .A1(ram[430]), .A2(n4820), .B1(n13150), .B2(n9209), .ZN(
        n4834) );
  INV_X1 U1387 ( .A(n4835), .ZN(n13149) );
  AOI22_X1 U1388 ( .A1(ram[431]), .A2(n4820), .B1(n13150), .B2(n9233), .ZN(
        n4835) );
  INV_X1 U1389 ( .A(n4853), .ZN(n13100) );
  AOI22_X1 U1390 ( .A1(ram[448]), .A2(n4854), .B1(n13116), .B2(n8872), .ZN(
        n4853) );
  INV_X1 U1391 ( .A(n4855), .ZN(n13101) );
  AOI22_X1 U1392 ( .A1(ram[449]), .A2(n4854), .B1(n13116), .B2(n8896), .ZN(
        n4855) );
  INV_X1 U1393 ( .A(n4856), .ZN(n13102) );
  AOI22_X1 U1394 ( .A1(ram[450]), .A2(n4854), .B1(n13116), .B2(n8920), .ZN(
        n4856) );
  INV_X1 U1395 ( .A(n4857), .ZN(n13103) );
  AOI22_X1 U1396 ( .A1(ram[451]), .A2(n4854), .B1(n13116), .B2(n8944), .ZN(
        n4857) );
  INV_X1 U1397 ( .A(n4858), .ZN(n13104) );
  AOI22_X1 U1398 ( .A1(ram[452]), .A2(n4854), .B1(n13116), .B2(n8968), .ZN(
        n4858) );
  INV_X1 U1399 ( .A(n4859), .ZN(n13105) );
  AOI22_X1 U1400 ( .A1(ram[453]), .A2(n4854), .B1(n13116), .B2(n8992), .ZN(
        n4859) );
  INV_X1 U1401 ( .A(n4860), .ZN(n13106) );
  AOI22_X1 U1402 ( .A1(ram[454]), .A2(n4854), .B1(n13116), .B2(n9016), .ZN(
        n4860) );
  INV_X1 U1403 ( .A(n4861), .ZN(n13107) );
  AOI22_X1 U1404 ( .A1(ram[455]), .A2(n4854), .B1(n13116), .B2(n9040), .ZN(
        n4861) );
  INV_X1 U1405 ( .A(n4862), .ZN(n13108) );
  AOI22_X1 U1406 ( .A1(ram[456]), .A2(n4854), .B1(n13116), .B2(n9064), .ZN(
        n4862) );
  INV_X1 U1407 ( .A(n4863), .ZN(n13109) );
  AOI22_X1 U1408 ( .A1(ram[457]), .A2(n4854), .B1(n13116), .B2(n9088), .ZN(
        n4863) );
  INV_X1 U1409 ( .A(n4864), .ZN(n13110) );
  AOI22_X1 U1410 ( .A1(ram[458]), .A2(n4854), .B1(n13116), .B2(n9112), .ZN(
        n4864) );
  INV_X1 U1411 ( .A(n4865), .ZN(n13111) );
  AOI22_X1 U1412 ( .A1(ram[459]), .A2(n4854), .B1(n13116), .B2(n9136), .ZN(
        n4865) );
  INV_X1 U1413 ( .A(n4866), .ZN(n13112) );
  AOI22_X1 U1414 ( .A1(ram[460]), .A2(n4854), .B1(n13116), .B2(n9160), .ZN(
        n4866) );
  INV_X1 U1415 ( .A(n4867), .ZN(n13113) );
  AOI22_X1 U1416 ( .A1(ram[461]), .A2(n4854), .B1(n13116), .B2(n9184), .ZN(
        n4867) );
  INV_X1 U1417 ( .A(n4868), .ZN(n13114) );
  AOI22_X1 U1418 ( .A1(ram[462]), .A2(n4854), .B1(n13116), .B2(n9208), .ZN(
        n4868) );
  INV_X1 U1419 ( .A(n4869), .ZN(n13115) );
  AOI22_X1 U1420 ( .A1(ram[463]), .A2(n4854), .B1(n13116), .B2(n9232), .ZN(
        n4869) );
  INV_X1 U1421 ( .A(n4887), .ZN(n13066) );
  AOI22_X1 U1422 ( .A1(ram[480]), .A2(n4888), .B1(n13082), .B2(n8872), .ZN(
        n4887) );
  INV_X1 U1423 ( .A(n4889), .ZN(n13067) );
  AOI22_X1 U1424 ( .A1(ram[481]), .A2(n4888), .B1(n13082), .B2(n8896), .ZN(
        n4889) );
  INV_X1 U1425 ( .A(n4890), .ZN(n13068) );
  AOI22_X1 U1426 ( .A1(ram[482]), .A2(n4888), .B1(n13082), .B2(n8920), .ZN(
        n4890) );
  INV_X1 U1427 ( .A(n4891), .ZN(n13069) );
  AOI22_X1 U1428 ( .A1(ram[483]), .A2(n4888), .B1(n13082), .B2(n8944), .ZN(
        n4891) );
  INV_X1 U1429 ( .A(n4892), .ZN(n13070) );
  AOI22_X1 U1430 ( .A1(ram[484]), .A2(n4888), .B1(n13082), .B2(n8968), .ZN(
        n4892) );
  INV_X1 U1431 ( .A(n4893), .ZN(n13071) );
  AOI22_X1 U1432 ( .A1(ram[485]), .A2(n4888), .B1(n13082), .B2(n8992), .ZN(
        n4893) );
  INV_X1 U1433 ( .A(n4894), .ZN(n13072) );
  AOI22_X1 U1434 ( .A1(ram[486]), .A2(n4888), .B1(n13082), .B2(n9016), .ZN(
        n4894) );
  INV_X1 U1435 ( .A(n4895), .ZN(n13073) );
  AOI22_X1 U1436 ( .A1(ram[487]), .A2(n4888), .B1(n13082), .B2(n9040), .ZN(
        n4895) );
  INV_X1 U1437 ( .A(n4896), .ZN(n13074) );
  AOI22_X1 U1438 ( .A1(ram[488]), .A2(n4888), .B1(n13082), .B2(n9064), .ZN(
        n4896) );
  INV_X1 U1439 ( .A(n4897), .ZN(n13075) );
  AOI22_X1 U1440 ( .A1(ram[489]), .A2(n4888), .B1(n13082), .B2(n9088), .ZN(
        n4897) );
  INV_X1 U1441 ( .A(n4898), .ZN(n13076) );
  AOI22_X1 U1442 ( .A1(ram[490]), .A2(n4888), .B1(n13082), .B2(n9112), .ZN(
        n4898) );
  INV_X1 U1443 ( .A(n4899), .ZN(n13077) );
  AOI22_X1 U1444 ( .A1(ram[491]), .A2(n4888), .B1(n13082), .B2(n9136), .ZN(
        n4899) );
  INV_X1 U1445 ( .A(n4900), .ZN(n13078) );
  AOI22_X1 U1446 ( .A1(ram[492]), .A2(n4888), .B1(n13082), .B2(n9160), .ZN(
        n4900) );
  INV_X1 U1447 ( .A(n4901), .ZN(n13079) );
  AOI22_X1 U1448 ( .A1(ram[493]), .A2(n4888), .B1(n13082), .B2(n9184), .ZN(
        n4901) );
  INV_X1 U1449 ( .A(n4902), .ZN(n13080) );
  AOI22_X1 U1450 ( .A1(ram[494]), .A2(n4888), .B1(n13082), .B2(n9208), .ZN(
        n4902) );
  INV_X1 U1451 ( .A(n4903), .ZN(n13081) );
  AOI22_X1 U1452 ( .A1(ram[495]), .A2(n4888), .B1(n13082), .B2(n9232), .ZN(
        n4903) );
  INV_X1 U1453 ( .A(n4922), .ZN(n13032) );
  AOI22_X1 U1454 ( .A1(ram[512]), .A2(n4923), .B1(n13048), .B2(n8872), .ZN(
        n4922) );
  INV_X1 U1455 ( .A(n4924), .ZN(n13033) );
  AOI22_X1 U1456 ( .A1(ram[513]), .A2(n4923), .B1(n13048), .B2(n8896), .ZN(
        n4924) );
  INV_X1 U1457 ( .A(n4925), .ZN(n13034) );
  AOI22_X1 U1458 ( .A1(ram[514]), .A2(n4923), .B1(n13048), .B2(n8920), .ZN(
        n4925) );
  INV_X1 U1459 ( .A(n4926), .ZN(n13035) );
  AOI22_X1 U1460 ( .A1(ram[515]), .A2(n4923), .B1(n13048), .B2(n8944), .ZN(
        n4926) );
  INV_X1 U1461 ( .A(n4927), .ZN(n13036) );
  AOI22_X1 U1462 ( .A1(ram[516]), .A2(n4923), .B1(n13048), .B2(n8968), .ZN(
        n4927) );
  INV_X1 U1463 ( .A(n4928), .ZN(n13037) );
  AOI22_X1 U1464 ( .A1(ram[517]), .A2(n4923), .B1(n13048), .B2(n8992), .ZN(
        n4928) );
  INV_X1 U1465 ( .A(n4929), .ZN(n13038) );
  AOI22_X1 U1466 ( .A1(ram[518]), .A2(n4923), .B1(n13048), .B2(n9016), .ZN(
        n4929) );
  INV_X1 U1467 ( .A(n4930), .ZN(n13039) );
  AOI22_X1 U1468 ( .A1(ram[519]), .A2(n4923), .B1(n13048), .B2(n9040), .ZN(
        n4930) );
  INV_X1 U1469 ( .A(n4931), .ZN(n13040) );
  AOI22_X1 U1470 ( .A1(ram[520]), .A2(n4923), .B1(n13048), .B2(n9064), .ZN(
        n4931) );
  INV_X1 U1471 ( .A(n4932), .ZN(n13041) );
  AOI22_X1 U1472 ( .A1(ram[521]), .A2(n4923), .B1(n13048), .B2(n9088), .ZN(
        n4932) );
  INV_X1 U1473 ( .A(n4933), .ZN(n13042) );
  AOI22_X1 U1474 ( .A1(ram[522]), .A2(n4923), .B1(n13048), .B2(n9112), .ZN(
        n4933) );
  INV_X1 U1475 ( .A(n4934), .ZN(n13043) );
  AOI22_X1 U1476 ( .A1(ram[523]), .A2(n4923), .B1(n13048), .B2(n9136), .ZN(
        n4934) );
  INV_X1 U1477 ( .A(n4935), .ZN(n13044) );
  AOI22_X1 U1478 ( .A1(ram[524]), .A2(n4923), .B1(n13048), .B2(n9160), .ZN(
        n4935) );
  INV_X1 U1479 ( .A(n4936), .ZN(n13045) );
  AOI22_X1 U1480 ( .A1(ram[525]), .A2(n4923), .B1(n13048), .B2(n9184), .ZN(
        n4936) );
  INV_X1 U1481 ( .A(n4937), .ZN(n13046) );
  AOI22_X1 U1482 ( .A1(ram[526]), .A2(n4923), .B1(n13048), .B2(n9208), .ZN(
        n4937) );
  INV_X1 U1483 ( .A(n4938), .ZN(n13047) );
  AOI22_X1 U1484 ( .A1(ram[527]), .A2(n4923), .B1(n13048), .B2(n9232), .ZN(
        n4938) );
  INV_X1 U1485 ( .A(n4957), .ZN(n12998) );
  AOI22_X1 U1486 ( .A1(ram[544]), .A2(n4958), .B1(n13014), .B2(n8872), .ZN(
        n4957) );
  INV_X1 U1487 ( .A(n4959), .ZN(n12999) );
  AOI22_X1 U1488 ( .A1(ram[545]), .A2(n4958), .B1(n13014), .B2(n8896), .ZN(
        n4959) );
  INV_X1 U1489 ( .A(n4960), .ZN(n13000) );
  AOI22_X1 U1490 ( .A1(ram[546]), .A2(n4958), .B1(n13014), .B2(n8920), .ZN(
        n4960) );
  INV_X1 U1491 ( .A(n4961), .ZN(n13001) );
  AOI22_X1 U1492 ( .A1(ram[547]), .A2(n4958), .B1(n13014), .B2(n8944), .ZN(
        n4961) );
  INV_X1 U1493 ( .A(n4962), .ZN(n13002) );
  AOI22_X1 U1494 ( .A1(ram[548]), .A2(n4958), .B1(n13014), .B2(n8968), .ZN(
        n4962) );
  INV_X1 U1495 ( .A(n4963), .ZN(n13003) );
  AOI22_X1 U1496 ( .A1(ram[549]), .A2(n4958), .B1(n13014), .B2(n8992), .ZN(
        n4963) );
  INV_X1 U1497 ( .A(n4964), .ZN(n13004) );
  AOI22_X1 U1498 ( .A1(ram[550]), .A2(n4958), .B1(n13014), .B2(n9016), .ZN(
        n4964) );
  INV_X1 U1499 ( .A(n4965), .ZN(n13005) );
  AOI22_X1 U1500 ( .A1(ram[551]), .A2(n4958), .B1(n13014), .B2(n9040), .ZN(
        n4965) );
  INV_X1 U1501 ( .A(n4966), .ZN(n13006) );
  AOI22_X1 U1502 ( .A1(ram[552]), .A2(n4958), .B1(n13014), .B2(n9064), .ZN(
        n4966) );
  INV_X1 U1503 ( .A(n4967), .ZN(n13007) );
  AOI22_X1 U1504 ( .A1(ram[553]), .A2(n4958), .B1(n13014), .B2(n9088), .ZN(
        n4967) );
  INV_X1 U1505 ( .A(n4968), .ZN(n13008) );
  AOI22_X1 U1506 ( .A1(ram[554]), .A2(n4958), .B1(n13014), .B2(n9112), .ZN(
        n4968) );
  INV_X1 U1507 ( .A(n4969), .ZN(n13009) );
  AOI22_X1 U1508 ( .A1(ram[555]), .A2(n4958), .B1(n13014), .B2(n9136), .ZN(
        n4969) );
  INV_X1 U1509 ( .A(n4970), .ZN(n13010) );
  AOI22_X1 U1510 ( .A1(ram[556]), .A2(n4958), .B1(n13014), .B2(n9160), .ZN(
        n4970) );
  INV_X1 U1511 ( .A(n4971), .ZN(n13011) );
  AOI22_X1 U1512 ( .A1(ram[557]), .A2(n4958), .B1(n13014), .B2(n9184), .ZN(
        n4971) );
  INV_X1 U1513 ( .A(n4972), .ZN(n13012) );
  AOI22_X1 U1514 ( .A1(ram[558]), .A2(n4958), .B1(n13014), .B2(n9208), .ZN(
        n4972) );
  INV_X1 U1515 ( .A(n4973), .ZN(n13013) );
  AOI22_X1 U1516 ( .A1(ram[559]), .A2(n4958), .B1(n13014), .B2(n9232), .ZN(
        n4973) );
  INV_X1 U1517 ( .A(n4991), .ZN(n12964) );
  AOI22_X1 U1518 ( .A1(ram[576]), .A2(n4992), .B1(n12980), .B2(n8872), .ZN(
        n4991) );
  INV_X1 U1519 ( .A(n4993), .ZN(n12965) );
  AOI22_X1 U1520 ( .A1(ram[577]), .A2(n4992), .B1(n12980), .B2(n8896), .ZN(
        n4993) );
  INV_X1 U1521 ( .A(n4994), .ZN(n12966) );
  AOI22_X1 U1522 ( .A1(ram[578]), .A2(n4992), .B1(n12980), .B2(n8920), .ZN(
        n4994) );
  INV_X1 U1523 ( .A(n4995), .ZN(n12967) );
  AOI22_X1 U1524 ( .A1(ram[579]), .A2(n4992), .B1(n12980), .B2(n8944), .ZN(
        n4995) );
  INV_X1 U1525 ( .A(n4996), .ZN(n12968) );
  AOI22_X1 U1526 ( .A1(ram[580]), .A2(n4992), .B1(n12980), .B2(n8968), .ZN(
        n4996) );
  INV_X1 U1527 ( .A(n4997), .ZN(n12969) );
  AOI22_X1 U1528 ( .A1(ram[581]), .A2(n4992), .B1(n12980), .B2(n8992), .ZN(
        n4997) );
  INV_X1 U1529 ( .A(n4998), .ZN(n12970) );
  AOI22_X1 U1530 ( .A1(ram[582]), .A2(n4992), .B1(n12980), .B2(n9016), .ZN(
        n4998) );
  INV_X1 U1531 ( .A(n4999), .ZN(n12971) );
  AOI22_X1 U1532 ( .A1(ram[583]), .A2(n4992), .B1(n12980), .B2(n9040), .ZN(
        n4999) );
  INV_X1 U1533 ( .A(n5000), .ZN(n12972) );
  AOI22_X1 U1534 ( .A1(ram[584]), .A2(n4992), .B1(n12980), .B2(n9064), .ZN(
        n5000) );
  INV_X1 U1535 ( .A(n5001), .ZN(n12973) );
  AOI22_X1 U1536 ( .A1(ram[585]), .A2(n4992), .B1(n12980), .B2(n9088), .ZN(
        n5001) );
  INV_X1 U1537 ( .A(n5002), .ZN(n12974) );
  AOI22_X1 U1538 ( .A1(ram[586]), .A2(n4992), .B1(n12980), .B2(n9112), .ZN(
        n5002) );
  INV_X1 U1539 ( .A(n5003), .ZN(n12975) );
  AOI22_X1 U1540 ( .A1(ram[587]), .A2(n4992), .B1(n12980), .B2(n9136), .ZN(
        n5003) );
  INV_X1 U1541 ( .A(n5004), .ZN(n12976) );
  AOI22_X1 U1542 ( .A1(ram[588]), .A2(n4992), .B1(n12980), .B2(n9160), .ZN(
        n5004) );
  INV_X1 U1543 ( .A(n5005), .ZN(n12977) );
  AOI22_X1 U1544 ( .A1(ram[589]), .A2(n4992), .B1(n12980), .B2(n9184), .ZN(
        n5005) );
  INV_X1 U1545 ( .A(n5006), .ZN(n12978) );
  AOI22_X1 U1546 ( .A1(ram[590]), .A2(n4992), .B1(n12980), .B2(n9208), .ZN(
        n5006) );
  INV_X1 U1547 ( .A(n5007), .ZN(n12979) );
  AOI22_X1 U1548 ( .A1(ram[591]), .A2(n4992), .B1(n12980), .B2(n9232), .ZN(
        n5007) );
  INV_X1 U1549 ( .A(n5025), .ZN(n12930) );
  AOI22_X1 U1550 ( .A1(ram[608]), .A2(n5026), .B1(n12946), .B2(n8872), .ZN(
        n5025) );
  INV_X1 U1551 ( .A(n5027), .ZN(n12931) );
  AOI22_X1 U1552 ( .A1(ram[609]), .A2(n5026), .B1(n12946), .B2(n8896), .ZN(
        n5027) );
  INV_X1 U1553 ( .A(n5028), .ZN(n12932) );
  AOI22_X1 U1554 ( .A1(ram[610]), .A2(n5026), .B1(n12946), .B2(n8920), .ZN(
        n5028) );
  INV_X1 U1555 ( .A(n5029), .ZN(n12933) );
  AOI22_X1 U1556 ( .A1(ram[611]), .A2(n5026), .B1(n12946), .B2(n8944), .ZN(
        n5029) );
  INV_X1 U1557 ( .A(n5030), .ZN(n12934) );
  AOI22_X1 U1558 ( .A1(ram[612]), .A2(n5026), .B1(n12946), .B2(n8968), .ZN(
        n5030) );
  INV_X1 U1559 ( .A(n5031), .ZN(n12935) );
  AOI22_X1 U1560 ( .A1(ram[613]), .A2(n5026), .B1(n12946), .B2(n8992), .ZN(
        n5031) );
  INV_X1 U1561 ( .A(n5032), .ZN(n12936) );
  AOI22_X1 U1562 ( .A1(ram[614]), .A2(n5026), .B1(n12946), .B2(n9016), .ZN(
        n5032) );
  INV_X1 U1563 ( .A(n5033), .ZN(n12937) );
  AOI22_X1 U1564 ( .A1(ram[615]), .A2(n5026), .B1(n12946), .B2(n9040), .ZN(
        n5033) );
  INV_X1 U1565 ( .A(n5034), .ZN(n12938) );
  AOI22_X1 U1566 ( .A1(ram[616]), .A2(n5026), .B1(n12946), .B2(n9064), .ZN(
        n5034) );
  INV_X1 U1567 ( .A(n5035), .ZN(n12939) );
  AOI22_X1 U1568 ( .A1(ram[617]), .A2(n5026), .B1(n12946), .B2(n9088), .ZN(
        n5035) );
  INV_X1 U1569 ( .A(n5036), .ZN(n12940) );
  AOI22_X1 U1570 ( .A1(ram[618]), .A2(n5026), .B1(n12946), .B2(n9112), .ZN(
        n5036) );
  INV_X1 U1571 ( .A(n5037), .ZN(n12941) );
  AOI22_X1 U1572 ( .A1(ram[619]), .A2(n5026), .B1(n12946), .B2(n9136), .ZN(
        n5037) );
  INV_X1 U1573 ( .A(n5038), .ZN(n12942) );
  AOI22_X1 U1574 ( .A1(ram[620]), .A2(n5026), .B1(n12946), .B2(n9160), .ZN(
        n5038) );
  INV_X1 U1575 ( .A(n5039), .ZN(n12943) );
  AOI22_X1 U1576 ( .A1(ram[621]), .A2(n5026), .B1(n12946), .B2(n9184), .ZN(
        n5039) );
  INV_X1 U1577 ( .A(n5040), .ZN(n12944) );
  AOI22_X1 U1578 ( .A1(ram[622]), .A2(n5026), .B1(n12946), .B2(n9208), .ZN(
        n5040) );
  INV_X1 U1579 ( .A(n5041), .ZN(n12945) );
  AOI22_X1 U1580 ( .A1(ram[623]), .A2(n5026), .B1(n12946), .B2(n9232), .ZN(
        n5041) );
  INV_X1 U1581 ( .A(n5059), .ZN(n12896) );
  AOI22_X1 U1582 ( .A1(ram[640]), .A2(n5060), .B1(n12912), .B2(n8871), .ZN(
        n5059) );
  INV_X1 U1583 ( .A(n5061), .ZN(n12897) );
  AOI22_X1 U1584 ( .A1(ram[641]), .A2(n5060), .B1(n12912), .B2(n8895), .ZN(
        n5061) );
  INV_X1 U1585 ( .A(n5062), .ZN(n12898) );
  AOI22_X1 U1586 ( .A1(ram[642]), .A2(n5060), .B1(n12912), .B2(n8919), .ZN(
        n5062) );
  INV_X1 U1587 ( .A(n5063), .ZN(n12899) );
  AOI22_X1 U1588 ( .A1(ram[643]), .A2(n5060), .B1(n12912), .B2(n8943), .ZN(
        n5063) );
  INV_X1 U1589 ( .A(n5064), .ZN(n12900) );
  AOI22_X1 U1590 ( .A1(ram[644]), .A2(n5060), .B1(n12912), .B2(n8967), .ZN(
        n5064) );
  INV_X1 U1591 ( .A(n5065), .ZN(n12901) );
  AOI22_X1 U1592 ( .A1(ram[645]), .A2(n5060), .B1(n12912), .B2(n8991), .ZN(
        n5065) );
  INV_X1 U1593 ( .A(n5066), .ZN(n12902) );
  AOI22_X1 U1594 ( .A1(ram[646]), .A2(n5060), .B1(n12912), .B2(n9015), .ZN(
        n5066) );
  INV_X1 U1595 ( .A(n5067), .ZN(n12903) );
  AOI22_X1 U1596 ( .A1(ram[647]), .A2(n5060), .B1(n12912), .B2(n9039), .ZN(
        n5067) );
  INV_X1 U1597 ( .A(n5068), .ZN(n12904) );
  AOI22_X1 U1598 ( .A1(ram[648]), .A2(n5060), .B1(n12912), .B2(n9063), .ZN(
        n5068) );
  INV_X1 U1599 ( .A(n5069), .ZN(n12905) );
  AOI22_X1 U1600 ( .A1(ram[649]), .A2(n5060), .B1(n12912), .B2(n9087), .ZN(
        n5069) );
  INV_X1 U1601 ( .A(n5070), .ZN(n12906) );
  AOI22_X1 U1602 ( .A1(ram[650]), .A2(n5060), .B1(n12912), .B2(n9111), .ZN(
        n5070) );
  INV_X1 U1603 ( .A(n5071), .ZN(n12907) );
  AOI22_X1 U1604 ( .A1(ram[651]), .A2(n5060), .B1(n12912), .B2(n9135), .ZN(
        n5071) );
  INV_X1 U1605 ( .A(n5072), .ZN(n12908) );
  AOI22_X1 U1606 ( .A1(ram[652]), .A2(n5060), .B1(n12912), .B2(n9159), .ZN(
        n5072) );
  INV_X1 U1607 ( .A(n5073), .ZN(n12909) );
  AOI22_X1 U1608 ( .A1(ram[653]), .A2(n5060), .B1(n12912), .B2(n9183), .ZN(
        n5073) );
  INV_X1 U1609 ( .A(n5074), .ZN(n12910) );
  AOI22_X1 U1610 ( .A1(ram[654]), .A2(n5060), .B1(n12912), .B2(n9207), .ZN(
        n5074) );
  INV_X1 U1611 ( .A(n5075), .ZN(n12911) );
  AOI22_X1 U1612 ( .A1(ram[655]), .A2(n5060), .B1(n12912), .B2(n9231), .ZN(
        n5075) );
  INV_X1 U1613 ( .A(n5093), .ZN(n12862) );
  AOI22_X1 U1614 ( .A1(ram[672]), .A2(n5094), .B1(n12878), .B2(n8871), .ZN(
        n5093) );
  INV_X1 U1615 ( .A(n5095), .ZN(n12863) );
  AOI22_X1 U1616 ( .A1(ram[673]), .A2(n5094), .B1(n12878), .B2(n8895), .ZN(
        n5095) );
  INV_X1 U1617 ( .A(n5096), .ZN(n12864) );
  AOI22_X1 U1618 ( .A1(ram[674]), .A2(n5094), .B1(n12878), .B2(n8919), .ZN(
        n5096) );
  INV_X1 U1619 ( .A(n5097), .ZN(n12865) );
  AOI22_X1 U1620 ( .A1(ram[675]), .A2(n5094), .B1(n12878), .B2(n8943), .ZN(
        n5097) );
  INV_X1 U1621 ( .A(n5098), .ZN(n12866) );
  AOI22_X1 U1622 ( .A1(ram[676]), .A2(n5094), .B1(n12878), .B2(n8967), .ZN(
        n5098) );
  INV_X1 U1623 ( .A(n5099), .ZN(n12867) );
  AOI22_X1 U1624 ( .A1(ram[677]), .A2(n5094), .B1(n12878), .B2(n8991), .ZN(
        n5099) );
  INV_X1 U1625 ( .A(n5100), .ZN(n12868) );
  AOI22_X1 U1626 ( .A1(ram[678]), .A2(n5094), .B1(n12878), .B2(n9015), .ZN(
        n5100) );
  INV_X1 U1627 ( .A(n5101), .ZN(n12869) );
  AOI22_X1 U1628 ( .A1(ram[679]), .A2(n5094), .B1(n12878), .B2(n9039), .ZN(
        n5101) );
  INV_X1 U1629 ( .A(n5102), .ZN(n12870) );
  AOI22_X1 U1630 ( .A1(ram[680]), .A2(n5094), .B1(n12878), .B2(n9063), .ZN(
        n5102) );
  INV_X1 U1631 ( .A(n5103), .ZN(n12871) );
  AOI22_X1 U1632 ( .A1(ram[681]), .A2(n5094), .B1(n12878), .B2(n9087), .ZN(
        n5103) );
  INV_X1 U1633 ( .A(n5104), .ZN(n12872) );
  AOI22_X1 U1634 ( .A1(ram[682]), .A2(n5094), .B1(n12878), .B2(n9111), .ZN(
        n5104) );
  INV_X1 U1635 ( .A(n5105), .ZN(n12873) );
  AOI22_X1 U1636 ( .A1(ram[683]), .A2(n5094), .B1(n12878), .B2(n9135), .ZN(
        n5105) );
  INV_X1 U1637 ( .A(n5106), .ZN(n12874) );
  AOI22_X1 U1638 ( .A1(ram[684]), .A2(n5094), .B1(n12878), .B2(n9159), .ZN(
        n5106) );
  INV_X1 U1639 ( .A(n5107), .ZN(n12875) );
  AOI22_X1 U1640 ( .A1(ram[685]), .A2(n5094), .B1(n12878), .B2(n9183), .ZN(
        n5107) );
  INV_X1 U1641 ( .A(n5108), .ZN(n12876) );
  AOI22_X1 U1642 ( .A1(ram[686]), .A2(n5094), .B1(n12878), .B2(n9207), .ZN(
        n5108) );
  INV_X1 U1643 ( .A(n5109), .ZN(n12877) );
  AOI22_X1 U1644 ( .A1(ram[687]), .A2(n5094), .B1(n12878), .B2(n9231), .ZN(
        n5109) );
  INV_X1 U1645 ( .A(n5127), .ZN(n12828) );
  AOI22_X1 U1646 ( .A1(ram[704]), .A2(n5128), .B1(n12844), .B2(n8871), .ZN(
        n5127) );
  INV_X1 U1647 ( .A(n5129), .ZN(n12829) );
  AOI22_X1 U1648 ( .A1(ram[705]), .A2(n5128), .B1(n12844), .B2(n8895), .ZN(
        n5129) );
  INV_X1 U1649 ( .A(n5130), .ZN(n12830) );
  AOI22_X1 U1650 ( .A1(ram[706]), .A2(n5128), .B1(n12844), .B2(n8919), .ZN(
        n5130) );
  INV_X1 U1651 ( .A(n5131), .ZN(n12831) );
  AOI22_X1 U1652 ( .A1(ram[707]), .A2(n5128), .B1(n12844), .B2(n8943), .ZN(
        n5131) );
  INV_X1 U1653 ( .A(n5132), .ZN(n12832) );
  AOI22_X1 U1654 ( .A1(ram[708]), .A2(n5128), .B1(n12844), .B2(n8967), .ZN(
        n5132) );
  INV_X1 U1655 ( .A(n5133), .ZN(n12833) );
  AOI22_X1 U1656 ( .A1(ram[709]), .A2(n5128), .B1(n12844), .B2(n8991), .ZN(
        n5133) );
  INV_X1 U1657 ( .A(n5134), .ZN(n12834) );
  AOI22_X1 U1658 ( .A1(ram[710]), .A2(n5128), .B1(n12844), .B2(n9015), .ZN(
        n5134) );
  INV_X1 U1659 ( .A(n5135), .ZN(n12835) );
  AOI22_X1 U1660 ( .A1(ram[711]), .A2(n5128), .B1(n12844), .B2(n9039), .ZN(
        n5135) );
  INV_X1 U1661 ( .A(n5136), .ZN(n12836) );
  AOI22_X1 U1662 ( .A1(ram[712]), .A2(n5128), .B1(n12844), .B2(n9063), .ZN(
        n5136) );
  INV_X1 U1663 ( .A(n5137), .ZN(n12837) );
  AOI22_X1 U1664 ( .A1(ram[713]), .A2(n5128), .B1(n12844), .B2(n9087), .ZN(
        n5137) );
  INV_X1 U1665 ( .A(n5138), .ZN(n12838) );
  AOI22_X1 U1666 ( .A1(ram[714]), .A2(n5128), .B1(n12844), .B2(n9111), .ZN(
        n5138) );
  INV_X1 U1667 ( .A(n5139), .ZN(n12839) );
  AOI22_X1 U1668 ( .A1(ram[715]), .A2(n5128), .B1(n12844), .B2(n9135), .ZN(
        n5139) );
  INV_X1 U1669 ( .A(n5140), .ZN(n12840) );
  AOI22_X1 U1670 ( .A1(ram[716]), .A2(n5128), .B1(n12844), .B2(n9159), .ZN(
        n5140) );
  INV_X1 U1671 ( .A(n5141), .ZN(n12841) );
  AOI22_X1 U1672 ( .A1(ram[717]), .A2(n5128), .B1(n12844), .B2(n9183), .ZN(
        n5141) );
  INV_X1 U1673 ( .A(n5142), .ZN(n12842) );
  AOI22_X1 U1674 ( .A1(ram[718]), .A2(n5128), .B1(n12844), .B2(n9207), .ZN(
        n5142) );
  INV_X1 U1675 ( .A(n5143), .ZN(n12843) );
  AOI22_X1 U1676 ( .A1(ram[719]), .A2(n5128), .B1(n12844), .B2(n9231), .ZN(
        n5143) );
  INV_X1 U1677 ( .A(n5161), .ZN(n12794) );
  AOI22_X1 U1678 ( .A1(ram[736]), .A2(n5162), .B1(n12810), .B2(n8871), .ZN(
        n5161) );
  INV_X1 U1679 ( .A(n5163), .ZN(n12795) );
  AOI22_X1 U1680 ( .A1(ram[737]), .A2(n5162), .B1(n12810), .B2(n8895), .ZN(
        n5163) );
  INV_X1 U1681 ( .A(n5164), .ZN(n12796) );
  AOI22_X1 U1682 ( .A1(ram[738]), .A2(n5162), .B1(n12810), .B2(n8919), .ZN(
        n5164) );
  INV_X1 U1683 ( .A(n5165), .ZN(n12797) );
  AOI22_X1 U1684 ( .A1(ram[739]), .A2(n5162), .B1(n12810), .B2(n8943), .ZN(
        n5165) );
  INV_X1 U1685 ( .A(n5166), .ZN(n12798) );
  AOI22_X1 U1686 ( .A1(ram[740]), .A2(n5162), .B1(n12810), .B2(n8967), .ZN(
        n5166) );
  INV_X1 U1687 ( .A(n5167), .ZN(n12799) );
  AOI22_X1 U1688 ( .A1(ram[741]), .A2(n5162), .B1(n12810), .B2(n8991), .ZN(
        n5167) );
  INV_X1 U1689 ( .A(n5168), .ZN(n12800) );
  AOI22_X1 U1690 ( .A1(ram[742]), .A2(n5162), .B1(n12810), .B2(n9015), .ZN(
        n5168) );
  INV_X1 U1691 ( .A(n5169), .ZN(n12801) );
  AOI22_X1 U1692 ( .A1(ram[743]), .A2(n5162), .B1(n12810), .B2(n9039), .ZN(
        n5169) );
  INV_X1 U1693 ( .A(n5170), .ZN(n12802) );
  AOI22_X1 U1694 ( .A1(ram[744]), .A2(n5162), .B1(n12810), .B2(n9063), .ZN(
        n5170) );
  INV_X1 U1695 ( .A(n5171), .ZN(n12803) );
  AOI22_X1 U1696 ( .A1(ram[745]), .A2(n5162), .B1(n12810), .B2(n9087), .ZN(
        n5171) );
  INV_X1 U1697 ( .A(n5172), .ZN(n12804) );
  AOI22_X1 U1698 ( .A1(ram[746]), .A2(n5162), .B1(n12810), .B2(n9111), .ZN(
        n5172) );
  INV_X1 U1699 ( .A(n5173), .ZN(n12805) );
  AOI22_X1 U1700 ( .A1(ram[747]), .A2(n5162), .B1(n12810), .B2(n9135), .ZN(
        n5173) );
  INV_X1 U1701 ( .A(n5174), .ZN(n12806) );
  AOI22_X1 U1702 ( .A1(ram[748]), .A2(n5162), .B1(n12810), .B2(n9159), .ZN(
        n5174) );
  INV_X1 U1703 ( .A(n5175), .ZN(n12807) );
  AOI22_X1 U1704 ( .A1(ram[749]), .A2(n5162), .B1(n12810), .B2(n9183), .ZN(
        n5175) );
  INV_X1 U1705 ( .A(n5176), .ZN(n12808) );
  AOI22_X1 U1706 ( .A1(ram[750]), .A2(n5162), .B1(n12810), .B2(n9207), .ZN(
        n5176) );
  INV_X1 U1707 ( .A(n5177), .ZN(n12809) );
  AOI22_X1 U1708 ( .A1(ram[751]), .A2(n5162), .B1(n12810), .B2(n9231), .ZN(
        n5177) );
  INV_X1 U1709 ( .A(n5196), .ZN(n12760) );
  AOI22_X1 U1710 ( .A1(ram[768]), .A2(n5197), .B1(n12776), .B2(n8871), .ZN(
        n5196) );
  INV_X1 U1711 ( .A(n5198), .ZN(n12761) );
  AOI22_X1 U1712 ( .A1(ram[769]), .A2(n5197), .B1(n12776), .B2(n8895), .ZN(
        n5198) );
  INV_X1 U1713 ( .A(n5199), .ZN(n12762) );
  AOI22_X1 U1714 ( .A1(ram[770]), .A2(n5197), .B1(n12776), .B2(n8919), .ZN(
        n5199) );
  INV_X1 U1715 ( .A(n5200), .ZN(n12763) );
  AOI22_X1 U1716 ( .A1(ram[771]), .A2(n5197), .B1(n12776), .B2(n8943), .ZN(
        n5200) );
  INV_X1 U1717 ( .A(n5201), .ZN(n12764) );
  AOI22_X1 U1718 ( .A1(ram[772]), .A2(n5197), .B1(n12776), .B2(n8967), .ZN(
        n5201) );
  INV_X1 U1719 ( .A(n5202), .ZN(n12765) );
  AOI22_X1 U1720 ( .A1(ram[773]), .A2(n5197), .B1(n12776), .B2(n8991), .ZN(
        n5202) );
  INV_X1 U1721 ( .A(n5203), .ZN(n12766) );
  AOI22_X1 U1722 ( .A1(ram[774]), .A2(n5197), .B1(n12776), .B2(n9015), .ZN(
        n5203) );
  INV_X1 U1723 ( .A(n5204), .ZN(n12767) );
  AOI22_X1 U1724 ( .A1(ram[775]), .A2(n5197), .B1(n12776), .B2(n9039), .ZN(
        n5204) );
  INV_X1 U1725 ( .A(n5205), .ZN(n12768) );
  AOI22_X1 U1726 ( .A1(ram[776]), .A2(n5197), .B1(n12776), .B2(n9063), .ZN(
        n5205) );
  INV_X1 U1727 ( .A(n5206), .ZN(n12769) );
  AOI22_X1 U1728 ( .A1(ram[777]), .A2(n5197), .B1(n12776), .B2(n9087), .ZN(
        n5206) );
  INV_X1 U1729 ( .A(n5207), .ZN(n12770) );
  AOI22_X1 U1730 ( .A1(ram[778]), .A2(n5197), .B1(n12776), .B2(n9111), .ZN(
        n5207) );
  INV_X1 U1731 ( .A(n5208), .ZN(n12771) );
  AOI22_X1 U1732 ( .A1(ram[779]), .A2(n5197), .B1(n12776), .B2(n9135), .ZN(
        n5208) );
  INV_X1 U1733 ( .A(n5209), .ZN(n12772) );
  AOI22_X1 U1734 ( .A1(ram[780]), .A2(n5197), .B1(n12776), .B2(n9159), .ZN(
        n5209) );
  INV_X1 U1735 ( .A(n5210), .ZN(n12773) );
  AOI22_X1 U1736 ( .A1(ram[781]), .A2(n5197), .B1(n12776), .B2(n9183), .ZN(
        n5210) );
  INV_X1 U1737 ( .A(n5211), .ZN(n12774) );
  AOI22_X1 U1738 ( .A1(ram[782]), .A2(n5197), .B1(n12776), .B2(n9207), .ZN(
        n5211) );
  INV_X1 U1739 ( .A(n5212), .ZN(n12775) );
  AOI22_X1 U1740 ( .A1(ram[783]), .A2(n5197), .B1(n12776), .B2(n9231), .ZN(
        n5212) );
  INV_X1 U1741 ( .A(n5231), .ZN(n12726) );
  AOI22_X1 U1742 ( .A1(ram[800]), .A2(n5232), .B1(n12742), .B2(n8871), .ZN(
        n5231) );
  INV_X1 U1743 ( .A(n5233), .ZN(n12727) );
  AOI22_X1 U1744 ( .A1(ram[801]), .A2(n5232), .B1(n12742), .B2(n8895), .ZN(
        n5233) );
  INV_X1 U1745 ( .A(n5234), .ZN(n12728) );
  AOI22_X1 U1746 ( .A1(ram[802]), .A2(n5232), .B1(n12742), .B2(n8919), .ZN(
        n5234) );
  INV_X1 U1747 ( .A(n5235), .ZN(n12729) );
  AOI22_X1 U1748 ( .A1(ram[803]), .A2(n5232), .B1(n12742), .B2(n8943), .ZN(
        n5235) );
  INV_X1 U1749 ( .A(n5236), .ZN(n12730) );
  AOI22_X1 U1750 ( .A1(ram[804]), .A2(n5232), .B1(n12742), .B2(n8967), .ZN(
        n5236) );
  INV_X1 U1751 ( .A(n5237), .ZN(n12731) );
  AOI22_X1 U1752 ( .A1(ram[805]), .A2(n5232), .B1(n12742), .B2(n8991), .ZN(
        n5237) );
  INV_X1 U1753 ( .A(n5238), .ZN(n12732) );
  AOI22_X1 U1754 ( .A1(ram[806]), .A2(n5232), .B1(n12742), .B2(n9015), .ZN(
        n5238) );
  INV_X1 U1755 ( .A(n5239), .ZN(n12733) );
  AOI22_X1 U1756 ( .A1(ram[807]), .A2(n5232), .B1(n12742), .B2(n9039), .ZN(
        n5239) );
  INV_X1 U1757 ( .A(n5240), .ZN(n12734) );
  AOI22_X1 U1758 ( .A1(ram[808]), .A2(n5232), .B1(n12742), .B2(n9063), .ZN(
        n5240) );
  INV_X1 U1759 ( .A(n5241), .ZN(n12735) );
  AOI22_X1 U1760 ( .A1(ram[809]), .A2(n5232), .B1(n12742), .B2(n9087), .ZN(
        n5241) );
  INV_X1 U1761 ( .A(n5242), .ZN(n12736) );
  AOI22_X1 U1762 ( .A1(ram[810]), .A2(n5232), .B1(n12742), .B2(n9111), .ZN(
        n5242) );
  INV_X1 U1763 ( .A(n5243), .ZN(n12737) );
  AOI22_X1 U1764 ( .A1(ram[811]), .A2(n5232), .B1(n12742), .B2(n9135), .ZN(
        n5243) );
  INV_X1 U1765 ( .A(n5244), .ZN(n12738) );
  AOI22_X1 U1766 ( .A1(ram[812]), .A2(n5232), .B1(n12742), .B2(n9159), .ZN(
        n5244) );
  INV_X1 U1767 ( .A(n5245), .ZN(n12739) );
  AOI22_X1 U1768 ( .A1(ram[813]), .A2(n5232), .B1(n12742), .B2(n9183), .ZN(
        n5245) );
  INV_X1 U1769 ( .A(n5246), .ZN(n12740) );
  AOI22_X1 U1770 ( .A1(ram[814]), .A2(n5232), .B1(n12742), .B2(n9207), .ZN(
        n5246) );
  INV_X1 U1771 ( .A(n5247), .ZN(n12741) );
  AOI22_X1 U1772 ( .A1(ram[815]), .A2(n5232), .B1(n12742), .B2(n9231), .ZN(
        n5247) );
  INV_X1 U1773 ( .A(n5265), .ZN(n12692) );
  AOI22_X1 U1774 ( .A1(ram[832]), .A2(n5266), .B1(n12708), .B2(n8870), .ZN(
        n5265) );
  INV_X1 U1775 ( .A(n5267), .ZN(n12693) );
  AOI22_X1 U1776 ( .A1(ram[833]), .A2(n5266), .B1(n12708), .B2(n8894), .ZN(
        n5267) );
  INV_X1 U1777 ( .A(n5268), .ZN(n12694) );
  AOI22_X1 U1778 ( .A1(ram[834]), .A2(n5266), .B1(n12708), .B2(n8918), .ZN(
        n5268) );
  INV_X1 U1779 ( .A(n5269), .ZN(n12695) );
  AOI22_X1 U1780 ( .A1(ram[835]), .A2(n5266), .B1(n12708), .B2(n8942), .ZN(
        n5269) );
  INV_X1 U1781 ( .A(n5270), .ZN(n12696) );
  AOI22_X1 U1782 ( .A1(ram[836]), .A2(n5266), .B1(n12708), .B2(n8966), .ZN(
        n5270) );
  INV_X1 U1783 ( .A(n5271), .ZN(n12697) );
  AOI22_X1 U1784 ( .A1(ram[837]), .A2(n5266), .B1(n12708), .B2(n8990), .ZN(
        n5271) );
  INV_X1 U1785 ( .A(n5272), .ZN(n12698) );
  AOI22_X1 U1786 ( .A1(ram[838]), .A2(n5266), .B1(n12708), .B2(n9014), .ZN(
        n5272) );
  INV_X1 U1787 ( .A(n5273), .ZN(n12699) );
  AOI22_X1 U1788 ( .A1(ram[839]), .A2(n5266), .B1(n12708), .B2(n9038), .ZN(
        n5273) );
  INV_X1 U1789 ( .A(n5274), .ZN(n12700) );
  AOI22_X1 U1790 ( .A1(ram[840]), .A2(n5266), .B1(n12708), .B2(n9062), .ZN(
        n5274) );
  INV_X1 U1791 ( .A(n5275), .ZN(n12701) );
  AOI22_X1 U1792 ( .A1(ram[841]), .A2(n5266), .B1(n12708), .B2(n9086), .ZN(
        n5275) );
  INV_X1 U1793 ( .A(n5276), .ZN(n12702) );
  AOI22_X1 U1794 ( .A1(ram[842]), .A2(n5266), .B1(n12708), .B2(n9110), .ZN(
        n5276) );
  INV_X1 U1795 ( .A(n5277), .ZN(n12703) );
  AOI22_X1 U1796 ( .A1(ram[843]), .A2(n5266), .B1(n12708), .B2(n9134), .ZN(
        n5277) );
  INV_X1 U1797 ( .A(n5278), .ZN(n12704) );
  AOI22_X1 U1798 ( .A1(ram[844]), .A2(n5266), .B1(n12708), .B2(n9158), .ZN(
        n5278) );
  INV_X1 U1799 ( .A(n5279), .ZN(n12705) );
  AOI22_X1 U1800 ( .A1(ram[845]), .A2(n5266), .B1(n12708), .B2(n9182), .ZN(
        n5279) );
  INV_X1 U1801 ( .A(n5280), .ZN(n12706) );
  AOI22_X1 U1802 ( .A1(ram[846]), .A2(n5266), .B1(n12708), .B2(n9206), .ZN(
        n5280) );
  INV_X1 U1803 ( .A(n5281), .ZN(n12707) );
  AOI22_X1 U1804 ( .A1(ram[847]), .A2(n5266), .B1(n12708), .B2(n9230), .ZN(
        n5281) );
  INV_X1 U1805 ( .A(n5299), .ZN(n12658) );
  AOI22_X1 U1806 ( .A1(ram[864]), .A2(n5300), .B1(n12674), .B2(n8870), .ZN(
        n5299) );
  INV_X1 U1807 ( .A(n5301), .ZN(n12659) );
  AOI22_X1 U1808 ( .A1(ram[865]), .A2(n5300), .B1(n12674), .B2(n8894), .ZN(
        n5301) );
  INV_X1 U1809 ( .A(n5302), .ZN(n12660) );
  AOI22_X1 U1810 ( .A1(ram[866]), .A2(n5300), .B1(n12674), .B2(n8918), .ZN(
        n5302) );
  INV_X1 U1811 ( .A(n5303), .ZN(n12661) );
  AOI22_X1 U1812 ( .A1(ram[867]), .A2(n5300), .B1(n12674), .B2(n8942), .ZN(
        n5303) );
  INV_X1 U1813 ( .A(n5304), .ZN(n12662) );
  AOI22_X1 U1814 ( .A1(ram[868]), .A2(n5300), .B1(n12674), .B2(n8966), .ZN(
        n5304) );
  INV_X1 U1815 ( .A(n5305), .ZN(n12663) );
  AOI22_X1 U1816 ( .A1(ram[869]), .A2(n5300), .B1(n12674), .B2(n8990), .ZN(
        n5305) );
  INV_X1 U1817 ( .A(n5306), .ZN(n12664) );
  AOI22_X1 U1818 ( .A1(ram[870]), .A2(n5300), .B1(n12674), .B2(n9014), .ZN(
        n5306) );
  INV_X1 U1819 ( .A(n5307), .ZN(n12665) );
  AOI22_X1 U1820 ( .A1(ram[871]), .A2(n5300), .B1(n12674), .B2(n9038), .ZN(
        n5307) );
  INV_X1 U1821 ( .A(n5308), .ZN(n12666) );
  AOI22_X1 U1822 ( .A1(ram[872]), .A2(n5300), .B1(n12674), .B2(n9062), .ZN(
        n5308) );
  INV_X1 U1823 ( .A(n5309), .ZN(n12667) );
  AOI22_X1 U1824 ( .A1(ram[873]), .A2(n5300), .B1(n12674), .B2(n9086), .ZN(
        n5309) );
  INV_X1 U1825 ( .A(n5310), .ZN(n12668) );
  AOI22_X1 U1826 ( .A1(ram[874]), .A2(n5300), .B1(n12674), .B2(n9110), .ZN(
        n5310) );
  INV_X1 U1827 ( .A(n5311), .ZN(n12669) );
  AOI22_X1 U1828 ( .A1(ram[875]), .A2(n5300), .B1(n12674), .B2(n9134), .ZN(
        n5311) );
  INV_X1 U1829 ( .A(n5312), .ZN(n12670) );
  AOI22_X1 U1830 ( .A1(ram[876]), .A2(n5300), .B1(n12674), .B2(n9158), .ZN(
        n5312) );
  INV_X1 U1831 ( .A(n5313), .ZN(n12671) );
  AOI22_X1 U1832 ( .A1(ram[877]), .A2(n5300), .B1(n12674), .B2(n9182), .ZN(
        n5313) );
  INV_X1 U1833 ( .A(n5314), .ZN(n12672) );
  AOI22_X1 U1834 ( .A1(ram[878]), .A2(n5300), .B1(n12674), .B2(n9206), .ZN(
        n5314) );
  INV_X1 U1835 ( .A(n5315), .ZN(n12673) );
  AOI22_X1 U1836 ( .A1(ram[879]), .A2(n5300), .B1(n12674), .B2(n9230), .ZN(
        n5315) );
  INV_X1 U1837 ( .A(n5333), .ZN(n12624) );
  AOI22_X1 U1838 ( .A1(ram[896]), .A2(n5334), .B1(n12640), .B2(n8870), .ZN(
        n5333) );
  INV_X1 U1839 ( .A(n5335), .ZN(n12625) );
  AOI22_X1 U1840 ( .A1(ram[897]), .A2(n5334), .B1(n12640), .B2(n8894), .ZN(
        n5335) );
  INV_X1 U1841 ( .A(n5336), .ZN(n12626) );
  AOI22_X1 U1842 ( .A1(ram[898]), .A2(n5334), .B1(n12640), .B2(n8918), .ZN(
        n5336) );
  INV_X1 U1843 ( .A(n5337), .ZN(n12627) );
  AOI22_X1 U1844 ( .A1(ram[899]), .A2(n5334), .B1(n12640), .B2(n8942), .ZN(
        n5337) );
  INV_X1 U1845 ( .A(n5338), .ZN(n12628) );
  AOI22_X1 U1846 ( .A1(ram[900]), .A2(n5334), .B1(n12640), .B2(n8966), .ZN(
        n5338) );
  INV_X1 U1847 ( .A(n5339), .ZN(n12629) );
  AOI22_X1 U1848 ( .A1(ram[901]), .A2(n5334), .B1(n12640), .B2(n8990), .ZN(
        n5339) );
  INV_X1 U1849 ( .A(n5340), .ZN(n12630) );
  AOI22_X1 U1850 ( .A1(ram[902]), .A2(n5334), .B1(n12640), .B2(n9014), .ZN(
        n5340) );
  INV_X1 U1851 ( .A(n5341), .ZN(n12631) );
  AOI22_X1 U1852 ( .A1(ram[903]), .A2(n5334), .B1(n12640), .B2(n9038), .ZN(
        n5341) );
  INV_X1 U1853 ( .A(n5342), .ZN(n12632) );
  AOI22_X1 U1854 ( .A1(ram[904]), .A2(n5334), .B1(n12640), .B2(n9062), .ZN(
        n5342) );
  INV_X1 U1855 ( .A(n5343), .ZN(n12633) );
  AOI22_X1 U1856 ( .A1(ram[905]), .A2(n5334), .B1(n12640), .B2(n9086), .ZN(
        n5343) );
  INV_X1 U1857 ( .A(n5344), .ZN(n12634) );
  AOI22_X1 U1858 ( .A1(ram[906]), .A2(n5334), .B1(n12640), .B2(n9110), .ZN(
        n5344) );
  INV_X1 U1859 ( .A(n5345), .ZN(n12635) );
  AOI22_X1 U1860 ( .A1(ram[907]), .A2(n5334), .B1(n12640), .B2(n9134), .ZN(
        n5345) );
  INV_X1 U1861 ( .A(n5346), .ZN(n12636) );
  AOI22_X1 U1862 ( .A1(ram[908]), .A2(n5334), .B1(n12640), .B2(n9158), .ZN(
        n5346) );
  INV_X1 U1863 ( .A(n5347), .ZN(n12637) );
  AOI22_X1 U1864 ( .A1(ram[909]), .A2(n5334), .B1(n12640), .B2(n9182), .ZN(
        n5347) );
  INV_X1 U1865 ( .A(n5348), .ZN(n12638) );
  AOI22_X1 U1866 ( .A1(ram[910]), .A2(n5334), .B1(n12640), .B2(n9206), .ZN(
        n5348) );
  INV_X1 U1867 ( .A(n5349), .ZN(n12639) );
  AOI22_X1 U1868 ( .A1(ram[911]), .A2(n5334), .B1(n12640), .B2(n9230), .ZN(
        n5349) );
  INV_X1 U1869 ( .A(n5367), .ZN(n12590) );
  AOI22_X1 U1870 ( .A1(ram[928]), .A2(n5368), .B1(n12606), .B2(n8870), .ZN(
        n5367) );
  INV_X1 U1871 ( .A(n5369), .ZN(n12591) );
  AOI22_X1 U1872 ( .A1(ram[929]), .A2(n5368), .B1(n12606), .B2(n8894), .ZN(
        n5369) );
  INV_X1 U1873 ( .A(n5370), .ZN(n12592) );
  AOI22_X1 U1874 ( .A1(ram[930]), .A2(n5368), .B1(n12606), .B2(n8918), .ZN(
        n5370) );
  INV_X1 U1875 ( .A(n5371), .ZN(n12593) );
  AOI22_X1 U1876 ( .A1(ram[931]), .A2(n5368), .B1(n12606), .B2(n8942), .ZN(
        n5371) );
  INV_X1 U1877 ( .A(n5372), .ZN(n12594) );
  AOI22_X1 U1878 ( .A1(ram[932]), .A2(n5368), .B1(n12606), .B2(n8966), .ZN(
        n5372) );
  INV_X1 U1879 ( .A(n5373), .ZN(n12595) );
  AOI22_X1 U1880 ( .A1(ram[933]), .A2(n5368), .B1(n12606), .B2(n8990), .ZN(
        n5373) );
  INV_X1 U1881 ( .A(n5374), .ZN(n12596) );
  AOI22_X1 U1882 ( .A1(ram[934]), .A2(n5368), .B1(n12606), .B2(n9014), .ZN(
        n5374) );
  INV_X1 U1883 ( .A(n5375), .ZN(n12597) );
  AOI22_X1 U1884 ( .A1(ram[935]), .A2(n5368), .B1(n12606), .B2(n9038), .ZN(
        n5375) );
  INV_X1 U1885 ( .A(n5376), .ZN(n12598) );
  AOI22_X1 U1886 ( .A1(ram[936]), .A2(n5368), .B1(n12606), .B2(n9062), .ZN(
        n5376) );
  INV_X1 U1887 ( .A(n5377), .ZN(n12599) );
  AOI22_X1 U1888 ( .A1(ram[937]), .A2(n5368), .B1(n12606), .B2(n9086), .ZN(
        n5377) );
  INV_X1 U1889 ( .A(n5378), .ZN(n12600) );
  AOI22_X1 U1890 ( .A1(ram[938]), .A2(n5368), .B1(n12606), .B2(n9110), .ZN(
        n5378) );
  INV_X1 U1891 ( .A(n5379), .ZN(n12601) );
  AOI22_X1 U1892 ( .A1(ram[939]), .A2(n5368), .B1(n12606), .B2(n9134), .ZN(
        n5379) );
  INV_X1 U1893 ( .A(n5380), .ZN(n12602) );
  AOI22_X1 U1894 ( .A1(ram[940]), .A2(n5368), .B1(n12606), .B2(n9158), .ZN(
        n5380) );
  INV_X1 U1895 ( .A(n5381), .ZN(n12603) );
  AOI22_X1 U1896 ( .A1(ram[941]), .A2(n5368), .B1(n12606), .B2(n9182), .ZN(
        n5381) );
  INV_X1 U1897 ( .A(n5382), .ZN(n12604) );
  AOI22_X1 U1898 ( .A1(ram[942]), .A2(n5368), .B1(n12606), .B2(n9206), .ZN(
        n5382) );
  INV_X1 U1899 ( .A(n5383), .ZN(n12605) );
  AOI22_X1 U1900 ( .A1(ram[943]), .A2(n5368), .B1(n12606), .B2(n9230), .ZN(
        n5383) );
  INV_X1 U1901 ( .A(n5401), .ZN(n12556) );
  AOI22_X1 U1902 ( .A1(ram[960]), .A2(n5402), .B1(n12572), .B2(n8870), .ZN(
        n5401) );
  INV_X1 U1903 ( .A(n5403), .ZN(n12557) );
  AOI22_X1 U1904 ( .A1(ram[961]), .A2(n5402), .B1(n12572), .B2(n8894), .ZN(
        n5403) );
  INV_X1 U1905 ( .A(n5404), .ZN(n12558) );
  AOI22_X1 U1906 ( .A1(ram[962]), .A2(n5402), .B1(n12572), .B2(n8918), .ZN(
        n5404) );
  INV_X1 U1907 ( .A(n5405), .ZN(n12559) );
  AOI22_X1 U1908 ( .A1(ram[963]), .A2(n5402), .B1(n12572), .B2(n8942), .ZN(
        n5405) );
  INV_X1 U1909 ( .A(n5406), .ZN(n12560) );
  AOI22_X1 U1910 ( .A1(ram[964]), .A2(n5402), .B1(n12572), .B2(n8966), .ZN(
        n5406) );
  INV_X1 U1911 ( .A(n5407), .ZN(n12561) );
  AOI22_X1 U1912 ( .A1(ram[965]), .A2(n5402), .B1(n12572), .B2(n8990), .ZN(
        n5407) );
  INV_X1 U1913 ( .A(n5408), .ZN(n12562) );
  AOI22_X1 U1914 ( .A1(ram[966]), .A2(n5402), .B1(n12572), .B2(n9014), .ZN(
        n5408) );
  INV_X1 U1915 ( .A(n5409), .ZN(n12563) );
  AOI22_X1 U1916 ( .A1(ram[967]), .A2(n5402), .B1(n12572), .B2(n9038), .ZN(
        n5409) );
  INV_X1 U1917 ( .A(n5410), .ZN(n12564) );
  AOI22_X1 U1918 ( .A1(ram[968]), .A2(n5402), .B1(n12572), .B2(n9062), .ZN(
        n5410) );
  INV_X1 U1919 ( .A(n5411), .ZN(n12565) );
  AOI22_X1 U1920 ( .A1(ram[969]), .A2(n5402), .B1(n12572), .B2(n9086), .ZN(
        n5411) );
  INV_X1 U1921 ( .A(n5412), .ZN(n12566) );
  AOI22_X1 U1922 ( .A1(ram[970]), .A2(n5402), .B1(n12572), .B2(n9110), .ZN(
        n5412) );
  INV_X1 U1923 ( .A(n5413), .ZN(n12567) );
  AOI22_X1 U1924 ( .A1(ram[971]), .A2(n5402), .B1(n12572), .B2(n9134), .ZN(
        n5413) );
  INV_X1 U1925 ( .A(n5414), .ZN(n12568) );
  AOI22_X1 U1926 ( .A1(ram[972]), .A2(n5402), .B1(n12572), .B2(n9158), .ZN(
        n5414) );
  INV_X1 U1927 ( .A(n5415), .ZN(n12569) );
  AOI22_X1 U1928 ( .A1(ram[973]), .A2(n5402), .B1(n12572), .B2(n9182), .ZN(
        n5415) );
  INV_X1 U1929 ( .A(n5416), .ZN(n12570) );
  AOI22_X1 U1930 ( .A1(ram[974]), .A2(n5402), .B1(n12572), .B2(n9206), .ZN(
        n5416) );
  INV_X1 U1931 ( .A(n5417), .ZN(n12571) );
  AOI22_X1 U1932 ( .A1(ram[975]), .A2(n5402), .B1(n12572), .B2(n9230), .ZN(
        n5417) );
  INV_X1 U1933 ( .A(n5435), .ZN(n12522) );
  AOI22_X1 U1934 ( .A1(ram[992]), .A2(n5436), .B1(n12538), .B2(n8870), .ZN(
        n5435) );
  INV_X1 U1935 ( .A(n5437), .ZN(n12523) );
  AOI22_X1 U1936 ( .A1(ram[993]), .A2(n5436), .B1(n12538), .B2(n8894), .ZN(
        n5437) );
  INV_X1 U1937 ( .A(n5438), .ZN(n12524) );
  AOI22_X1 U1938 ( .A1(ram[994]), .A2(n5436), .B1(n12538), .B2(n8918), .ZN(
        n5438) );
  INV_X1 U1939 ( .A(n5439), .ZN(n12525) );
  AOI22_X1 U1940 ( .A1(ram[995]), .A2(n5436), .B1(n12538), .B2(n8942), .ZN(
        n5439) );
  INV_X1 U1941 ( .A(n5440), .ZN(n12526) );
  AOI22_X1 U1942 ( .A1(ram[996]), .A2(n5436), .B1(n12538), .B2(n8966), .ZN(
        n5440) );
  INV_X1 U1943 ( .A(n5441), .ZN(n12527) );
  AOI22_X1 U1944 ( .A1(ram[997]), .A2(n5436), .B1(n12538), .B2(n8990), .ZN(
        n5441) );
  INV_X1 U1945 ( .A(n5442), .ZN(n12528) );
  AOI22_X1 U1946 ( .A1(ram[998]), .A2(n5436), .B1(n12538), .B2(n9014), .ZN(
        n5442) );
  INV_X1 U1947 ( .A(n5443), .ZN(n12529) );
  AOI22_X1 U1948 ( .A1(ram[999]), .A2(n5436), .B1(n12538), .B2(n9038), .ZN(
        n5443) );
  INV_X1 U1949 ( .A(n5444), .ZN(n12530) );
  AOI22_X1 U1950 ( .A1(ram[1000]), .A2(n5436), .B1(n12538), .B2(n9062), .ZN(
        n5444) );
  INV_X1 U1951 ( .A(n5445), .ZN(n12531) );
  AOI22_X1 U1952 ( .A1(ram[1001]), .A2(n5436), .B1(n12538), .B2(n9086), .ZN(
        n5445) );
  INV_X1 U1953 ( .A(n5446), .ZN(n12532) );
  AOI22_X1 U1954 ( .A1(ram[1002]), .A2(n5436), .B1(n12538), .B2(n9110), .ZN(
        n5446) );
  INV_X1 U1955 ( .A(n5447), .ZN(n12533) );
  AOI22_X1 U1956 ( .A1(ram[1003]), .A2(n5436), .B1(n12538), .B2(n9134), .ZN(
        n5447) );
  INV_X1 U1957 ( .A(n5448), .ZN(n12534) );
  AOI22_X1 U1958 ( .A1(ram[1004]), .A2(n5436), .B1(n12538), .B2(n9158), .ZN(
        n5448) );
  INV_X1 U1959 ( .A(n5449), .ZN(n12535) );
  AOI22_X1 U1960 ( .A1(ram[1005]), .A2(n5436), .B1(n12538), .B2(n9182), .ZN(
        n5449) );
  INV_X1 U1961 ( .A(n5450), .ZN(n12536) );
  AOI22_X1 U1962 ( .A1(ram[1006]), .A2(n5436), .B1(n12538), .B2(n9206), .ZN(
        n5450) );
  INV_X1 U1963 ( .A(n5451), .ZN(n12537) );
  AOI22_X1 U1964 ( .A1(ram[1007]), .A2(n5436), .B1(n12538), .B2(n9230), .ZN(
        n5451) );
  INV_X1 U1965 ( .A(n5470), .ZN(n12488) );
  AOI22_X1 U1966 ( .A1(ram[1024]), .A2(n5471), .B1(n12504), .B2(n8869), .ZN(
        n5470) );
  INV_X1 U1967 ( .A(n5472), .ZN(n12489) );
  AOI22_X1 U1968 ( .A1(ram[1025]), .A2(n5471), .B1(n12504), .B2(n8893), .ZN(
        n5472) );
  INV_X1 U1969 ( .A(n5473), .ZN(n12490) );
  AOI22_X1 U1970 ( .A1(ram[1026]), .A2(n5471), .B1(n12504), .B2(n8917), .ZN(
        n5473) );
  INV_X1 U1971 ( .A(n5474), .ZN(n12491) );
  AOI22_X1 U1972 ( .A1(ram[1027]), .A2(n5471), .B1(n12504), .B2(n8941), .ZN(
        n5474) );
  INV_X1 U1973 ( .A(n5475), .ZN(n12492) );
  AOI22_X1 U1974 ( .A1(ram[1028]), .A2(n5471), .B1(n12504), .B2(n8965), .ZN(
        n5475) );
  INV_X1 U1975 ( .A(n5476), .ZN(n12493) );
  AOI22_X1 U1976 ( .A1(ram[1029]), .A2(n5471), .B1(n12504), .B2(n8989), .ZN(
        n5476) );
  INV_X1 U1977 ( .A(n5477), .ZN(n12494) );
  AOI22_X1 U1978 ( .A1(ram[1030]), .A2(n5471), .B1(n12504), .B2(n9013), .ZN(
        n5477) );
  INV_X1 U1979 ( .A(n5478), .ZN(n12495) );
  AOI22_X1 U1980 ( .A1(ram[1031]), .A2(n5471), .B1(n12504), .B2(n9037), .ZN(
        n5478) );
  INV_X1 U1981 ( .A(n5479), .ZN(n12496) );
  AOI22_X1 U1982 ( .A1(ram[1032]), .A2(n5471), .B1(n12504), .B2(n9061), .ZN(
        n5479) );
  INV_X1 U1983 ( .A(n5480), .ZN(n12497) );
  AOI22_X1 U1984 ( .A1(ram[1033]), .A2(n5471), .B1(n12504), .B2(n9085), .ZN(
        n5480) );
  INV_X1 U1985 ( .A(n5481), .ZN(n12498) );
  AOI22_X1 U1986 ( .A1(ram[1034]), .A2(n5471), .B1(n12504), .B2(n9109), .ZN(
        n5481) );
  INV_X1 U1987 ( .A(n5482), .ZN(n12499) );
  AOI22_X1 U1988 ( .A1(ram[1035]), .A2(n5471), .B1(n12504), .B2(n9133), .ZN(
        n5482) );
  INV_X1 U1989 ( .A(n5483), .ZN(n12500) );
  AOI22_X1 U1990 ( .A1(ram[1036]), .A2(n5471), .B1(n12504), .B2(n9157), .ZN(
        n5483) );
  INV_X1 U1991 ( .A(n5484), .ZN(n12501) );
  AOI22_X1 U1992 ( .A1(ram[1037]), .A2(n5471), .B1(n12504), .B2(n9181), .ZN(
        n5484) );
  INV_X1 U1993 ( .A(n5485), .ZN(n12502) );
  AOI22_X1 U1994 ( .A1(ram[1038]), .A2(n5471), .B1(n12504), .B2(n9205), .ZN(
        n5485) );
  INV_X1 U1995 ( .A(n5486), .ZN(n12503) );
  AOI22_X1 U1996 ( .A1(ram[1039]), .A2(n5471), .B1(n12504), .B2(n9229), .ZN(
        n5486) );
  INV_X1 U1997 ( .A(n5505), .ZN(n12454) );
  AOI22_X1 U1998 ( .A1(ram[1056]), .A2(n5506), .B1(n12470), .B2(n8869), .ZN(
        n5505) );
  INV_X1 U1999 ( .A(n5507), .ZN(n12455) );
  AOI22_X1 U2000 ( .A1(ram[1057]), .A2(n5506), .B1(n12470), .B2(n8893), .ZN(
        n5507) );
  INV_X1 U2001 ( .A(n5508), .ZN(n12456) );
  AOI22_X1 U2002 ( .A1(ram[1058]), .A2(n5506), .B1(n12470), .B2(n8917), .ZN(
        n5508) );
  INV_X1 U2003 ( .A(n5509), .ZN(n12457) );
  AOI22_X1 U2004 ( .A1(ram[1059]), .A2(n5506), .B1(n12470), .B2(n8941), .ZN(
        n5509) );
  INV_X1 U2005 ( .A(n5510), .ZN(n12458) );
  AOI22_X1 U2006 ( .A1(ram[1060]), .A2(n5506), .B1(n12470), .B2(n8965), .ZN(
        n5510) );
  INV_X1 U2007 ( .A(n5511), .ZN(n12459) );
  AOI22_X1 U2008 ( .A1(ram[1061]), .A2(n5506), .B1(n12470), .B2(n8989), .ZN(
        n5511) );
  INV_X1 U2009 ( .A(n5512), .ZN(n12460) );
  AOI22_X1 U2010 ( .A1(ram[1062]), .A2(n5506), .B1(n12470), .B2(n9013), .ZN(
        n5512) );
  INV_X1 U2011 ( .A(n5513), .ZN(n12461) );
  AOI22_X1 U2012 ( .A1(ram[1063]), .A2(n5506), .B1(n12470), .B2(n9037), .ZN(
        n5513) );
  INV_X1 U2013 ( .A(n5514), .ZN(n12462) );
  AOI22_X1 U2014 ( .A1(ram[1064]), .A2(n5506), .B1(n12470), .B2(n9061), .ZN(
        n5514) );
  INV_X1 U2015 ( .A(n5515), .ZN(n12463) );
  AOI22_X1 U2016 ( .A1(ram[1065]), .A2(n5506), .B1(n12470), .B2(n9085), .ZN(
        n5515) );
  INV_X1 U2017 ( .A(n5516), .ZN(n12464) );
  AOI22_X1 U2018 ( .A1(ram[1066]), .A2(n5506), .B1(n12470), .B2(n9109), .ZN(
        n5516) );
  INV_X1 U2019 ( .A(n5517), .ZN(n12465) );
  AOI22_X1 U2020 ( .A1(ram[1067]), .A2(n5506), .B1(n12470), .B2(n9133), .ZN(
        n5517) );
  INV_X1 U2021 ( .A(n5518), .ZN(n12466) );
  AOI22_X1 U2022 ( .A1(ram[1068]), .A2(n5506), .B1(n12470), .B2(n9157), .ZN(
        n5518) );
  INV_X1 U2023 ( .A(n5519), .ZN(n12467) );
  AOI22_X1 U2024 ( .A1(ram[1069]), .A2(n5506), .B1(n12470), .B2(n9181), .ZN(
        n5519) );
  INV_X1 U2025 ( .A(n5520), .ZN(n12468) );
  AOI22_X1 U2026 ( .A1(ram[1070]), .A2(n5506), .B1(n12470), .B2(n9205), .ZN(
        n5520) );
  INV_X1 U2027 ( .A(n5521), .ZN(n12469) );
  AOI22_X1 U2028 ( .A1(ram[1071]), .A2(n5506), .B1(n12470), .B2(n9229), .ZN(
        n5521) );
  INV_X1 U2029 ( .A(n5539), .ZN(n12420) );
  AOI22_X1 U2030 ( .A1(ram[1088]), .A2(n5540), .B1(n12436), .B2(n8869), .ZN(
        n5539) );
  INV_X1 U2031 ( .A(n5541), .ZN(n12421) );
  AOI22_X1 U2032 ( .A1(ram[1089]), .A2(n5540), .B1(n12436), .B2(n8893), .ZN(
        n5541) );
  INV_X1 U2033 ( .A(n5542), .ZN(n12422) );
  AOI22_X1 U2034 ( .A1(ram[1090]), .A2(n5540), .B1(n12436), .B2(n8917), .ZN(
        n5542) );
  INV_X1 U2035 ( .A(n5543), .ZN(n12423) );
  AOI22_X1 U2036 ( .A1(ram[1091]), .A2(n5540), .B1(n12436), .B2(n8941), .ZN(
        n5543) );
  INV_X1 U2037 ( .A(n5544), .ZN(n12424) );
  AOI22_X1 U2038 ( .A1(ram[1092]), .A2(n5540), .B1(n12436), .B2(n8965), .ZN(
        n5544) );
  INV_X1 U2039 ( .A(n5545), .ZN(n12425) );
  AOI22_X1 U2040 ( .A1(ram[1093]), .A2(n5540), .B1(n12436), .B2(n8989), .ZN(
        n5545) );
  INV_X1 U2041 ( .A(n5546), .ZN(n12426) );
  AOI22_X1 U2042 ( .A1(ram[1094]), .A2(n5540), .B1(n12436), .B2(n9013), .ZN(
        n5546) );
  INV_X1 U2043 ( .A(n5547), .ZN(n12427) );
  AOI22_X1 U2044 ( .A1(ram[1095]), .A2(n5540), .B1(n12436), .B2(n9037), .ZN(
        n5547) );
  INV_X1 U2045 ( .A(n5548), .ZN(n12428) );
  AOI22_X1 U2046 ( .A1(ram[1096]), .A2(n5540), .B1(n12436), .B2(n9061), .ZN(
        n5548) );
  INV_X1 U2047 ( .A(n5549), .ZN(n12429) );
  AOI22_X1 U2048 ( .A1(ram[1097]), .A2(n5540), .B1(n12436), .B2(n9085), .ZN(
        n5549) );
  INV_X1 U2049 ( .A(n5550), .ZN(n12430) );
  AOI22_X1 U2050 ( .A1(ram[1098]), .A2(n5540), .B1(n12436), .B2(n9109), .ZN(
        n5550) );
  INV_X1 U2051 ( .A(n5551), .ZN(n12431) );
  AOI22_X1 U2052 ( .A1(ram[1099]), .A2(n5540), .B1(n12436), .B2(n9133), .ZN(
        n5551) );
  INV_X1 U2053 ( .A(n5552), .ZN(n12432) );
  AOI22_X1 U2054 ( .A1(ram[1100]), .A2(n5540), .B1(n12436), .B2(n9157), .ZN(
        n5552) );
  INV_X1 U2055 ( .A(n5553), .ZN(n12433) );
  AOI22_X1 U2056 ( .A1(ram[1101]), .A2(n5540), .B1(n12436), .B2(n9181), .ZN(
        n5553) );
  INV_X1 U2057 ( .A(n5554), .ZN(n12434) );
  AOI22_X1 U2058 ( .A1(ram[1102]), .A2(n5540), .B1(n12436), .B2(n9205), .ZN(
        n5554) );
  INV_X1 U2059 ( .A(n5555), .ZN(n12435) );
  AOI22_X1 U2060 ( .A1(ram[1103]), .A2(n5540), .B1(n12436), .B2(n9229), .ZN(
        n5555) );
  INV_X1 U2061 ( .A(n5573), .ZN(n12386) );
  AOI22_X1 U2062 ( .A1(ram[1120]), .A2(n5574), .B1(n12402), .B2(n8869), .ZN(
        n5573) );
  INV_X1 U2063 ( .A(n5575), .ZN(n12387) );
  AOI22_X1 U2064 ( .A1(ram[1121]), .A2(n5574), .B1(n12402), .B2(n8893), .ZN(
        n5575) );
  INV_X1 U2065 ( .A(n5576), .ZN(n12388) );
  AOI22_X1 U2066 ( .A1(ram[1122]), .A2(n5574), .B1(n12402), .B2(n8917), .ZN(
        n5576) );
  INV_X1 U2067 ( .A(n5577), .ZN(n12389) );
  AOI22_X1 U2068 ( .A1(ram[1123]), .A2(n5574), .B1(n12402), .B2(n8941), .ZN(
        n5577) );
  INV_X1 U2069 ( .A(n5578), .ZN(n12390) );
  AOI22_X1 U2070 ( .A1(ram[1124]), .A2(n5574), .B1(n12402), .B2(n8965), .ZN(
        n5578) );
  INV_X1 U2071 ( .A(n5579), .ZN(n12391) );
  AOI22_X1 U2072 ( .A1(ram[1125]), .A2(n5574), .B1(n12402), .B2(n8989), .ZN(
        n5579) );
  INV_X1 U2073 ( .A(n5580), .ZN(n12392) );
  AOI22_X1 U2074 ( .A1(ram[1126]), .A2(n5574), .B1(n12402), .B2(n9013), .ZN(
        n5580) );
  INV_X1 U2075 ( .A(n5581), .ZN(n12393) );
  AOI22_X1 U2076 ( .A1(ram[1127]), .A2(n5574), .B1(n12402), .B2(n9037), .ZN(
        n5581) );
  INV_X1 U2077 ( .A(n5582), .ZN(n12394) );
  AOI22_X1 U2078 ( .A1(ram[1128]), .A2(n5574), .B1(n12402), .B2(n9061), .ZN(
        n5582) );
  INV_X1 U2079 ( .A(n5583), .ZN(n12395) );
  AOI22_X1 U2080 ( .A1(ram[1129]), .A2(n5574), .B1(n12402), .B2(n9085), .ZN(
        n5583) );
  INV_X1 U2081 ( .A(n5584), .ZN(n12396) );
  AOI22_X1 U2082 ( .A1(ram[1130]), .A2(n5574), .B1(n12402), .B2(n9109), .ZN(
        n5584) );
  INV_X1 U2083 ( .A(n5585), .ZN(n12397) );
  AOI22_X1 U2084 ( .A1(ram[1131]), .A2(n5574), .B1(n12402), .B2(n9133), .ZN(
        n5585) );
  INV_X1 U2085 ( .A(n5586), .ZN(n12398) );
  AOI22_X1 U2086 ( .A1(ram[1132]), .A2(n5574), .B1(n12402), .B2(n9157), .ZN(
        n5586) );
  INV_X1 U2087 ( .A(n5587), .ZN(n12399) );
  AOI22_X1 U2088 ( .A1(ram[1133]), .A2(n5574), .B1(n12402), .B2(n9181), .ZN(
        n5587) );
  INV_X1 U2089 ( .A(n5588), .ZN(n12400) );
  AOI22_X1 U2090 ( .A1(ram[1134]), .A2(n5574), .B1(n12402), .B2(n9205), .ZN(
        n5588) );
  INV_X1 U2091 ( .A(n5589), .ZN(n12401) );
  AOI22_X1 U2092 ( .A1(ram[1135]), .A2(n5574), .B1(n12402), .B2(n9229), .ZN(
        n5589) );
  INV_X1 U2093 ( .A(n5607), .ZN(n12352) );
  AOI22_X1 U2094 ( .A1(ram[1152]), .A2(n5608), .B1(n12368), .B2(n8869), .ZN(
        n5607) );
  INV_X1 U2095 ( .A(n5609), .ZN(n12353) );
  AOI22_X1 U2096 ( .A1(ram[1153]), .A2(n5608), .B1(n12368), .B2(n8893), .ZN(
        n5609) );
  INV_X1 U2097 ( .A(n5610), .ZN(n12354) );
  AOI22_X1 U2098 ( .A1(ram[1154]), .A2(n5608), .B1(n12368), .B2(n8917), .ZN(
        n5610) );
  INV_X1 U2099 ( .A(n5611), .ZN(n12355) );
  AOI22_X1 U2100 ( .A1(ram[1155]), .A2(n5608), .B1(n12368), .B2(n8941), .ZN(
        n5611) );
  INV_X1 U2101 ( .A(n5612), .ZN(n12356) );
  AOI22_X1 U2102 ( .A1(ram[1156]), .A2(n5608), .B1(n12368), .B2(n8965), .ZN(
        n5612) );
  INV_X1 U2103 ( .A(n5613), .ZN(n12357) );
  AOI22_X1 U2104 ( .A1(ram[1157]), .A2(n5608), .B1(n12368), .B2(n8989), .ZN(
        n5613) );
  INV_X1 U2105 ( .A(n5614), .ZN(n12358) );
  AOI22_X1 U2106 ( .A1(ram[1158]), .A2(n5608), .B1(n12368), .B2(n9013), .ZN(
        n5614) );
  INV_X1 U2107 ( .A(n5615), .ZN(n12359) );
  AOI22_X1 U2108 ( .A1(ram[1159]), .A2(n5608), .B1(n12368), .B2(n9037), .ZN(
        n5615) );
  INV_X1 U2109 ( .A(n5616), .ZN(n12360) );
  AOI22_X1 U2110 ( .A1(ram[1160]), .A2(n5608), .B1(n12368), .B2(n9061), .ZN(
        n5616) );
  INV_X1 U2111 ( .A(n5617), .ZN(n12361) );
  AOI22_X1 U2112 ( .A1(ram[1161]), .A2(n5608), .B1(n12368), .B2(n9085), .ZN(
        n5617) );
  INV_X1 U2113 ( .A(n5618), .ZN(n12362) );
  AOI22_X1 U2114 ( .A1(ram[1162]), .A2(n5608), .B1(n12368), .B2(n9109), .ZN(
        n5618) );
  INV_X1 U2115 ( .A(n5619), .ZN(n12363) );
  AOI22_X1 U2116 ( .A1(ram[1163]), .A2(n5608), .B1(n12368), .B2(n9133), .ZN(
        n5619) );
  INV_X1 U2117 ( .A(n5620), .ZN(n12364) );
  AOI22_X1 U2118 ( .A1(ram[1164]), .A2(n5608), .B1(n12368), .B2(n9157), .ZN(
        n5620) );
  INV_X1 U2119 ( .A(n5621), .ZN(n12365) );
  AOI22_X1 U2120 ( .A1(ram[1165]), .A2(n5608), .B1(n12368), .B2(n9181), .ZN(
        n5621) );
  INV_X1 U2121 ( .A(n5622), .ZN(n12366) );
  AOI22_X1 U2122 ( .A1(ram[1166]), .A2(n5608), .B1(n12368), .B2(n9205), .ZN(
        n5622) );
  INV_X1 U2123 ( .A(n5623), .ZN(n12367) );
  AOI22_X1 U2124 ( .A1(ram[1167]), .A2(n5608), .B1(n12368), .B2(n9229), .ZN(
        n5623) );
  INV_X1 U2125 ( .A(n5641), .ZN(n12318) );
  AOI22_X1 U2126 ( .A1(ram[1184]), .A2(n5642), .B1(n12334), .B2(n8869), .ZN(
        n5641) );
  INV_X1 U2127 ( .A(n5643), .ZN(n12319) );
  AOI22_X1 U2128 ( .A1(ram[1185]), .A2(n5642), .B1(n12334), .B2(n8893), .ZN(
        n5643) );
  INV_X1 U2129 ( .A(n5644), .ZN(n12320) );
  AOI22_X1 U2130 ( .A1(ram[1186]), .A2(n5642), .B1(n12334), .B2(n8917), .ZN(
        n5644) );
  INV_X1 U2131 ( .A(n5645), .ZN(n12321) );
  AOI22_X1 U2132 ( .A1(ram[1187]), .A2(n5642), .B1(n12334), .B2(n8941), .ZN(
        n5645) );
  INV_X1 U2133 ( .A(n5646), .ZN(n12322) );
  AOI22_X1 U2134 ( .A1(ram[1188]), .A2(n5642), .B1(n12334), .B2(n8965), .ZN(
        n5646) );
  INV_X1 U2135 ( .A(n5647), .ZN(n12323) );
  AOI22_X1 U2136 ( .A1(ram[1189]), .A2(n5642), .B1(n12334), .B2(n8989), .ZN(
        n5647) );
  INV_X1 U2137 ( .A(n5648), .ZN(n12324) );
  AOI22_X1 U2138 ( .A1(ram[1190]), .A2(n5642), .B1(n12334), .B2(n9013), .ZN(
        n5648) );
  INV_X1 U2139 ( .A(n5649), .ZN(n12325) );
  AOI22_X1 U2140 ( .A1(ram[1191]), .A2(n5642), .B1(n12334), .B2(n9037), .ZN(
        n5649) );
  INV_X1 U2141 ( .A(n5650), .ZN(n12326) );
  AOI22_X1 U2142 ( .A1(ram[1192]), .A2(n5642), .B1(n12334), .B2(n9061), .ZN(
        n5650) );
  INV_X1 U2143 ( .A(n5651), .ZN(n12327) );
  AOI22_X1 U2144 ( .A1(ram[1193]), .A2(n5642), .B1(n12334), .B2(n9085), .ZN(
        n5651) );
  INV_X1 U2145 ( .A(n5652), .ZN(n12328) );
  AOI22_X1 U2146 ( .A1(ram[1194]), .A2(n5642), .B1(n12334), .B2(n9109), .ZN(
        n5652) );
  INV_X1 U2147 ( .A(n5653), .ZN(n12329) );
  AOI22_X1 U2148 ( .A1(ram[1195]), .A2(n5642), .B1(n12334), .B2(n9133), .ZN(
        n5653) );
  INV_X1 U2149 ( .A(n5654), .ZN(n12330) );
  AOI22_X1 U2150 ( .A1(ram[1196]), .A2(n5642), .B1(n12334), .B2(n9157), .ZN(
        n5654) );
  INV_X1 U2151 ( .A(n5655), .ZN(n12331) );
  AOI22_X1 U2152 ( .A1(ram[1197]), .A2(n5642), .B1(n12334), .B2(n9181), .ZN(
        n5655) );
  INV_X1 U2153 ( .A(n5656), .ZN(n12332) );
  AOI22_X1 U2154 ( .A1(ram[1198]), .A2(n5642), .B1(n12334), .B2(n9205), .ZN(
        n5656) );
  INV_X1 U2155 ( .A(n5657), .ZN(n12333) );
  AOI22_X1 U2156 ( .A1(ram[1199]), .A2(n5642), .B1(n12334), .B2(n9229), .ZN(
        n5657) );
  INV_X1 U2157 ( .A(n5675), .ZN(n12284) );
  AOI22_X1 U2158 ( .A1(ram[1216]), .A2(n5676), .B1(n12300), .B2(n8868), .ZN(
        n5675) );
  INV_X1 U2159 ( .A(n5677), .ZN(n12285) );
  AOI22_X1 U2160 ( .A1(ram[1217]), .A2(n5676), .B1(n12300), .B2(n8892), .ZN(
        n5677) );
  INV_X1 U2161 ( .A(n5678), .ZN(n12286) );
  AOI22_X1 U2162 ( .A1(ram[1218]), .A2(n5676), .B1(n12300), .B2(n8916), .ZN(
        n5678) );
  INV_X1 U2163 ( .A(n5679), .ZN(n12287) );
  AOI22_X1 U2164 ( .A1(ram[1219]), .A2(n5676), .B1(n12300), .B2(n8940), .ZN(
        n5679) );
  INV_X1 U2165 ( .A(n5680), .ZN(n12288) );
  AOI22_X1 U2166 ( .A1(ram[1220]), .A2(n5676), .B1(n12300), .B2(n8964), .ZN(
        n5680) );
  INV_X1 U2167 ( .A(n5681), .ZN(n12289) );
  AOI22_X1 U2168 ( .A1(ram[1221]), .A2(n5676), .B1(n12300), .B2(n8988), .ZN(
        n5681) );
  INV_X1 U2169 ( .A(n5682), .ZN(n12290) );
  AOI22_X1 U2170 ( .A1(ram[1222]), .A2(n5676), .B1(n12300), .B2(n9012), .ZN(
        n5682) );
  INV_X1 U2171 ( .A(n5683), .ZN(n12291) );
  AOI22_X1 U2172 ( .A1(ram[1223]), .A2(n5676), .B1(n12300), .B2(n9036), .ZN(
        n5683) );
  INV_X1 U2173 ( .A(n5684), .ZN(n12292) );
  AOI22_X1 U2174 ( .A1(ram[1224]), .A2(n5676), .B1(n12300), .B2(n9060), .ZN(
        n5684) );
  INV_X1 U2175 ( .A(n5685), .ZN(n12293) );
  AOI22_X1 U2176 ( .A1(ram[1225]), .A2(n5676), .B1(n12300), .B2(n9084), .ZN(
        n5685) );
  INV_X1 U2177 ( .A(n5686), .ZN(n12294) );
  AOI22_X1 U2178 ( .A1(ram[1226]), .A2(n5676), .B1(n12300), .B2(n9108), .ZN(
        n5686) );
  INV_X1 U2179 ( .A(n5687), .ZN(n12295) );
  AOI22_X1 U2180 ( .A1(ram[1227]), .A2(n5676), .B1(n12300), .B2(n9132), .ZN(
        n5687) );
  INV_X1 U2181 ( .A(n5688), .ZN(n12296) );
  AOI22_X1 U2182 ( .A1(ram[1228]), .A2(n5676), .B1(n12300), .B2(n9156), .ZN(
        n5688) );
  INV_X1 U2183 ( .A(n5689), .ZN(n12297) );
  AOI22_X1 U2184 ( .A1(ram[1229]), .A2(n5676), .B1(n12300), .B2(n9180), .ZN(
        n5689) );
  INV_X1 U2185 ( .A(n5690), .ZN(n12298) );
  AOI22_X1 U2186 ( .A1(ram[1230]), .A2(n5676), .B1(n12300), .B2(n9204), .ZN(
        n5690) );
  INV_X1 U2187 ( .A(n5691), .ZN(n12299) );
  AOI22_X1 U2188 ( .A1(ram[1231]), .A2(n5676), .B1(n12300), .B2(n9228), .ZN(
        n5691) );
  INV_X1 U2189 ( .A(n5709), .ZN(n12250) );
  AOI22_X1 U2190 ( .A1(ram[1248]), .A2(n5710), .B1(n12266), .B2(n8868), .ZN(
        n5709) );
  INV_X1 U2191 ( .A(n5711), .ZN(n12251) );
  AOI22_X1 U2192 ( .A1(ram[1249]), .A2(n5710), .B1(n12266), .B2(n8892), .ZN(
        n5711) );
  INV_X1 U2193 ( .A(n5712), .ZN(n12252) );
  AOI22_X1 U2194 ( .A1(ram[1250]), .A2(n5710), .B1(n12266), .B2(n8916), .ZN(
        n5712) );
  INV_X1 U2195 ( .A(n5713), .ZN(n12253) );
  AOI22_X1 U2196 ( .A1(ram[1251]), .A2(n5710), .B1(n12266), .B2(n8940), .ZN(
        n5713) );
  INV_X1 U2197 ( .A(n5714), .ZN(n12254) );
  AOI22_X1 U2198 ( .A1(ram[1252]), .A2(n5710), .B1(n12266), .B2(n8964), .ZN(
        n5714) );
  INV_X1 U2199 ( .A(n5715), .ZN(n12255) );
  AOI22_X1 U2200 ( .A1(ram[1253]), .A2(n5710), .B1(n12266), .B2(n8988), .ZN(
        n5715) );
  INV_X1 U2201 ( .A(n5716), .ZN(n12256) );
  AOI22_X1 U2202 ( .A1(ram[1254]), .A2(n5710), .B1(n12266), .B2(n9012), .ZN(
        n5716) );
  INV_X1 U2203 ( .A(n5717), .ZN(n12257) );
  AOI22_X1 U2204 ( .A1(ram[1255]), .A2(n5710), .B1(n12266), .B2(n9036), .ZN(
        n5717) );
  INV_X1 U2205 ( .A(n5718), .ZN(n12258) );
  AOI22_X1 U2206 ( .A1(ram[1256]), .A2(n5710), .B1(n12266), .B2(n9060), .ZN(
        n5718) );
  INV_X1 U2207 ( .A(n5719), .ZN(n12259) );
  AOI22_X1 U2208 ( .A1(ram[1257]), .A2(n5710), .B1(n12266), .B2(n9084), .ZN(
        n5719) );
  INV_X1 U2209 ( .A(n5720), .ZN(n12260) );
  AOI22_X1 U2210 ( .A1(ram[1258]), .A2(n5710), .B1(n12266), .B2(n9108), .ZN(
        n5720) );
  INV_X1 U2211 ( .A(n5721), .ZN(n12261) );
  AOI22_X1 U2212 ( .A1(ram[1259]), .A2(n5710), .B1(n12266), .B2(n9132), .ZN(
        n5721) );
  INV_X1 U2213 ( .A(n5722), .ZN(n12262) );
  AOI22_X1 U2214 ( .A1(ram[1260]), .A2(n5710), .B1(n12266), .B2(n9156), .ZN(
        n5722) );
  INV_X1 U2215 ( .A(n5723), .ZN(n12263) );
  AOI22_X1 U2216 ( .A1(ram[1261]), .A2(n5710), .B1(n12266), .B2(n9180), .ZN(
        n5723) );
  INV_X1 U2217 ( .A(n5724), .ZN(n12264) );
  AOI22_X1 U2218 ( .A1(ram[1262]), .A2(n5710), .B1(n12266), .B2(n9204), .ZN(
        n5724) );
  INV_X1 U2219 ( .A(n5725), .ZN(n12265) );
  AOI22_X1 U2220 ( .A1(ram[1263]), .A2(n5710), .B1(n12266), .B2(n9228), .ZN(
        n5725) );
  INV_X1 U2221 ( .A(n5744), .ZN(n12216) );
  AOI22_X1 U2222 ( .A1(ram[1280]), .A2(n5745), .B1(n12232), .B2(n8868), .ZN(
        n5744) );
  INV_X1 U2223 ( .A(n5746), .ZN(n12217) );
  AOI22_X1 U2224 ( .A1(ram[1281]), .A2(n5745), .B1(n12232), .B2(n8892), .ZN(
        n5746) );
  INV_X1 U2225 ( .A(n5747), .ZN(n12218) );
  AOI22_X1 U2226 ( .A1(ram[1282]), .A2(n5745), .B1(n12232), .B2(n8916), .ZN(
        n5747) );
  INV_X1 U2227 ( .A(n5748), .ZN(n12219) );
  AOI22_X1 U2228 ( .A1(ram[1283]), .A2(n5745), .B1(n12232), .B2(n8940), .ZN(
        n5748) );
  INV_X1 U2229 ( .A(n5749), .ZN(n12220) );
  AOI22_X1 U2230 ( .A1(ram[1284]), .A2(n5745), .B1(n12232), .B2(n8964), .ZN(
        n5749) );
  INV_X1 U2231 ( .A(n5750), .ZN(n12221) );
  AOI22_X1 U2232 ( .A1(ram[1285]), .A2(n5745), .B1(n12232), .B2(n8988), .ZN(
        n5750) );
  INV_X1 U2233 ( .A(n5751), .ZN(n12222) );
  AOI22_X1 U2234 ( .A1(ram[1286]), .A2(n5745), .B1(n12232), .B2(n9012), .ZN(
        n5751) );
  INV_X1 U2235 ( .A(n5752), .ZN(n12223) );
  AOI22_X1 U2236 ( .A1(ram[1287]), .A2(n5745), .B1(n12232), .B2(n9036), .ZN(
        n5752) );
  INV_X1 U2237 ( .A(n5753), .ZN(n12224) );
  AOI22_X1 U2238 ( .A1(ram[1288]), .A2(n5745), .B1(n12232), .B2(n9060), .ZN(
        n5753) );
  INV_X1 U2239 ( .A(n5754), .ZN(n12225) );
  AOI22_X1 U2240 ( .A1(ram[1289]), .A2(n5745), .B1(n12232), .B2(n9084), .ZN(
        n5754) );
  INV_X1 U2241 ( .A(n5755), .ZN(n12226) );
  AOI22_X1 U2242 ( .A1(ram[1290]), .A2(n5745), .B1(n12232), .B2(n9108), .ZN(
        n5755) );
  INV_X1 U2243 ( .A(n5756), .ZN(n12227) );
  AOI22_X1 U2244 ( .A1(ram[1291]), .A2(n5745), .B1(n12232), .B2(n9132), .ZN(
        n5756) );
  INV_X1 U2245 ( .A(n5757), .ZN(n12228) );
  AOI22_X1 U2246 ( .A1(ram[1292]), .A2(n5745), .B1(n12232), .B2(n9156), .ZN(
        n5757) );
  INV_X1 U2247 ( .A(n5758), .ZN(n12229) );
  AOI22_X1 U2248 ( .A1(ram[1293]), .A2(n5745), .B1(n12232), .B2(n9180), .ZN(
        n5758) );
  INV_X1 U2249 ( .A(n5759), .ZN(n12230) );
  AOI22_X1 U2250 ( .A1(ram[1294]), .A2(n5745), .B1(n12232), .B2(n9204), .ZN(
        n5759) );
  INV_X1 U2251 ( .A(n5760), .ZN(n12231) );
  AOI22_X1 U2252 ( .A1(ram[1295]), .A2(n5745), .B1(n12232), .B2(n9228), .ZN(
        n5760) );
  INV_X1 U2253 ( .A(n5779), .ZN(n12182) );
  AOI22_X1 U2254 ( .A1(ram[1312]), .A2(n5780), .B1(n12198), .B2(n8868), .ZN(
        n5779) );
  INV_X1 U2255 ( .A(n5781), .ZN(n12183) );
  AOI22_X1 U2256 ( .A1(ram[1313]), .A2(n5780), .B1(n12198), .B2(n8892), .ZN(
        n5781) );
  INV_X1 U2257 ( .A(n5782), .ZN(n12184) );
  AOI22_X1 U2258 ( .A1(ram[1314]), .A2(n5780), .B1(n12198), .B2(n8916), .ZN(
        n5782) );
  INV_X1 U2259 ( .A(n5783), .ZN(n12185) );
  AOI22_X1 U2260 ( .A1(ram[1315]), .A2(n5780), .B1(n12198), .B2(n8940), .ZN(
        n5783) );
  INV_X1 U2261 ( .A(n5784), .ZN(n12186) );
  AOI22_X1 U2262 ( .A1(ram[1316]), .A2(n5780), .B1(n12198), .B2(n8964), .ZN(
        n5784) );
  INV_X1 U2263 ( .A(n5785), .ZN(n12187) );
  AOI22_X1 U2264 ( .A1(ram[1317]), .A2(n5780), .B1(n12198), .B2(n8988), .ZN(
        n5785) );
  INV_X1 U2265 ( .A(n5786), .ZN(n12188) );
  AOI22_X1 U2266 ( .A1(ram[1318]), .A2(n5780), .B1(n12198), .B2(n9012), .ZN(
        n5786) );
  INV_X1 U2267 ( .A(n5787), .ZN(n12189) );
  AOI22_X1 U2268 ( .A1(ram[1319]), .A2(n5780), .B1(n12198), .B2(n9036), .ZN(
        n5787) );
  INV_X1 U2269 ( .A(n5788), .ZN(n12190) );
  AOI22_X1 U2270 ( .A1(ram[1320]), .A2(n5780), .B1(n12198), .B2(n9060), .ZN(
        n5788) );
  INV_X1 U2271 ( .A(n5789), .ZN(n12191) );
  AOI22_X1 U2272 ( .A1(ram[1321]), .A2(n5780), .B1(n12198), .B2(n9084), .ZN(
        n5789) );
  INV_X1 U2273 ( .A(n5790), .ZN(n12192) );
  AOI22_X1 U2274 ( .A1(ram[1322]), .A2(n5780), .B1(n12198), .B2(n9108), .ZN(
        n5790) );
  INV_X1 U2275 ( .A(n5791), .ZN(n12193) );
  AOI22_X1 U2276 ( .A1(ram[1323]), .A2(n5780), .B1(n12198), .B2(n9132), .ZN(
        n5791) );
  INV_X1 U2277 ( .A(n5792), .ZN(n12194) );
  AOI22_X1 U2278 ( .A1(ram[1324]), .A2(n5780), .B1(n12198), .B2(n9156), .ZN(
        n5792) );
  INV_X1 U2279 ( .A(n5793), .ZN(n12195) );
  AOI22_X1 U2280 ( .A1(ram[1325]), .A2(n5780), .B1(n12198), .B2(n9180), .ZN(
        n5793) );
  INV_X1 U2281 ( .A(n5794), .ZN(n12196) );
  AOI22_X1 U2282 ( .A1(ram[1326]), .A2(n5780), .B1(n12198), .B2(n9204), .ZN(
        n5794) );
  INV_X1 U2283 ( .A(n5795), .ZN(n12197) );
  AOI22_X1 U2284 ( .A1(ram[1327]), .A2(n5780), .B1(n12198), .B2(n9228), .ZN(
        n5795) );
  INV_X1 U2285 ( .A(n5813), .ZN(n12148) );
  AOI22_X1 U2286 ( .A1(ram[1344]), .A2(n5814), .B1(n12164), .B2(n8868), .ZN(
        n5813) );
  INV_X1 U2287 ( .A(n5815), .ZN(n12149) );
  AOI22_X1 U2288 ( .A1(ram[1345]), .A2(n5814), .B1(n12164), .B2(n8892), .ZN(
        n5815) );
  INV_X1 U2289 ( .A(n5816), .ZN(n12150) );
  AOI22_X1 U2290 ( .A1(ram[1346]), .A2(n5814), .B1(n12164), .B2(n8916), .ZN(
        n5816) );
  INV_X1 U2291 ( .A(n5817), .ZN(n12151) );
  AOI22_X1 U2292 ( .A1(ram[1347]), .A2(n5814), .B1(n12164), .B2(n8940), .ZN(
        n5817) );
  INV_X1 U2293 ( .A(n5818), .ZN(n12152) );
  AOI22_X1 U2294 ( .A1(ram[1348]), .A2(n5814), .B1(n12164), .B2(n8964), .ZN(
        n5818) );
  INV_X1 U2295 ( .A(n5819), .ZN(n12153) );
  AOI22_X1 U2296 ( .A1(ram[1349]), .A2(n5814), .B1(n12164), .B2(n8988), .ZN(
        n5819) );
  INV_X1 U2297 ( .A(n5820), .ZN(n12154) );
  AOI22_X1 U2298 ( .A1(ram[1350]), .A2(n5814), .B1(n12164), .B2(n9012), .ZN(
        n5820) );
  INV_X1 U2299 ( .A(n5821), .ZN(n12155) );
  AOI22_X1 U2300 ( .A1(ram[1351]), .A2(n5814), .B1(n12164), .B2(n9036), .ZN(
        n5821) );
  INV_X1 U2301 ( .A(n5822), .ZN(n12156) );
  AOI22_X1 U2302 ( .A1(ram[1352]), .A2(n5814), .B1(n12164), .B2(n9060), .ZN(
        n5822) );
  INV_X1 U2303 ( .A(n5823), .ZN(n12157) );
  AOI22_X1 U2304 ( .A1(ram[1353]), .A2(n5814), .B1(n12164), .B2(n9084), .ZN(
        n5823) );
  INV_X1 U2305 ( .A(n5824), .ZN(n12158) );
  AOI22_X1 U2306 ( .A1(ram[1354]), .A2(n5814), .B1(n12164), .B2(n9108), .ZN(
        n5824) );
  INV_X1 U2307 ( .A(n5825), .ZN(n12159) );
  AOI22_X1 U2308 ( .A1(ram[1355]), .A2(n5814), .B1(n12164), .B2(n9132), .ZN(
        n5825) );
  INV_X1 U2309 ( .A(n5826), .ZN(n12160) );
  AOI22_X1 U2310 ( .A1(ram[1356]), .A2(n5814), .B1(n12164), .B2(n9156), .ZN(
        n5826) );
  INV_X1 U2311 ( .A(n5827), .ZN(n12161) );
  AOI22_X1 U2312 ( .A1(ram[1357]), .A2(n5814), .B1(n12164), .B2(n9180), .ZN(
        n5827) );
  INV_X1 U2313 ( .A(n5828), .ZN(n12162) );
  AOI22_X1 U2314 ( .A1(ram[1358]), .A2(n5814), .B1(n12164), .B2(n9204), .ZN(
        n5828) );
  INV_X1 U2315 ( .A(n5829), .ZN(n12163) );
  AOI22_X1 U2316 ( .A1(ram[1359]), .A2(n5814), .B1(n12164), .B2(n9228), .ZN(
        n5829) );
  INV_X1 U2317 ( .A(n5847), .ZN(n12114) );
  AOI22_X1 U2318 ( .A1(ram[1376]), .A2(n5848), .B1(n12130), .B2(n8868), .ZN(
        n5847) );
  INV_X1 U2319 ( .A(n5849), .ZN(n12115) );
  AOI22_X1 U2320 ( .A1(ram[1377]), .A2(n5848), .B1(n12130), .B2(n8892), .ZN(
        n5849) );
  INV_X1 U2321 ( .A(n5850), .ZN(n12116) );
  AOI22_X1 U2322 ( .A1(ram[1378]), .A2(n5848), .B1(n12130), .B2(n8916), .ZN(
        n5850) );
  INV_X1 U2323 ( .A(n5851), .ZN(n12117) );
  AOI22_X1 U2324 ( .A1(ram[1379]), .A2(n5848), .B1(n12130), .B2(n8940), .ZN(
        n5851) );
  INV_X1 U2325 ( .A(n5852), .ZN(n12118) );
  AOI22_X1 U2326 ( .A1(ram[1380]), .A2(n5848), .B1(n12130), .B2(n8964), .ZN(
        n5852) );
  INV_X1 U2327 ( .A(n5853), .ZN(n12119) );
  AOI22_X1 U2328 ( .A1(ram[1381]), .A2(n5848), .B1(n12130), .B2(n8988), .ZN(
        n5853) );
  INV_X1 U2329 ( .A(n5854), .ZN(n12120) );
  AOI22_X1 U2330 ( .A1(ram[1382]), .A2(n5848), .B1(n12130), .B2(n9012), .ZN(
        n5854) );
  INV_X1 U2331 ( .A(n5855), .ZN(n12121) );
  AOI22_X1 U2332 ( .A1(ram[1383]), .A2(n5848), .B1(n12130), .B2(n9036), .ZN(
        n5855) );
  INV_X1 U2333 ( .A(n5856), .ZN(n12122) );
  AOI22_X1 U2334 ( .A1(ram[1384]), .A2(n5848), .B1(n12130), .B2(n9060), .ZN(
        n5856) );
  INV_X1 U2335 ( .A(n5857), .ZN(n12123) );
  AOI22_X1 U2336 ( .A1(ram[1385]), .A2(n5848), .B1(n12130), .B2(n9084), .ZN(
        n5857) );
  INV_X1 U2337 ( .A(n5858), .ZN(n12124) );
  AOI22_X1 U2338 ( .A1(ram[1386]), .A2(n5848), .B1(n12130), .B2(n9108), .ZN(
        n5858) );
  INV_X1 U2339 ( .A(n5859), .ZN(n12125) );
  AOI22_X1 U2340 ( .A1(ram[1387]), .A2(n5848), .B1(n12130), .B2(n9132), .ZN(
        n5859) );
  INV_X1 U2341 ( .A(n5860), .ZN(n12126) );
  AOI22_X1 U2342 ( .A1(ram[1388]), .A2(n5848), .B1(n12130), .B2(n9156), .ZN(
        n5860) );
  INV_X1 U2343 ( .A(n5861), .ZN(n12127) );
  AOI22_X1 U2344 ( .A1(ram[1389]), .A2(n5848), .B1(n12130), .B2(n9180), .ZN(
        n5861) );
  INV_X1 U2345 ( .A(n5862), .ZN(n12128) );
  AOI22_X1 U2346 ( .A1(ram[1390]), .A2(n5848), .B1(n12130), .B2(n9204), .ZN(
        n5862) );
  INV_X1 U2347 ( .A(n5863), .ZN(n12129) );
  AOI22_X1 U2348 ( .A1(ram[1391]), .A2(n5848), .B1(n12130), .B2(n9228), .ZN(
        n5863) );
  INV_X1 U2349 ( .A(n5881), .ZN(n12080) );
  AOI22_X1 U2350 ( .A1(ram[1408]), .A2(n5882), .B1(n12096), .B2(n8867), .ZN(
        n5881) );
  INV_X1 U2351 ( .A(n5883), .ZN(n12081) );
  AOI22_X1 U2352 ( .A1(ram[1409]), .A2(n5882), .B1(n12096), .B2(n8891), .ZN(
        n5883) );
  INV_X1 U2353 ( .A(n5884), .ZN(n12082) );
  AOI22_X1 U2354 ( .A1(ram[1410]), .A2(n5882), .B1(n12096), .B2(n8915), .ZN(
        n5884) );
  INV_X1 U2355 ( .A(n5885), .ZN(n12083) );
  AOI22_X1 U2356 ( .A1(ram[1411]), .A2(n5882), .B1(n12096), .B2(n8939), .ZN(
        n5885) );
  INV_X1 U2357 ( .A(n5886), .ZN(n12084) );
  AOI22_X1 U2358 ( .A1(ram[1412]), .A2(n5882), .B1(n12096), .B2(n8963), .ZN(
        n5886) );
  INV_X1 U2359 ( .A(n5887), .ZN(n12085) );
  AOI22_X1 U2360 ( .A1(ram[1413]), .A2(n5882), .B1(n12096), .B2(n8987), .ZN(
        n5887) );
  INV_X1 U2361 ( .A(n5888), .ZN(n12086) );
  AOI22_X1 U2362 ( .A1(ram[1414]), .A2(n5882), .B1(n12096), .B2(n9011), .ZN(
        n5888) );
  INV_X1 U2363 ( .A(n5889), .ZN(n12087) );
  AOI22_X1 U2364 ( .A1(ram[1415]), .A2(n5882), .B1(n12096), .B2(n9035), .ZN(
        n5889) );
  INV_X1 U2365 ( .A(n5890), .ZN(n12088) );
  AOI22_X1 U2366 ( .A1(ram[1416]), .A2(n5882), .B1(n12096), .B2(n9059), .ZN(
        n5890) );
  INV_X1 U2367 ( .A(n5891), .ZN(n12089) );
  AOI22_X1 U2368 ( .A1(ram[1417]), .A2(n5882), .B1(n12096), .B2(n9083), .ZN(
        n5891) );
  INV_X1 U2369 ( .A(n5892), .ZN(n12090) );
  AOI22_X1 U2370 ( .A1(ram[1418]), .A2(n5882), .B1(n12096), .B2(n9107), .ZN(
        n5892) );
  INV_X1 U2371 ( .A(n5893), .ZN(n12091) );
  AOI22_X1 U2372 ( .A1(ram[1419]), .A2(n5882), .B1(n12096), .B2(n9131), .ZN(
        n5893) );
  INV_X1 U2373 ( .A(n5894), .ZN(n12092) );
  AOI22_X1 U2374 ( .A1(ram[1420]), .A2(n5882), .B1(n12096), .B2(n9155), .ZN(
        n5894) );
  INV_X1 U2375 ( .A(n5895), .ZN(n12093) );
  AOI22_X1 U2376 ( .A1(ram[1421]), .A2(n5882), .B1(n12096), .B2(n9179), .ZN(
        n5895) );
  INV_X1 U2377 ( .A(n5896), .ZN(n12094) );
  AOI22_X1 U2378 ( .A1(ram[1422]), .A2(n5882), .B1(n12096), .B2(n9203), .ZN(
        n5896) );
  INV_X1 U2379 ( .A(n5897), .ZN(n12095) );
  AOI22_X1 U2380 ( .A1(ram[1423]), .A2(n5882), .B1(n12096), .B2(n9227), .ZN(
        n5897) );
  INV_X1 U2381 ( .A(n5915), .ZN(n12046) );
  AOI22_X1 U2382 ( .A1(ram[1440]), .A2(n5916), .B1(n12062), .B2(n8867), .ZN(
        n5915) );
  INV_X1 U2383 ( .A(n5917), .ZN(n12047) );
  AOI22_X1 U2384 ( .A1(ram[1441]), .A2(n5916), .B1(n12062), .B2(n8891), .ZN(
        n5917) );
  INV_X1 U2385 ( .A(n5918), .ZN(n12048) );
  AOI22_X1 U2386 ( .A1(ram[1442]), .A2(n5916), .B1(n12062), .B2(n8915), .ZN(
        n5918) );
  INV_X1 U2387 ( .A(n5919), .ZN(n12049) );
  AOI22_X1 U2388 ( .A1(ram[1443]), .A2(n5916), .B1(n12062), .B2(n8939), .ZN(
        n5919) );
  INV_X1 U2389 ( .A(n5920), .ZN(n12050) );
  AOI22_X1 U2390 ( .A1(ram[1444]), .A2(n5916), .B1(n12062), .B2(n8963), .ZN(
        n5920) );
  INV_X1 U2391 ( .A(n5921), .ZN(n12051) );
  AOI22_X1 U2392 ( .A1(ram[1445]), .A2(n5916), .B1(n12062), .B2(n8987), .ZN(
        n5921) );
  INV_X1 U2393 ( .A(n5922), .ZN(n12052) );
  AOI22_X1 U2394 ( .A1(ram[1446]), .A2(n5916), .B1(n12062), .B2(n9011), .ZN(
        n5922) );
  INV_X1 U2395 ( .A(n5923), .ZN(n12053) );
  AOI22_X1 U2396 ( .A1(ram[1447]), .A2(n5916), .B1(n12062), .B2(n9035), .ZN(
        n5923) );
  INV_X1 U2397 ( .A(n5924), .ZN(n12054) );
  AOI22_X1 U2398 ( .A1(ram[1448]), .A2(n5916), .B1(n12062), .B2(n9059), .ZN(
        n5924) );
  INV_X1 U2399 ( .A(n5925), .ZN(n12055) );
  AOI22_X1 U2400 ( .A1(ram[1449]), .A2(n5916), .B1(n12062), .B2(n9083), .ZN(
        n5925) );
  INV_X1 U2401 ( .A(n5926), .ZN(n12056) );
  AOI22_X1 U2402 ( .A1(ram[1450]), .A2(n5916), .B1(n12062), .B2(n9107), .ZN(
        n5926) );
  INV_X1 U2403 ( .A(n5927), .ZN(n12057) );
  AOI22_X1 U2404 ( .A1(ram[1451]), .A2(n5916), .B1(n12062), .B2(n9131), .ZN(
        n5927) );
  INV_X1 U2405 ( .A(n5928), .ZN(n12058) );
  AOI22_X1 U2406 ( .A1(ram[1452]), .A2(n5916), .B1(n12062), .B2(n9155), .ZN(
        n5928) );
  INV_X1 U2407 ( .A(n5929), .ZN(n12059) );
  AOI22_X1 U2408 ( .A1(ram[1453]), .A2(n5916), .B1(n12062), .B2(n9179), .ZN(
        n5929) );
  INV_X1 U2409 ( .A(n5930), .ZN(n12060) );
  AOI22_X1 U2410 ( .A1(ram[1454]), .A2(n5916), .B1(n12062), .B2(n9203), .ZN(
        n5930) );
  INV_X1 U2411 ( .A(n5931), .ZN(n12061) );
  AOI22_X1 U2412 ( .A1(ram[1455]), .A2(n5916), .B1(n12062), .B2(n9227), .ZN(
        n5931) );
  INV_X1 U2413 ( .A(n5949), .ZN(n12012) );
  AOI22_X1 U2414 ( .A1(ram[1472]), .A2(n5950), .B1(n12028), .B2(n8867), .ZN(
        n5949) );
  INV_X1 U2415 ( .A(n5951), .ZN(n12013) );
  AOI22_X1 U2416 ( .A1(ram[1473]), .A2(n5950), .B1(n12028), .B2(n8891), .ZN(
        n5951) );
  INV_X1 U2417 ( .A(n5952), .ZN(n12014) );
  AOI22_X1 U2418 ( .A1(ram[1474]), .A2(n5950), .B1(n12028), .B2(n8915), .ZN(
        n5952) );
  INV_X1 U2419 ( .A(n5953), .ZN(n12015) );
  AOI22_X1 U2420 ( .A1(ram[1475]), .A2(n5950), .B1(n12028), .B2(n8939), .ZN(
        n5953) );
  INV_X1 U2421 ( .A(n5954), .ZN(n12016) );
  AOI22_X1 U2422 ( .A1(ram[1476]), .A2(n5950), .B1(n12028), .B2(n8963), .ZN(
        n5954) );
  INV_X1 U2423 ( .A(n5955), .ZN(n12017) );
  AOI22_X1 U2424 ( .A1(ram[1477]), .A2(n5950), .B1(n12028), .B2(n8987), .ZN(
        n5955) );
  INV_X1 U2425 ( .A(n5956), .ZN(n12018) );
  AOI22_X1 U2426 ( .A1(ram[1478]), .A2(n5950), .B1(n12028), .B2(n9011), .ZN(
        n5956) );
  INV_X1 U2427 ( .A(n5957), .ZN(n12019) );
  AOI22_X1 U2428 ( .A1(ram[1479]), .A2(n5950), .B1(n12028), .B2(n9035), .ZN(
        n5957) );
  INV_X1 U2429 ( .A(n5958), .ZN(n12020) );
  AOI22_X1 U2430 ( .A1(ram[1480]), .A2(n5950), .B1(n12028), .B2(n9059), .ZN(
        n5958) );
  INV_X1 U2431 ( .A(n5959), .ZN(n12021) );
  AOI22_X1 U2432 ( .A1(ram[1481]), .A2(n5950), .B1(n12028), .B2(n9083), .ZN(
        n5959) );
  INV_X1 U2433 ( .A(n5960), .ZN(n12022) );
  AOI22_X1 U2434 ( .A1(ram[1482]), .A2(n5950), .B1(n12028), .B2(n9107), .ZN(
        n5960) );
  INV_X1 U2435 ( .A(n5961), .ZN(n12023) );
  AOI22_X1 U2436 ( .A1(ram[1483]), .A2(n5950), .B1(n12028), .B2(n9131), .ZN(
        n5961) );
  INV_X1 U2437 ( .A(n5962), .ZN(n12024) );
  AOI22_X1 U2438 ( .A1(ram[1484]), .A2(n5950), .B1(n12028), .B2(n9155), .ZN(
        n5962) );
  INV_X1 U2439 ( .A(n5963), .ZN(n12025) );
  AOI22_X1 U2440 ( .A1(ram[1485]), .A2(n5950), .B1(n12028), .B2(n9179), .ZN(
        n5963) );
  INV_X1 U2441 ( .A(n5964), .ZN(n12026) );
  AOI22_X1 U2442 ( .A1(ram[1486]), .A2(n5950), .B1(n12028), .B2(n9203), .ZN(
        n5964) );
  INV_X1 U2443 ( .A(n5965), .ZN(n12027) );
  AOI22_X1 U2444 ( .A1(ram[1487]), .A2(n5950), .B1(n12028), .B2(n9227), .ZN(
        n5965) );
  INV_X1 U2445 ( .A(n5983), .ZN(n11978) );
  AOI22_X1 U2446 ( .A1(ram[1504]), .A2(n5984), .B1(n11994), .B2(n8867), .ZN(
        n5983) );
  INV_X1 U2447 ( .A(n5985), .ZN(n11979) );
  AOI22_X1 U2448 ( .A1(ram[1505]), .A2(n5984), .B1(n11994), .B2(n8891), .ZN(
        n5985) );
  INV_X1 U2449 ( .A(n5986), .ZN(n11980) );
  AOI22_X1 U2450 ( .A1(ram[1506]), .A2(n5984), .B1(n11994), .B2(n8915), .ZN(
        n5986) );
  INV_X1 U2451 ( .A(n5987), .ZN(n11981) );
  AOI22_X1 U2452 ( .A1(ram[1507]), .A2(n5984), .B1(n11994), .B2(n8939), .ZN(
        n5987) );
  INV_X1 U2453 ( .A(n5988), .ZN(n11982) );
  AOI22_X1 U2454 ( .A1(ram[1508]), .A2(n5984), .B1(n11994), .B2(n8963), .ZN(
        n5988) );
  INV_X1 U2455 ( .A(n5989), .ZN(n11983) );
  AOI22_X1 U2456 ( .A1(ram[1509]), .A2(n5984), .B1(n11994), .B2(n8987), .ZN(
        n5989) );
  INV_X1 U2457 ( .A(n5990), .ZN(n11984) );
  AOI22_X1 U2458 ( .A1(ram[1510]), .A2(n5984), .B1(n11994), .B2(n9011), .ZN(
        n5990) );
  INV_X1 U2459 ( .A(n5991), .ZN(n11985) );
  AOI22_X1 U2460 ( .A1(ram[1511]), .A2(n5984), .B1(n11994), .B2(n9035), .ZN(
        n5991) );
  INV_X1 U2461 ( .A(n5992), .ZN(n11986) );
  AOI22_X1 U2462 ( .A1(ram[1512]), .A2(n5984), .B1(n11994), .B2(n9059), .ZN(
        n5992) );
  INV_X1 U2463 ( .A(n5993), .ZN(n11987) );
  AOI22_X1 U2464 ( .A1(ram[1513]), .A2(n5984), .B1(n11994), .B2(n9083), .ZN(
        n5993) );
  INV_X1 U2465 ( .A(n5994), .ZN(n11988) );
  AOI22_X1 U2466 ( .A1(ram[1514]), .A2(n5984), .B1(n11994), .B2(n9107), .ZN(
        n5994) );
  INV_X1 U2467 ( .A(n5995), .ZN(n11989) );
  AOI22_X1 U2468 ( .A1(ram[1515]), .A2(n5984), .B1(n11994), .B2(n9131), .ZN(
        n5995) );
  INV_X1 U2469 ( .A(n5996), .ZN(n11990) );
  AOI22_X1 U2470 ( .A1(ram[1516]), .A2(n5984), .B1(n11994), .B2(n9155), .ZN(
        n5996) );
  INV_X1 U2471 ( .A(n5997), .ZN(n11991) );
  AOI22_X1 U2472 ( .A1(ram[1517]), .A2(n5984), .B1(n11994), .B2(n9179), .ZN(
        n5997) );
  INV_X1 U2473 ( .A(n5998), .ZN(n11992) );
  AOI22_X1 U2474 ( .A1(ram[1518]), .A2(n5984), .B1(n11994), .B2(n9203), .ZN(
        n5998) );
  INV_X1 U2475 ( .A(n5999), .ZN(n11993) );
  AOI22_X1 U2476 ( .A1(ram[1519]), .A2(n5984), .B1(n11994), .B2(n9227), .ZN(
        n5999) );
  INV_X1 U2477 ( .A(n6017), .ZN(n11944) );
  AOI22_X1 U2478 ( .A1(ram[1536]), .A2(n6018), .B1(n11960), .B2(n8867), .ZN(
        n6017) );
  INV_X1 U2479 ( .A(n6019), .ZN(n11945) );
  AOI22_X1 U2480 ( .A1(ram[1537]), .A2(n6018), .B1(n11960), .B2(n8891), .ZN(
        n6019) );
  INV_X1 U2481 ( .A(n6020), .ZN(n11946) );
  AOI22_X1 U2482 ( .A1(ram[1538]), .A2(n6018), .B1(n11960), .B2(n8915), .ZN(
        n6020) );
  INV_X1 U2483 ( .A(n6021), .ZN(n11947) );
  AOI22_X1 U2484 ( .A1(ram[1539]), .A2(n6018), .B1(n11960), .B2(n8939), .ZN(
        n6021) );
  INV_X1 U2485 ( .A(n6022), .ZN(n11948) );
  AOI22_X1 U2486 ( .A1(ram[1540]), .A2(n6018), .B1(n11960), .B2(n8963), .ZN(
        n6022) );
  INV_X1 U2487 ( .A(n6023), .ZN(n11949) );
  AOI22_X1 U2488 ( .A1(ram[1541]), .A2(n6018), .B1(n11960), .B2(n8987), .ZN(
        n6023) );
  INV_X1 U2489 ( .A(n6024), .ZN(n11950) );
  AOI22_X1 U2490 ( .A1(ram[1542]), .A2(n6018), .B1(n11960), .B2(n9011), .ZN(
        n6024) );
  INV_X1 U2491 ( .A(n6025), .ZN(n11951) );
  AOI22_X1 U2492 ( .A1(ram[1543]), .A2(n6018), .B1(n11960), .B2(n9035), .ZN(
        n6025) );
  INV_X1 U2493 ( .A(n6026), .ZN(n11952) );
  AOI22_X1 U2494 ( .A1(ram[1544]), .A2(n6018), .B1(n11960), .B2(n9059), .ZN(
        n6026) );
  INV_X1 U2495 ( .A(n6027), .ZN(n11953) );
  AOI22_X1 U2496 ( .A1(ram[1545]), .A2(n6018), .B1(n11960), .B2(n9083), .ZN(
        n6027) );
  INV_X1 U2497 ( .A(n6028), .ZN(n11954) );
  AOI22_X1 U2498 ( .A1(ram[1546]), .A2(n6018), .B1(n11960), .B2(n9107), .ZN(
        n6028) );
  INV_X1 U2499 ( .A(n6029), .ZN(n11955) );
  AOI22_X1 U2500 ( .A1(ram[1547]), .A2(n6018), .B1(n11960), .B2(n9131), .ZN(
        n6029) );
  INV_X1 U2501 ( .A(n6030), .ZN(n11956) );
  AOI22_X1 U2502 ( .A1(ram[1548]), .A2(n6018), .B1(n11960), .B2(n9155), .ZN(
        n6030) );
  INV_X1 U2503 ( .A(n6031), .ZN(n11957) );
  AOI22_X1 U2504 ( .A1(ram[1549]), .A2(n6018), .B1(n11960), .B2(n9179), .ZN(
        n6031) );
  INV_X1 U2505 ( .A(n6032), .ZN(n11958) );
  AOI22_X1 U2506 ( .A1(ram[1550]), .A2(n6018), .B1(n11960), .B2(n9203), .ZN(
        n6032) );
  INV_X1 U2507 ( .A(n6033), .ZN(n11959) );
  AOI22_X1 U2508 ( .A1(ram[1551]), .A2(n6018), .B1(n11960), .B2(n9227), .ZN(
        n6033) );
  INV_X1 U2509 ( .A(n6052), .ZN(n11910) );
  AOI22_X1 U2510 ( .A1(ram[1568]), .A2(n6053), .B1(n11926), .B2(n8867), .ZN(
        n6052) );
  INV_X1 U2511 ( .A(n6054), .ZN(n11911) );
  AOI22_X1 U2512 ( .A1(ram[1569]), .A2(n6053), .B1(n11926), .B2(n8891), .ZN(
        n6054) );
  INV_X1 U2513 ( .A(n6055), .ZN(n11912) );
  AOI22_X1 U2514 ( .A1(ram[1570]), .A2(n6053), .B1(n11926), .B2(n8915), .ZN(
        n6055) );
  INV_X1 U2515 ( .A(n6056), .ZN(n11913) );
  AOI22_X1 U2516 ( .A1(ram[1571]), .A2(n6053), .B1(n11926), .B2(n8939), .ZN(
        n6056) );
  INV_X1 U2517 ( .A(n6057), .ZN(n11914) );
  AOI22_X1 U2518 ( .A1(ram[1572]), .A2(n6053), .B1(n11926), .B2(n8963), .ZN(
        n6057) );
  INV_X1 U2519 ( .A(n6058), .ZN(n11915) );
  AOI22_X1 U2520 ( .A1(ram[1573]), .A2(n6053), .B1(n11926), .B2(n8987), .ZN(
        n6058) );
  INV_X1 U2521 ( .A(n6059), .ZN(n11916) );
  AOI22_X1 U2522 ( .A1(ram[1574]), .A2(n6053), .B1(n11926), .B2(n9011), .ZN(
        n6059) );
  INV_X1 U2523 ( .A(n6060), .ZN(n11917) );
  AOI22_X1 U2524 ( .A1(ram[1575]), .A2(n6053), .B1(n11926), .B2(n9035), .ZN(
        n6060) );
  INV_X1 U2525 ( .A(n6061), .ZN(n11918) );
  AOI22_X1 U2526 ( .A1(ram[1576]), .A2(n6053), .B1(n11926), .B2(n9059), .ZN(
        n6061) );
  INV_X1 U2527 ( .A(n6062), .ZN(n11919) );
  AOI22_X1 U2528 ( .A1(ram[1577]), .A2(n6053), .B1(n11926), .B2(n9083), .ZN(
        n6062) );
  INV_X1 U2529 ( .A(n6063), .ZN(n11920) );
  AOI22_X1 U2530 ( .A1(ram[1578]), .A2(n6053), .B1(n11926), .B2(n9107), .ZN(
        n6063) );
  INV_X1 U2531 ( .A(n6064), .ZN(n11921) );
  AOI22_X1 U2532 ( .A1(ram[1579]), .A2(n6053), .B1(n11926), .B2(n9131), .ZN(
        n6064) );
  INV_X1 U2533 ( .A(n6065), .ZN(n11922) );
  AOI22_X1 U2534 ( .A1(ram[1580]), .A2(n6053), .B1(n11926), .B2(n9155), .ZN(
        n6065) );
  INV_X1 U2535 ( .A(n6066), .ZN(n11923) );
  AOI22_X1 U2536 ( .A1(ram[1581]), .A2(n6053), .B1(n11926), .B2(n9179), .ZN(
        n6066) );
  INV_X1 U2537 ( .A(n6067), .ZN(n11924) );
  AOI22_X1 U2538 ( .A1(ram[1582]), .A2(n6053), .B1(n11926), .B2(n9203), .ZN(
        n6067) );
  INV_X1 U2539 ( .A(n6068), .ZN(n11925) );
  AOI22_X1 U2540 ( .A1(ram[1583]), .A2(n6053), .B1(n11926), .B2(n9227), .ZN(
        n6068) );
  INV_X1 U2541 ( .A(n6086), .ZN(n11876) );
  AOI22_X1 U2542 ( .A1(ram[1600]), .A2(n6087), .B1(n11892), .B2(n8866), .ZN(
        n6086) );
  INV_X1 U2543 ( .A(n6088), .ZN(n11877) );
  AOI22_X1 U2544 ( .A1(ram[1601]), .A2(n6087), .B1(n11892), .B2(n8890), .ZN(
        n6088) );
  INV_X1 U2545 ( .A(n6089), .ZN(n11878) );
  AOI22_X1 U2546 ( .A1(ram[1602]), .A2(n6087), .B1(n11892), .B2(n8914), .ZN(
        n6089) );
  INV_X1 U2547 ( .A(n6090), .ZN(n11879) );
  AOI22_X1 U2548 ( .A1(ram[1603]), .A2(n6087), .B1(n11892), .B2(n8938), .ZN(
        n6090) );
  INV_X1 U2549 ( .A(n6091), .ZN(n11880) );
  AOI22_X1 U2550 ( .A1(ram[1604]), .A2(n6087), .B1(n11892), .B2(n8962), .ZN(
        n6091) );
  INV_X1 U2551 ( .A(n6092), .ZN(n11881) );
  AOI22_X1 U2552 ( .A1(ram[1605]), .A2(n6087), .B1(n11892), .B2(n8986), .ZN(
        n6092) );
  INV_X1 U2553 ( .A(n6093), .ZN(n11882) );
  AOI22_X1 U2554 ( .A1(ram[1606]), .A2(n6087), .B1(n11892), .B2(n9010), .ZN(
        n6093) );
  INV_X1 U2555 ( .A(n6094), .ZN(n11883) );
  AOI22_X1 U2556 ( .A1(ram[1607]), .A2(n6087), .B1(n11892), .B2(n9034), .ZN(
        n6094) );
  INV_X1 U2557 ( .A(n6095), .ZN(n11884) );
  AOI22_X1 U2558 ( .A1(ram[1608]), .A2(n6087), .B1(n11892), .B2(n9058), .ZN(
        n6095) );
  INV_X1 U2559 ( .A(n6096), .ZN(n11885) );
  AOI22_X1 U2560 ( .A1(ram[1609]), .A2(n6087), .B1(n11892), .B2(n9082), .ZN(
        n6096) );
  INV_X1 U2561 ( .A(n6097), .ZN(n11886) );
  AOI22_X1 U2562 ( .A1(ram[1610]), .A2(n6087), .B1(n11892), .B2(n9106), .ZN(
        n6097) );
  INV_X1 U2563 ( .A(n6098), .ZN(n11887) );
  AOI22_X1 U2564 ( .A1(ram[1611]), .A2(n6087), .B1(n11892), .B2(n9130), .ZN(
        n6098) );
  INV_X1 U2565 ( .A(n6099), .ZN(n11888) );
  AOI22_X1 U2566 ( .A1(ram[1612]), .A2(n6087), .B1(n11892), .B2(n9154), .ZN(
        n6099) );
  INV_X1 U2567 ( .A(n6100), .ZN(n11889) );
  AOI22_X1 U2568 ( .A1(ram[1613]), .A2(n6087), .B1(n11892), .B2(n9178), .ZN(
        n6100) );
  INV_X1 U2569 ( .A(n6101), .ZN(n11890) );
  AOI22_X1 U2570 ( .A1(ram[1614]), .A2(n6087), .B1(n11892), .B2(n9202), .ZN(
        n6101) );
  INV_X1 U2571 ( .A(n6102), .ZN(n11891) );
  AOI22_X1 U2572 ( .A1(ram[1615]), .A2(n6087), .B1(n11892), .B2(n9226), .ZN(
        n6102) );
  INV_X1 U2573 ( .A(n6120), .ZN(n11842) );
  AOI22_X1 U2574 ( .A1(ram[1632]), .A2(n6121), .B1(n11858), .B2(n8866), .ZN(
        n6120) );
  INV_X1 U2575 ( .A(n6122), .ZN(n11843) );
  AOI22_X1 U2576 ( .A1(ram[1633]), .A2(n6121), .B1(n11858), .B2(n8890), .ZN(
        n6122) );
  INV_X1 U2577 ( .A(n6123), .ZN(n11844) );
  AOI22_X1 U2578 ( .A1(ram[1634]), .A2(n6121), .B1(n11858), .B2(n8914), .ZN(
        n6123) );
  INV_X1 U2579 ( .A(n6124), .ZN(n11845) );
  AOI22_X1 U2580 ( .A1(ram[1635]), .A2(n6121), .B1(n11858), .B2(n8938), .ZN(
        n6124) );
  INV_X1 U2581 ( .A(n6125), .ZN(n11846) );
  AOI22_X1 U2582 ( .A1(ram[1636]), .A2(n6121), .B1(n11858), .B2(n8962), .ZN(
        n6125) );
  INV_X1 U2583 ( .A(n6126), .ZN(n11847) );
  AOI22_X1 U2584 ( .A1(ram[1637]), .A2(n6121), .B1(n11858), .B2(n8986), .ZN(
        n6126) );
  INV_X1 U2585 ( .A(n6127), .ZN(n11848) );
  AOI22_X1 U2586 ( .A1(ram[1638]), .A2(n6121), .B1(n11858), .B2(n9010), .ZN(
        n6127) );
  INV_X1 U2587 ( .A(n6128), .ZN(n11849) );
  AOI22_X1 U2588 ( .A1(ram[1639]), .A2(n6121), .B1(n11858), .B2(n9034), .ZN(
        n6128) );
  INV_X1 U2589 ( .A(n6129), .ZN(n11850) );
  AOI22_X1 U2590 ( .A1(ram[1640]), .A2(n6121), .B1(n11858), .B2(n9058), .ZN(
        n6129) );
  INV_X1 U2591 ( .A(n6130), .ZN(n11851) );
  AOI22_X1 U2592 ( .A1(ram[1641]), .A2(n6121), .B1(n11858), .B2(n9082), .ZN(
        n6130) );
  INV_X1 U2593 ( .A(n6131), .ZN(n11852) );
  AOI22_X1 U2594 ( .A1(ram[1642]), .A2(n6121), .B1(n11858), .B2(n9106), .ZN(
        n6131) );
  INV_X1 U2595 ( .A(n6132), .ZN(n11853) );
  AOI22_X1 U2596 ( .A1(ram[1643]), .A2(n6121), .B1(n11858), .B2(n9130), .ZN(
        n6132) );
  INV_X1 U2597 ( .A(n6133), .ZN(n11854) );
  AOI22_X1 U2598 ( .A1(ram[1644]), .A2(n6121), .B1(n11858), .B2(n9154), .ZN(
        n6133) );
  INV_X1 U2599 ( .A(n6134), .ZN(n11855) );
  AOI22_X1 U2600 ( .A1(ram[1645]), .A2(n6121), .B1(n11858), .B2(n9178), .ZN(
        n6134) );
  INV_X1 U2601 ( .A(n6135), .ZN(n11856) );
  AOI22_X1 U2602 ( .A1(ram[1646]), .A2(n6121), .B1(n11858), .B2(n9202), .ZN(
        n6135) );
  INV_X1 U2603 ( .A(n6136), .ZN(n11857) );
  AOI22_X1 U2604 ( .A1(ram[1647]), .A2(n6121), .B1(n11858), .B2(n9226), .ZN(
        n6136) );
  INV_X1 U2605 ( .A(n6154), .ZN(n11808) );
  AOI22_X1 U2606 ( .A1(ram[1664]), .A2(n6155), .B1(n11824), .B2(n8866), .ZN(
        n6154) );
  INV_X1 U2607 ( .A(n6156), .ZN(n11809) );
  AOI22_X1 U2608 ( .A1(ram[1665]), .A2(n6155), .B1(n11824), .B2(n8890), .ZN(
        n6156) );
  INV_X1 U2609 ( .A(n6157), .ZN(n11810) );
  AOI22_X1 U2610 ( .A1(ram[1666]), .A2(n6155), .B1(n11824), .B2(n8914), .ZN(
        n6157) );
  INV_X1 U2611 ( .A(n6158), .ZN(n11811) );
  AOI22_X1 U2612 ( .A1(ram[1667]), .A2(n6155), .B1(n11824), .B2(n8938), .ZN(
        n6158) );
  INV_X1 U2613 ( .A(n6159), .ZN(n11812) );
  AOI22_X1 U2614 ( .A1(ram[1668]), .A2(n6155), .B1(n11824), .B2(n8962), .ZN(
        n6159) );
  INV_X1 U2615 ( .A(n6160), .ZN(n11813) );
  AOI22_X1 U2616 ( .A1(ram[1669]), .A2(n6155), .B1(n11824), .B2(n8986), .ZN(
        n6160) );
  INV_X1 U2617 ( .A(n6161), .ZN(n11814) );
  AOI22_X1 U2618 ( .A1(ram[1670]), .A2(n6155), .B1(n11824), .B2(n9010), .ZN(
        n6161) );
  INV_X1 U2619 ( .A(n6162), .ZN(n11815) );
  AOI22_X1 U2620 ( .A1(ram[1671]), .A2(n6155), .B1(n11824), .B2(n9034), .ZN(
        n6162) );
  INV_X1 U2621 ( .A(n6163), .ZN(n11816) );
  AOI22_X1 U2622 ( .A1(ram[1672]), .A2(n6155), .B1(n11824), .B2(n9058), .ZN(
        n6163) );
  INV_X1 U2623 ( .A(n6164), .ZN(n11817) );
  AOI22_X1 U2624 ( .A1(ram[1673]), .A2(n6155), .B1(n11824), .B2(n9082), .ZN(
        n6164) );
  INV_X1 U2625 ( .A(n6165), .ZN(n11818) );
  AOI22_X1 U2626 ( .A1(ram[1674]), .A2(n6155), .B1(n11824), .B2(n9106), .ZN(
        n6165) );
  INV_X1 U2627 ( .A(n6166), .ZN(n11819) );
  AOI22_X1 U2628 ( .A1(ram[1675]), .A2(n6155), .B1(n11824), .B2(n9130), .ZN(
        n6166) );
  INV_X1 U2629 ( .A(n6167), .ZN(n11820) );
  AOI22_X1 U2630 ( .A1(ram[1676]), .A2(n6155), .B1(n11824), .B2(n9154), .ZN(
        n6167) );
  INV_X1 U2631 ( .A(n6168), .ZN(n11821) );
  AOI22_X1 U2632 ( .A1(ram[1677]), .A2(n6155), .B1(n11824), .B2(n9178), .ZN(
        n6168) );
  INV_X1 U2633 ( .A(n6169), .ZN(n11822) );
  AOI22_X1 U2634 ( .A1(ram[1678]), .A2(n6155), .B1(n11824), .B2(n9202), .ZN(
        n6169) );
  INV_X1 U2635 ( .A(n6170), .ZN(n11823) );
  AOI22_X1 U2636 ( .A1(ram[1679]), .A2(n6155), .B1(n11824), .B2(n9226), .ZN(
        n6170) );
  INV_X1 U2637 ( .A(n6188), .ZN(n11774) );
  AOI22_X1 U2638 ( .A1(ram[1696]), .A2(n6189), .B1(n11790), .B2(n8866), .ZN(
        n6188) );
  INV_X1 U2639 ( .A(n6190), .ZN(n11775) );
  AOI22_X1 U2640 ( .A1(ram[1697]), .A2(n6189), .B1(n11790), .B2(n8890), .ZN(
        n6190) );
  INV_X1 U2641 ( .A(n6191), .ZN(n11776) );
  AOI22_X1 U2642 ( .A1(ram[1698]), .A2(n6189), .B1(n11790), .B2(n8914), .ZN(
        n6191) );
  INV_X1 U2643 ( .A(n6192), .ZN(n11777) );
  AOI22_X1 U2644 ( .A1(ram[1699]), .A2(n6189), .B1(n11790), .B2(n8938), .ZN(
        n6192) );
  INV_X1 U2645 ( .A(n6193), .ZN(n11778) );
  AOI22_X1 U2646 ( .A1(ram[1700]), .A2(n6189), .B1(n11790), .B2(n8962), .ZN(
        n6193) );
  INV_X1 U2647 ( .A(n6194), .ZN(n11779) );
  AOI22_X1 U2648 ( .A1(ram[1701]), .A2(n6189), .B1(n11790), .B2(n8986), .ZN(
        n6194) );
  INV_X1 U2649 ( .A(n6195), .ZN(n11780) );
  AOI22_X1 U2650 ( .A1(ram[1702]), .A2(n6189), .B1(n11790), .B2(n9010), .ZN(
        n6195) );
  INV_X1 U2651 ( .A(n6196), .ZN(n11781) );
  AOI22_X1 U2652 ( .A1(ram[1703]), .A2(n6189), .B1(n11790), .B2(n9034), .ZN(
        n6196) );
  INV_X1 U2653 ( .A(n6197), .ZN(n11782) );
  AOI22_X1 U2654 ( .A1(ram[1704]), .A2(n6189), .B1(n11790), .B2(n9058), .ZN(
        n6197) );
  INV_X1 U2655 ( .A(n6198), .ZN(n11783) );
  AOI22_X1 U2656 ( .A1(ram[1705]), .A2(n6189), .B1(n11790), .B2(n9082), .ZN(
        n6198) );
  INV_X1 U2657 ( .A(n6199), .ZN(n11784) );
  AOI22_X1 U2658 ( .A1(ram[1706]), .A2(n6189), .B1(n11790), .B2(n9106), .ZN(
        n6199) );
  INV_X1 U2659 ( .A(n6200), .ZN(n11785) );
  AOI22_X1 U2660 ( .A1(ram[1707]), .A2(n6189), .B1(n11790), .B2(n9130), .ZN(
        n6200) );
  INV_X1 U2661 ( .A(n6201), .ZN(n11786) );
  AOI22_X1 U2662 ( .A1(ram[1708]), .A2(n6189), .B1(n11790), .B2(n9154), .ZN(
        n6201) );
  INV_X1 U2663 ( .A(n6202), .ZN(n11787) );
  AOI22_X1 U2664 ( .A1(ram[1709]), .A2(n6189), .B1(n11790), .B2(n9178), .ZN(
        n6202) );
  INV_X1 U2665 ( .A(n6203), .ZN(n11788) );
  AOI22_X1 U2666 ( .A1(ram[1710]), .A2(n6189), .B1(n11790), .B2(n9202), .ZN(
        n6203) );
  INV_X1 U2667 ( .A(n6204), .ZN(n11789) );
  AOI22_X1 U2668 ( .A1(ram[1711]), .A2(n6189), .B1(n11790), .B2(n9226), .ZN(
        n6204) );
  INV_X1 U2669 ( .A(n6222), .ZN(n11740) );
  AOI22_X1 U2670 ( .A1(ram[1728]), .A2(n6223), .B1(n11756), .B2(n8866), .ZN(
        n6222) );
  INV_X1 U2671 ( .A(n6224), .ZN(n11741) );
  AOI22_X1 U2672 ( .A1(ram[1729]), .A2(n6223), .B1(n11756), .B2(n8890), .ZN(
        n6224) );
  INV_X1 U2673 ( .A(n6225), .ZN(n11742) );
  AOI22_X1 U2674 ( .A1(ram[1730]), .A2(n6223), .B1(n11756), .B2(n8914), .ZN(
        n6225) );
  INV_X1 U2675 ( .A(n6226), .ZN(n11743) );
  AOI22_X1 U2676 ( .A1(ram[1731]), .A2(n6223), .B1(n11756), .B2(n8938), .ZN(
        n6226) );
  INV_X1 U2677 ( .A(n6227), .ZN(n11744) );
  AOI22_X1 U2678 ( .A1(ram[1732]), .A2(n6223), .B1(n11756), .B2(n8962), .ZN(
        n6227) );
  INV_X1 U2679 ( .A(n6228), .ZN(n11745) );
  AOI22_X1 U2680 ( .A1(ram[1733]), .A2(n6223), .B1(n11756), .B2(n8986), .ZN(
        n6228) );
  INV_X1 U2681 ( .A(n6229), .ZN(n11746) );
  AOI22_X1 U2682 ( .A1(ram[1734]), .A2(n6223), .B1(n11756), .B2(n9010), .ZN(
        n6229) );
  INV_X1 U2683 ( .A(n6230), .ZN(n11747) );
  AOI22_X1 U2684 ( .A1(ram[1735]), .A2(n6223), .B1(n11756), .B2(n9034), .ZN(
        n6230) );
  INV_X1 U2685 ( .A(n6231), .ZN(n11748) );
  AOI22_X1 U2686 ( .A1(ram[1736]), .A2(n6223), .B1(n11756), .B2(n9058), .ZN(
        n6231) );
  INV_X1 U2687 ( .A(n6232), .ZN(n11749) );
  AOI22_X1 U2688 ( .A1(ram[1737]), .A2(n6223), .B1(n11756), .B2(n9082), .ZN(
        n6232) );
  INV_X1 U2689 ( .A(n6233), .ZN(n11750) );
  AOI22_X1 U2690 ( .A1(ram[1738]), .A2(n6223), .B1(n11756), .B2(n9106), .ZN(
        n6233) );
  INV_X1 U2691 ( .A(n6234), .ZN(n11751) );
  AOI22_X1 U2692 ( .A1(ram[1739]), .A2(n6223), .B1(n11756), .B2(n9130), .ZN(
        n6234) );
  INV_X1 U2693 ( .A(n6235), .ZN(n11752) );
  AOI22_X1 U2694 ( .A1(ram[1740]), .A2(n6223), .B1(n11756), .B2(n9154), .ZN(
        n6235) );
  INV_X1 U2695 ( .A(n6236), .ZN(n11753) );
  AOI22_X1 U2696 ( .A1(ram[1741]), .A2(n6223), .B1(n11756), .B2(n9178), .ZN(
        n6236) );
  INV_X1 U2697 ( .A(n6237), .ZN(n11754) );
  AOI22_X1 U2698 ( .A1(ram[1742]), .A2(n6223), .B1(n11756), .B2(n9202), .ZN(
        n6237) );
  INV_X1 U2699 ( .A(n6238), .ZN(n11755) );
  AOI22_X1 U2700 ( .A1(ram[1743]), .A2(n6223), .B1(n11756), .B2(n9226), .ZN(
        n6238) );
  INV_X1 U2701 ( .A(n6256), .ZN(n11706) );
  AOI22_X1 U2702 ( .A1(ram[1760]), .A2(n6257), .B1(n11722), .B2(n8866), .ZN(
        n6256) );
  INV_X1 U2703 ( .A(n6258), .ZN(n11707) );
  AOI22_X1 U2704 ( .A1(ram[1761]), .A2(n6257), .B1(n11722), .B2(n8890), .ZN(
        n6258) );
  INV_X1 U2705 ( .A(n6259), .ZN(n11708) );
  AOI22_X1 U2706 ( .A1(ram[1762]), .A2(n6257), .B1(n11722), .B2(n8914), .ZN(
        n6259) );
  INV_X1 U2707 ( .A(n6260), .ZN(n11709) );
  AOI22_X1 U2708 ( .A1(ram[1763]), .A2(n6257), .B1(n11722), .B2(n8938), .ZN(
        n6260) );
  INV_X1 U2709 ( .A(n6261), .ZN(n11710) );
  AOI22_X1 U2710 ( .A1(ram[1764]), .A2(n6257), .B1(n11722), .B2(n8962), .ZN(
        n6261) );
  INV_X1 U2711 ( .A(n6262), .ZN(n11711) );
  AOI22_X1 U2712 ( .A1(ram[1765]), .A2(n6257), .B1(n11722), .B2(n8986), .ZN(
        n6262) );
  INV_X1 U2713 ( .A(n6263), .ZN(n11712) );
  AOI22_X1 U2714 ( .A1(ram[1766]), .A2(n6257), .B1(n11722), .B2(n9010), .ZN(
        n6263) );
  INV_X1 U2715 ( .A(n6264), .ZN(n11713) );
  AOI22_X1 U2716 ( .A1(ram[1767]), .A2(n6257), .B1(n11722), .B2(n9034), .ZN(
        n6264) );
  INV_X1 U2717 ( .A(n6265), .ZN(n11714) );
  AOI22_X1 U2718 ( .A1(ram[1768]), .A2(n6257), .B1(n11722), .B2(n9058), .ZN(
        n6265) );
  INV_X1 U2719 ( .A(n6266), .ZN(n11715) );
  AOI22_X1 U2720 ( .A1(ram[1769]), .A2(n6257), .B1(n11722), .B2(n9082), .ZN(
        n6266) );
  INV_X1 U2721 ( .A(n6267), .ZN(n11716) );
  AOI22_X1 U2722 ( .A1(ram[1770]), .A2(n6257), .B1(n11722), .B2(n9106), .ZN(
        n6267) );
  INV_X1 U2723 ( .A(n6268), .ZN(n11717) );
  AOI22_X1 U2724 ( .A1(ram[1771]), .A2(n6257), .B1(n11722), .B2(n9130), .ZN(
        n6268) );
  INV_X1 U2725 ( .A(n6269), .ZN(n11718) );
  AOI22_X1 U2726 ( .A1(ram[1772]), .A2(n6257), .B1(n11722), .B2(n9154), .ZN(
        n6269) );
  INV_X1 U2727 ( .A(n6270), .ZN(n11719) );
  AOI22_X1 U2728 ( .A1(ram[1773]), .A2(n6257), .B1(n11722), .B2(n9178), .ZN(
        n6270) );
  INV_X1 U2729 ( .A(n6271), .ZN(n11720) );
  AOI22_X1 U2730 ( .A1(ram[1774]), .A2(n6257), .B1(n11722), .B2(n9202), .ZN(
        n6271) );
  INV_X1 U2731 ( .A(n6272), .ZN(n11721) );
  AOI22_X1 U2732 ( .A1(ram[1775]), .A2(n6257), .B1(n11722), .B2(n9226), .ZN(
        n6272) );
  INV_X1 U2733 ( .A(n6290), .ZN(n11672) );
  AOI22_X1 U2734 ( .A1(ram[1792]), .A2(n6291), .B1(n11688), .B2(n8865), .ZN(
        n6290) );
  INV_X1 U2735 ( .A(n6292), .ZN(n11673) );
  AOI22_X1 U2736 ( .A1(ram[1793]), .A2(n6291), .B1(n11688), .B2(n8889), .ZN(
        n6292) );
  INV_X1 U2737 ( .A(n6293), .ZN(n11674) );
  AOI22_X1 U2738 ( .A1(ram[1794]), .A2(n6291), .B1(n11688), .B2(n8913), .ZN(
        n6293) );
  INV_X1 U2739 ( .A(n6294), .ZN(n11675) );
  AOI22_X1 U2740 ( .A1(ram[1795]), .A2(n6291), .B1(n11688), .B2(n8937), .ZN(
        n6294) );
  INV_X1 U2741 ( .A(n6295), .ZN(n11676) );
  AOI22_X1 U2742 ( .A1(ram[1796]), .A2(n6291), .B1(n11688), .B2(n8961), .ZN(
        n6295) );
  INV_X1 U2743 ( .A(n6296), .ZN(n11677) );
  AOI22_X1 U2744 ( .A1(ram[1797]), .A2(n6291), .B1(n11688), .B2(n8985), .ZN(
        n6296) );
  INV_X1 U2745 ( .A(n6297), .ZN(n11678) );
  AOI22_X1 U2746 ( .A1(ram[1798]), .A2(n6291), .B1(n11688), .B2(n9009), .ZN(
        n6297) );
  INV_X1 U2747 ( .A(n6298), .ZN(n11679) );
  AOI22_X1 U2748 ( .A1(ram[1799]), .A2(n6291), .B1(n11688), .B2(n9033), .ZN(
        n6298) );
  INV_X1 U2749 ( .A(n6299), .ZN(n11680) );
  AOI22_X1 U2750 ( .A1(ram[1800]), .A2(n6291), .B1(n11688), .B2(n9057), .ZN(
        n6299) );
  INV_X1 U2751 ( .A(n6300), .ZN(n11681) );
  AOI22_X1 U2752 ( .A1(ram[1801]), .A2(n6291), .B1(n11688), .B2(n9081), .ZN(
        n6300) );
  INV_X1 U2753 ( .A(n6301), .ZN(n11682) );
  AOI22_X1 U2754 ( .A1(ram[1802]), .A2(n6291), .B1(n11688), .B2(n9105), .ZN(
        n6301) );
  INV_X1 U2755 ( .A(n6302), .ZN(n11683) );
  AOI22_X1 U2756 ( .A1(ram[1803]), .A2(n6291), .B1(n11688), .B2(n9129), .ZN(
        n6302) );
  INV_X1 U2757 ( .A(n6303), .ZN(n11684) );
  AOI22_X1 U2758 ( .A1(ram[1804]), .A2(n6291), .B1(n11688), .B2(n9153), .ZN(
        n6303) );
  INV_X1 U2759 ( .A(n6304), .ZN(n11685) );
  AOI22_X1 U2760 ( .A1(ram[1805]), .A2(n6291), .B1(n11688), .B2(n9177), .ZN(
        n6304) );
  INV_X1 U2761 ( .A(n6305), .ZN(n11686) );
  AOI22_X1 U2762 ( .A1(ram[1806]), .A2(n6291), .B1(n11688), .B2(n9201), .ZN(
        n6305) );
  INV_X1 U2763 ( .A(n6306), .ZN(n11687) );
  AOI22_X1 U2764 ( .A1(ram[1807]), .A2(n6291), .B1(n11688), .B2(n9225), .ZN(
        n6306) );
  INV_X1 U2765 ( .A(n6325), .ZN(n11638) );
  AOI22_X1 U2766 ( .A1(ram[1824]), .A2(n6326), .B1(n11654), .B2(n8865), .ZN(
        n6325) );
  INV_X1 U2767 ( .A(n6327), .ZN(n11639) );
  AOI22_X1 U2768 ( .A1(ram[1825]), .A2(n6326), .B1(n11654), .B2(n8889), .ZN(
        n6327) );
  INV_X1 U2769 ( .A(n6328), .ZN(n11640) );
  AOI22_X1 U2770 ( .A1(ram[1826]), .A2(n6326), .B1(n11654), .B2(n8913), .ZN(
        n6328) );
  INV_X1 U2771 ( .A(n6329), .ZN(n11641) );
  AOI22_X1 U2772 ( .A1(ram[1827]), .A2(n6326), .B1(n11654), .B2(n8937), .ZN(
        n6329) );
  INV_X1 U2773 ( .A(n6330), .ZN(n11642) );
  AOI22_X1 U2774 ( .A1(ram[1828]), .A2(n6326), .B1(n11654), .B2(n8961), .ZN(
        n6330) );
  INV_X1 U2775 ( .A(n6331), .ZN(n11643) );
  AOI22_X1 U2776 ( .A1(ram[1829]), .A2(n6326), .B1(n11654), .B2(n8985), .ZN(
        n6331) );
  INV_X1 U2777 ( .A(n6332), .ZN(n11644) );
  AOI22_X1 U2778 ( .A1(ram[1830]), .A2(n6326), .B1(n11654), .B2(n9009), .ZN(
        n6332) );
  INV_X1 U2779 ( .A(n6333), .ZN(n11645) );
  AOI22_X1 U2780 ( .A1(ram[1831]), .A2(n6326), .B1(n11654), .B2(n9033), .ZN(
        n6333) );
  INV_X1 U2781 ( .A(n6334), .ZN(n11646) );
  AOI22_X1 U2782 ( .A1(ram[1832]), .A2(n6326), .B1(n11654), .B2(n9057), .ZN(
        n6334) );
  INV_X1 U2783 ( .A(n6335), .ZN(n11647) );
  AOI22_X1 U2784 ( .A1(ram[1833]), .A2(n6326), .B1(n11654), .B2(n9081), .ZN(
        n6335) );
  INV_X1 U2785 ( .A(n6336), .ZN(n11648) );
  AOI22_X1 U2786 ( .A1(ram[1834]), .A2(n6326), .B1(n11654), .B2(n9105), .ZN(
        n6336) );
  INV_X1 U2787 ( .A(n6337), .ZN(n11649) );
  AOI22_X1 U2788 ( .A1(ram[1835]), .A2(n6326), .B1(n11654), .B2(n9129), .ZN(
        n6337) );
  INV_X1 U2789 ( .A(n6338), .ZN(n11650) );
  AOI22_X1 U2790 ( .A1(ram[1836]), .A2(n6326), .B1(n11654), .B2(n9153), .ZN(
        n6338) );
  INV_X1 U2791 ( .A(n6339), .ZN(n11651) );
  AOI22_X1 U2792 ( .A1(ram[1837]), .A2(n6326), .B1(n11654), .B2(n9177), .ZN(
        n6339) );
  INV_X1 U2793 ( .A(n6340), .ZN(n11652) );
  AOI22_X1 U2794 ( .A1(ram[1838]), .A2(n6326), .B1(n11654), .B2(n9201), .ZN(
        n6340) );
  INV_X1 U2795 ( .A(n6341), .ZN(n11653) );
  AOI22_X1 U2796 ( .A1(ram[1839]), .A2(n6326), .B1(n11654), .B2(n9225), .ZN(
        n6341) );
  INV_X1 U2797 ( .A(n6359), .ZN(n11604) );
  AOI22_X1 U2798 ( .A1(ram[1856]), .A2(n6360), .B1(n11620), .B2(n8865), .ZN(
        n6359) );
  INV_X1 U2799 ( .A(n6361), .ZN(n11605) );
  AOI22_X1 U2800 ( .A1(ram[1857]), .A2(n6360), .B1(n11620), .B2(n8889), .ZN(
        n6361) );
  INV_X1 U2801 ( .A(n6362), .ZN(n11606) );
  AOI22_X1 U2802 ( .A1(ram[1858]), .A2(n6360), .B1(n11620), .B2(n8913), .ZN(
        n6362) );
  INV_X1 U2803 ( .A(n6363), .ZN(n11607) );
  AOI22_X1 U2804 ( .A1(ram[1859]), .A2(n6360), .B1(n11620), .B2(n8937), .ZN(
        n6363) );
  INV_X1 U2805 ( .A(n6364), .ZN(n11608) );
  AOI22_X1 U2806 ( .A1(ram[1860]), .A2(n6360), .B1(n11620), .B2(n8961), .ZN(
        n6364) );
  INV_X1 U2807 ( .A(n6365), .ZN(n11609) );
  AOI22_X1 U2808 ( .A1(ram[1861]), .A2(n6360), .B1(n11620), .B2(n8985), .ZN(
        n6365) );
  INV_X1 U2809 ( .A(n6366), .ZN(n11610) );
  AOI22_X1 U2810 ( .A1(ram[1862]), .A2(n6360), .B1(n11620), .B2(n9009), .ZN(
        n6366) );
  INV_X1 U2811 ( .A(n6367), .ZN(n11611) );
  AOI22_X1 U2812 ( .A1(ram[1863]), .A2(n6360), .B1(n11620), .B2(n9033), .ZN(
        n6367) );
  INV_X1 U2813 ( .A(n6368), .ZN(n11612) );
  AOI22_X1 U2814 ( .A1(ram[1864]), .A2(n6360), .B1(n11620), .B2(n9057), .ZN(
        n6368) );
  INV_X1 U2815 ( .A(n6369), .ZN(n11613) );
  AOI22_X1 U2816 ( .A1(ram[1865]), .A2(n6360), .B1(n11620), .B2(n9081), .ZN(
        n6369) );
  INV_X1 U2817 ( .A(n6370), .ZN(n11614) );
  AOI22_X1 U2818 ( .A1(ram[1866]), .A2(n6360), .B1(n11620), .B2(n9105), .ZN(
        n6370) );
  INV_X1 U2819 ( .A(n6371), .ZN(n11615) );
  AOI22_X1 U2820 ( .A1(ram[1867]), .A2(n6360), .B1(n11620), .B2(n9129), .ZN(
        n6371) );
  INV_X1 U2821 ( .A(n6372), .ZN(n11616) );
  AOI22_X1 U2822 ( .A1(ram[1868]), .A2(n6360), .B1(n11620), .B2(n9153), .ZN(
        n6372) );
  INV_X1 U2823 ( .A(n6373), .ZN(n11617) );
  AOI22_X1 U2824 ( .A1(ram[1869]), .A2(n6360), .B1(n11620), .B2(n9177), .ZN(
        n6373) );
  INV_X1 U2825 ( .A(n6374), .ZN(n11618) );
  AOI22_X1 U2826 ( .A1(ram[1870]), .A2(n6360), .B1(n11620), .B2(n9201), .ZN(
        n6374) );
  INV_X1 U2827 ( .A(n6375), .ZN(n11619) );
  AOI22_X1 U2828 ( .A1(ram[1871]), .A2(n6360), .B1(n11620), .B2(n9225), .ZN(
        n6375) );
  INV_X1 U2829 ( .A(n6393), .ZN(n11570) );
  AOI22_X1 U2830 ( .A1(ram[1888]), .A2(n6394), .B1(n11586), .B2(n8865), .ZN(
        n6393) );
  INV_X1 U2831 ( .A(n6395), .ZN(n11571) );
  AOI22_X1 U2832 ( .A1(ram[1889]), .A2(n6394), .B1(n11586), .B2(n8889), .ZN(
        n6395) );
  INV_X1 U2833 ( .A(n6396), .ZN(n11572) );
  AOI22_X1 U2834 ( .A1(ram[1890]), .A2(n6394), .B1(n11586), .B2(n8913), .ZN(
        n6396) );
  INV_X1 U2835 ( .A(n6397), .ZN(n11573) );
  AOI22_X1 U2836 ( .A1(ram[1891]), .A2(n6394), .B1(n11586), .B2(n8937), .ZN(
        n6397) );
  INV_X1 U2837 ( .A(n6398), .ZN(n11574) );
  AOI22_X1 U2838 ( .A1(ram[1892]), .A2(n6394), .B1(n11586), .B2(n8961), .ZN(
        n6398) );
  INV_X1 U2839 ( .A(n6399), .ZN(n11575) );
  AOI22_X1 U2840 ( .A1(ram[1893]), .A2(n6394), .B1(n11586), .B2(n8985), .ZN(
        n6399) );
  INV_X1 U2841 ( .A(n6400), .ZN(n11576) );
  AOI22_X1 U2842 ( .A1(ram[1894]), .A2(n6394), .B1(n11586), .B2(n9009), .ZN(
        n6400) );
  INV_X1 U2843 ( .A(n6401), .ZN(n11577) );
  AOI22_X1 U2844 ( .A1(ram[1895]), .A2(n6394), .B1(n11586), .B2(n9033), .ZN(
        n6401) );
  INV_X1 U2845 ( .A(n6402), .ZN(n11578) );
  AOI22_X1 U2846 ( .A1(ram[1896]), .A2(n6394), .B1(n11586), .B2(n9057), .ZN(
        n6402) );
  INV_X1 U2847 ( .A(n6403), .ZN(n11579) );
  AOI22_X1 U2848 ( .A1(ram[1897]), .A2(n6394), .B1(n11586), .B2(n9081), .ZN(
        n6403) );
  INV_X1 U2849 ( .A(n6404), .ZN(n11580) );
  AOI22_X1 U2850 ( .A1(ram[1898]), .A2(n6394), .B1(n11586), .B2(n9105), .ZN(
        n6404) );
  INV_X1 U2851 ( .A(n6405), .ZN(n11581) );
  AOI22_X1 U2852 ( .A1(ram[1899]), .A2(n6394), .B1(n11586), .B2(n9129), .ZN(
        n6405) );
  INV_X1 U2853 ( .A(n6406), .ZN(n11582) );
  AOI22_X1 U2854 ( .A1(ram[1900]), .A2(n6394), .B1(n11586), .B2(n9153), .ZN(
        n6406) );
  INV_X1 U2855 ( .A(n6407), .ZN(n11583) );
  AOI22_X1 U2856 ( .A1(ram[1901]), .A2(n6394), .B1(n11586), .B2(n9177), .ZN(
        n6407) );
  INV_X1 U2857 ( .A(n6408), .ZN(n11584) );
  AOI22_X1 U2858 ( .A1(ram[1902]), .A2(n6394), .B1(n11586), .B2(n9201), .ZN(
        n6408) );
  INV_X1 U2859 ( .A(n6409), .ZN(n11585) );
  AOI22_X1 U2860 ( .A1(ram[1903]), .A2(n6394), .B1(n11586), .B2(n9225), .ZN(
        n6409) );
  INV_X1 U2861 ( .A(n6427), .ZN(n11536) );
  AOI22_X1 U2862 ( .A1(ram[1920]), .A2(n6428), .B1(n11552), .B2(n8865), .ZN(
        n6427) );
  INV_X1 U2863 ( .A(n6429), .ZN(n11537) );
  AOI22_X1 U2864 ( .A1(ram[1921]), .A2(n6428), .B1(n11552), .B2(n8889), .ZN(
        n6429) );
  INV_X1 U2865 ( .A(n6430), .ZN(n11538) );
  AOI22_X1 U2866 ( .A1(ram[1922]), .A2(n6428), .B1(n11552), .B2(n8913), .ZN(
        n6430) );
  INV_X1 U2867 ( .A(n6431), .ZN(n11539) );
  AOI22_X1 U2868 ( .A1(ram[1923]), .A2(n6428), .B1(n11552), .B2(n8937), .ZN(
        n6431) );
  INV_X1 U2869 ( .A(n6432), .ZN(n11540) );
  AOI22_X1 U2870 ( .A1(ram[1924]), .A2(n6428), .B1(n11552), .B2(n8961), .ZN(
        n6432) );
  INV_X1 U2871 ( .A(n6433), .ZN(n11541) );
  AOI22_X1 U2872 ( .A1(ram[1925]), .A2(n6428), .B1(n11552), .B2(n8985), .ZN(
        n6433) );
  INV_X1 U2873 ( .A(n6434), .ZN(n11542) );
  AOI22_X1 U2874 ( .A1(ram[1926]), .A2(n6428), .B1(n11552), .B2(n9009), .ZN(
        n6434) );
  INV_X1 U2875 ( .A(n6435), .ZN(n11543) );
  AOI22_X1 U2876 ( .A1(ram[1927]), .A2(n6428), .B1(n11552), .B2(n9033), .ZN(
        n6435) );
  INV_X1 U2877 ( .A(n6436), .ZN(n11544) );
  AOI22_X1 U2878 ( .A1(ram[1928]), .A2(n6428), .B1(n11552), .B2(n9057), .ZN(
        n6436) );
  INV_X1 U2879 ( .A(n6437), .ZN(n11545) );
  AOI22_X1 U2880 ( .A1(ram[1929]), .A2(n6428), .B1(n11552), .B2(n9081), .ZN(
        n6437) );
  INV_X1 U2881 ( .A(n6438), .ZN(n11546) );
  AOI22_X1 U2882 ( .A1(ram[1930]), .A2(n6428), .B1(n11552), .B2(n9105), .ZN(
        n6438) );
  INV_X1 U2883 ( .A(n6439), .ZN(n11547) );
  AOI22_X1 U2884 ( .A1(ram[1931]), .A2(n6428), .B1(n11552), .B2(n9129), .ZN(
        n6439) );
  INV_X1 U2885 ( .A(n6440), .ZN(n11548) );
  AOI22_X1 U2886 ( .A1(ram[1932]), .A2(n6428), .B1(n11552), .B2(n9153), .ZN(
        n6440) );
  INV_X1 U2887 ( .A(n6441), .ZN(n11549) );
  AOI22_X1 U2888 ( .A1(ram[1933]), .A2(n6428), .B1(n11552), .B2(n9177), .ZN(
        n6441) );
  INV_X1 U2889 ( .A(n6442), .ZN(n11550) );
  AOI22_X1 U2890 ( .A1(ram[1934]), .A2(n6428), .B1(n11552), .B2(n9201), .ZN(
        n6442) );
  INV_X1 U2891 ( .A(n6443), .ZN(n11551) );
  AOI22_X1 U2892 ( .A1(ram[1935]), .A2(n6428), .B1(n11552), .B2(n9225), .ZN(
        n6443) );
  INV_X1 U2893 ( .A(n6461), .ZN(n11502) );
  AOI22_X1 U2894 ( .A1(ram[1952]), .A2(n6462), .B1(n11518), .B2(n8865), .ZN(
        n6461) );
  INV_X1 U2895 ( .A(n6463), .ZN(n11503) );
  AOI22_X1 U2896 ( .A1(ram[1953]), .A2(n6462), .B1(n11518), .B2(n8889), .ZN(
        n6463) );
  INV_X1 U2897 ( .A(n6464), .ZN(n11504) );
  AOI22_X1 U2898 ( .A1(ram[1954]), .A2(n6462), .B1(n11518), .B2(n8913), .ZN(
        n6464) );
  INV_X1 U2899 ( .A(n6465), .ZN(n11505) );
  AOI22_X1 U2900 ( .A1(ram[1955]), .A2(n6462), .B1(n11518), .B2(n8937), .ZN(
        n6465) );
  INV_X1 U2901 ( .A(n6466), .ZN(n11506) );
  AOI22_X1 U2902 ( .A1(ram[1956]), .A2(n6462), .B1(n11518), .B2(n8961), .ZN(
        n6466) );
  INV_X1 U2903 ( .A(n6467), .ZN(n11507) );
  AOI22_X1 U2904 ( .A1(ram[1957]), .A2(n6462), .B1(n11518), .B2(n8985), .ZN(
        n6467) );
  INV_X1 U2905 ( .A(n6468), .ZN(n11508) );
  AOI22_X1 U2906 ( .A1(ram[1958]), .A2(n6462), .B1(n11518), .B2(n9009), .ZN(
        n6468) );
  INV_X1 U2907 ( .A(n6469), .ZN(n11509) );
  AOI22_X1 U2908 ( .A1(ram[1959]), .A2(n6462), .B1(n11518), .B2(n9033), .ZN(
        n6469) );
  INV_X1 U2909 ( .A(n6470), .ZN(n11510) );
  AOI22_X1 U2910 ( .A1(ram[1960]), .A2(n6462), .B1(n11518), .B2(n9057), .ZN(
        n6470) );
  INV_X1 U2911 ( .A(n6471), .ZN(n11511) );
  AOI22_X1 U2912 ( .A1(ram[1961]), .A2(n6462), .B1(n11518), .B2(n9081), .ZN(
        n6471) );
  INV_X1 U2913 ( .A(n6472), .ZN(n11512) );
  AOI22_X1 U2914 ( .A1(ram[1962]), .A2(n6462), .B1(n11518), .B2(n9105), .ZN(
        n6472) );
  INV_X1 U2915 ( .A(n6473), .ZN(n11513) );
  AOI22_X1 U2916 ( .A1(ram[1963]), .A2(n6462), .B1(n11518), .B2(n9129), .ZN(
        n6473) );
  INV_X1 U2917 ( .A(n6474), .ZN(n11514) );
  AOI22_X1 U2918 ( .A1(ram[1964]), .A2(n6462), .B1(n11518), .B2(n9153), .ZN(
        n6474) );
  INV_X1 U2919 ( .A(n6475), .ZN(n11515) );
  AOI22_X1 U2920 ( .A1(ram[1965]), .A2(n6462), .B1(n11518), .B2(n9177), .ZN(
        n6475) );
  INV_X1 U2921 ( .A(n6476), .ZN(n11516) );
  AOI22_X1 U2922 ( .A1(ram[1966]), .A2(n6462), .B1(n11518), .B2(n9201), .ZN(
        n6476) );
  INV_X1 U2923 ( .A(n6477), .ZN(n11517) );
  AOI22_X1 U2924 ( .A1(ram[1967]), .A2(n6462), .B1(n11518), .B2(n9225), .ZN(
        n6477) );
  INV_X1 U2925 ( .A(n6495), .ZN(n11468) );
  AOI22_X1 U2926 ( .A1(ram[1984]), .A2(n6496), .B1(n11484), .B2(n8864), .ZN(
        n6495) );
  INV_X1 U2927 ( .A(n6497), .ZN(n11469) );
  AOI22_X1 U2928 ( .A1(ram[1985]), .A2(n6496), .B1(n11484), .B2(n8888), .ZN(
        n6497) );
  INV_X1 U2929 ( .A(n6498), .ZN(n11470) );
  AOI22_X1 U2930 ( .A1(ram[1986]), .A2(n6496), .B1(n11484), .B2(n8912), .ZN(
        n6498) );
  INV_X1 U2931 ( .A(n6499), .ZN(n11471) );
  AOI22_X1 U2932 ( .A1(ram[1987]), .A2(n6496), .B1(n11484), .B2(n8936), .ZN(
        n6499) );
  INV_X1 U2933 ( .A(n6500), .ZN(n11472) );
  AOI22_X1 U2934 ( .A1(ram[1988]), .A2(n6496), .B1(n11484), .B2(n8960), .ZN(
        n6500) );
  INV_X1 U2935 ( .A(n6501), .ZN(n11473) );
  AOI22_X1 U2936 ( .A1(ram[1989]), .A2(n6496), .B1(n11484), .B2(n8984), .ZN(
        n6501) );
  INV_X1 U2937 ( .A(n6502), .ZN(n11474) );
  AOI22_X1 U2938 ( .A1(ram[1990]), .A2(n6496), .B1(n11484), .B2(n9008), .ZN(
        n6502) );
  INV_X1 U2939 ( .A(n6503), .ZN(n11475) );
  AOI22_X1 U2940 ( .A1(ram[1991]), .A2(n6496), .B1(n11484), .B2(n9032), .ZN(
        n6503) );
  INV_X1 U2941 ( .A(n6504), .ZN(n11476) );
  AOI22_X1 U2942 ( .A1(ram[1992]), .A2(n6496), .B1(n11484), .B2(n9056), .ZN(
        n6504) );
  INV_X1 U2943 ( .A(n6505), .ZN(n11477) );
  AOI22_X1 U2944 ( .A1(ram[1993]), .A2(n6496), .B1(n11484), .B2(n9080), .ZN(
        n6505) );
  INV_X1 U2945 ( .A(n6506), .ZN(n11478) );
  AOI22_X1 U2946 ( .A1(ram[1994]), .A2(n6496), .B1(n11484), .B2(n9104), .ZN(
        n6506) );
  INV_X1 U2947 ( .A(n6507), .ZN(n11479) );
  AOI22_X1 U2948 ( .A1(ram[1995]), .A2(n6496), .B1(n11484), .B2(n9128), .ZN(
        n6507) );
  INV_X1 U2949 ( .A(n6508), .ZN(n11480) );
  AOI22_X1 U2950 ( .A1(ram[1996]), .A2(n6496), .B1(n11484), .B2(n9152), .ZN(
        n6508) );
  INV_X1 U2951 ( .A(n6509), .ZN(n11481) );
  AOI22_X1 U2952 ( .A1(ram[1997]), .A2(n6496), .B1(n11484), .B2(n9176), .ZN(
        n6509) );
  INV_X1 U2953 ( .A(n6510), .ZN(n11482) );
  AOI22_X1 U2954 ( .A1(ram[1998]), .A2(n6496), .B1(n11484), .B2(n9200), .ZN(
        n6510) );
  INV_X1 U2955 ( .A(n6511), .ZN(n11483) );
  AOI22_X1 U2956 ( .A1(ram[1999]), .A2(n6496), .B1(n11484), .B2(n9224), .ZN(
        n6511) );
  INV_X1 U2957 ( .A(n6529), .ZN(n11434) );
  AOI22_X1 U2958 ( .A1(ram[2016]), .A2(n6530), .B1(n11450), .B2(n8864), .ZN(
        n6529) );
  INV_X1 U2959 ( .A(n6531), .ZN(n11435) );
  AOI22_X1 U2960 ( .A1(ram[2017]), .A2(n6530), .B1(n11450), .B2(n8888), .ZN(
        n6531) );
  INV_X1 U2961 ( .A(n6532), .ZN(n11436) );
  AOI22_X1 U2962 ( .A1(ram[2018]), .A2(n6530), .B1(n11450), .B2(n8912), .ZN(
        n6532) );
  INV_X1 U2963 ( .A(n6533), .ZN(n11437) );
  AOI22_X1 U2964 ( .A1(ram[2019]), .A2(n6530), .B1(n11450), .B2(n8936), .ZN(
        n6533) );
  INV_X1 U2965 ( .A(n6534), .ZN(n11438) );
  AOI22_X1 U2966 ( .A1(ram[2020]), .A2(n6530), .B1(n11450), .B2(n8960), .ZN(
        n6534) );
  INV_X1 U2967 ( .A(n6535), .ZN(n11439) );
  AOI22_X1 U2968 ( .A1(ram[2021]), .A2(n6530), .B1(n11450), .B2(n8984), .ZN(
        n6535) );
  INV_X1 U2969 ( .A(n6536), .ZN(n11440) );
  AOI22_X1 U2970 ( .A1(ram[2022]), .A2(n6530), .B1(n11450), .B2(n9008), .ZN(
        n6536) );
  INV_X1 U2971 ( .A(n6537), .ZN(n11441) );
  AOI22_X1 U2972 ( .A1(ram[2023]), .A2(n6530), .B1(n11450), .B2(n9032), .ZN(
        n6537) );
  INV_X1 U2973 ( .A(n6538), .ZN(n11442) );
  AOI22_X1 U2974 ( .A1(ram[2024]), .A2(n6530), .B1(n11450), .B2(n9056), .ZN(
        n6538) );
  INV_X1 U2975 ( .A(n6539), .ZN(n11443) );
  AOI22_X1 U2976 ( .A1(ram[2025]), .A2(n6530), .B1(n11450), .B2(n9080), .ZN(
        n6539) );
  INV_X1 U2977 ( .A(n6540), .ZN(n11444) );
  AOI22_X1 U2978 ( .A1(ram[2026]), .A2(n6530), .B1(n11450), .B2(n9104), .ZN(
        n6540) );
  INV_X1 U2979 ( .A(n6541), .ZN(n11445) );
  AOI22_X1 U2980 ( .A1(ram[2027]), .A2(n6530), .B1(n11450), .B2(n9128), .ZN(
        n6541) );
  INV_X1 U2981 ( .A(n6542), .ZN(n11446) );
  AOI22_X1 U2982 ( .A1(ram[2028]), .A2(n6530), .B1(n11450), .B2(n9152), .ZN(
        n6542) );
  INV_X1 U2983 ( .A(n6543), .ZN(n11447) );
  AOI22_X1 U2984 ( .A1(ram[2029]), .A2(n6530), .B1(n11450), .B2(n9176), .ZN(
        n6543) );
  INV_X1 U2985 ( .A(n6544), .ZN(n11448) );
  AOI22_X1 U2986 ( .A1(ram[2030]), .A2(n6530), .B1(n11450), .B2(n9200), .ZN(
        n6544) );
  INV_X1 U2987 ( .A(n6545), .ZN(n11449) );
  AOI22_X1 U2988 ( .A1(ram[2031]), .A2(n6530), .B1(n11450), .B2(n9224), .ZN(
        n6545) );
  INV_X1 U2989 ( .A(n6563), .ZN(n11400) );
  AOI22_X1 U2990 ( .A1(ram[2048]), .A2(n6564), .B1(n11416), .B2(n8864), .ZN(
        n6563) );
  INV_X1 U2991 ( .A(n6565), .ZN(n11401) );
  AOI22_X1 U2992 ( .A1(ram[2049]), .A2(n6564), .B1(n11416), .B2(n8888), .ZN(
        n6565) );
  INV_X1 U2993 ( .A(n6566), .ZN(n11402) );
  AOI22_X1 U2994 ( .A1(ram[2050]), .A2(n6564), .B1(n11416), .B2(n8912), .ZN(
        n6566) );
  INV_X1 U2995 ( .A(n6567), .ZN(n11403) );
  AOI22_X1 U2996 ( .A1(ram[2051]), .A2(n6564), .B1(n11416), .B2(n8936), .ZN(
        n6567) );
  INV_X1 U2997 ( .A(n6568), .ZN(n11404) );
  AOI22_X1 U2998 ( .A1(ram[2052]), .A2(n6564), .B1(n11416), .B2(n8960), .ZN(
        n6568) );
  INV_X1 U2999 ( .A(n6569), .ZN(n11405) );
  AOI22_X1 U3000 ( .A1(ram[2053]), .A2(n6564), .B1(n11416), .B2(n8984), .ZN(
        n6569) );
  INV_X1 U3001 ( .A(n6570), .ZN(n11406) );
  AOI22_X1 U3002 ( .A1(ram[2054]), .A2(n6564), .B1(n11416), .B2(n9008), .ZN(
        n6570) );
  INV_X1 U3003 ( .A(n6571), .ZN(n11407) );
  AOI22_X1 U3004 ( .A1(ram[2055]), .A2(n6564), .B1(n11416), .B2(n9032), .ZN(
        n6571) );
  INV_X1 U3005 ( .A(n6572), .ZN(n11408) );
  AOI22_X1 U3006 ( .A1(ram[2056]), .A2(n6564), .B1(n11416), .B2(n9056), .ZN(
        n6572) );
  INV_X1 U3007 ( .A(n6573), .ZN(n11409) );
  AOI22_X1 U3008 ( .A1(ram[2057]), .A2(n6564), .B1(n11416), .B2(n9080), .ZN(
        n6573) );
  INV_X1 U3009 ( .A(n6574), .ZN(n11410) );
  AOI22_X1 U3010 ( .A1(ram[2058]), .A2(n6564), .B1(n11416), .B2(n9104), .ZN(
        n6574) );
  INV_X1 U3011 ( .A(n6575), .ZN(n11411) );
  AOI22_X1 U3012 ( .A1(ram[2059]), .A2(n6564), .B1(n11416), .B2(n9128), .ZN(
        n6575) );
  INV_X1 U3013 ( .A(n6576), .ZN(n11412) );
  AOI22_X1 U3014 ( .A1(ram[2060]), .A2(n6564), .B1(n11416), .B2(n9152), .ZN(
        n6576) );
  INV_X1 U3015 ( .A(n6577), .ZN(n11413) );
  AOI22_X1 U3016 ( .A1(ram[2061]), .A2(n6564), .B1(n11416), .B2(n9176), .ZN(
        n6577) );
  INV_X1 U3017 ( .A(n6578), .ZN(n11414) );
  AOI22_X1 U3018 ( .A1(ram[2062]), .A2(n6564), .B1(n11416), .B2(n9200), .ZN(
        n6578) );
  INV_X1 U3019 ( .A(n6579), .ZN(n11415) );
  AOI22_X1 U3020 ( .A1(ram[2063]), .A2(n6564), .B1(n11416), .B2(n9224), .ZN(
        n6579) );
  INV_X1 U3021 ( .A(n6598), .ZN(n11366) );
  AOI22_X1 U3022 ( .A1(ram[2080]), .A2(n6599), .B1(n11382), .B2(n8864), .ZN(
        n6598) );
  INV_X1 U3023 ( .A(n6600), .ZN(n11367) );
  AOI22_X1 U3024 ( .A1(ram[2081]), .A2(n6599), .B1(n11382), .B2(n8888), .ZN(
        n6600) );
  INV_X1 U3025 ( .A(n6601), .ZN(n11368) );
  AOI22_X1 U3026 ( .A1(ram[2082]), .A2(n6599), .B1(n11382), .B2(n8912), .ZN(
        n6601) );
  INV_X1 U3027 ( .A(n6602), .ZN(n11369) );
  AOI22_X1 U3028 ( .A1(ram[2083]), .A2(n6599), .B1(n11382), .B2(n8936), .ZN(
        n6602) );
  INV_X1 U3029 ( .A(n6603), .ZN(n11370) );
  AOI22_X1 U3030 ( .A1(ram[2084]), .A2(n6599), .B1(n11382), .B2(n8960), .ZN(
        n6603) );
  INV_X1 U3031 ( .A(n6604), .ZN(n11371) );
  AOI22_X1 U3032 ( .A1(ram[2085]), .A2(n6599), .B1(n11382), .B2(n8984), .ZN(
        n6604) );
  INV_X1 U3033 ( .A(n6605), .ZN(n11372) );
  AOI22_X1 U3034 ( .A1(ram[2086]), .A2(n6599), .B1(n11382), .B2(n9008), .ZN(
        n6605) );
  INV_X1 U3035 ( .A(n6606), .ZN(n11373) );
  AOI22_X1 U3036 ( .A1(ram[2087]), .A2(n6599), .B1(n11382), .B2(n9032), .ZN(
        n6606) );
  INV_X1 U3037 ( .A(n6607), .ZN(n11374) );
  AOI22_X1 U3038 ( .A1(ram[2088]), .A2(n6599), .B1(n11382), .B2(n9056), .ZN(
        n6607) );
  INV_X1 U3039 ( .A(n6608), .ZN(n11375) );
  AOI22_X1 U3040 ( .A1(ram[2089]), .A2(n6599), .B1(n11382), .B2(n9080), .ZN(
        n6608) );
  INV_X1 U3041 ( .A(n6609), .ZN(n11376) );
  AOI22_X1 U3042 ( .A1(ram[2090]), .A2(n6599), .B1(n11382), .B2(n9104), .ZN(
        n6609) );
  INV_X1 U3043 ( .A(n6610), .ZN(n11377) );
  AOI22_X1 U3044 ( .A1(ram[2091]), .A2(n6599), .B1(n11382), .B2(n9128), .ZN(
        n6610) );
  INV_X1 U3045 ( .A(n6611), .ZN(n11378) );
  AOI22_X1 U3046 ( .A1(ram[2092]), .A2(n6599), .B1(n11382), .B2(n9152), .ZN(
        n6611) );
  INV_X1 U3047 ( .A(n6612), .ZN(n11379) );
  AOI22_X1 U3048 ( .A1(ram[2093]), .A2(n6599), .B1(n11382), .B2(n9176), .ZN(
        n6612) );
  INV_X1 U3049 ( .A(n6613), .ZN(n11380) );
  AOI22_X1 U3050 ( .A1(ram[2094]), .A2(n6599), .B1(n11382), .B2(n9200), .ZN(
        n6613) );
  INV_X1 U3051 ( .A(n6614), .ZN(n11381) );
  AOI22_X1 U3052 ( .A1(ram[2095]), .A2(n6599), .B1(n11382), .B2(n9224), .ZN(
        n6614) );
  INV_X1 U3053 ( .A(n6632), .ZN(n11332) );
  AOI22_X1 U3054 ( .A1(ram[2112]), .A2(n6633), .B1(n11348), .B2(n8864), .ZN(
        n6632) );
  INV_X1 U3055 ( .A(n6634), .ZN(n11333) );
  AOI22_X1 U3056 ( .A1(ram[2113]), .A2(n6633), .B1(n11348), .B2(n8888), .ZN(
        n6634) );
  INV_X1 U3057 ( .A(n6635), .ZN(n11334) );
  AOI22_X1 U3058 ( .A1(ram[2114]), .A2(n6633), .B1(n11348), .B2(n8912), .ZN(
        n6635) );
  INV_X1 U3059 ( .A(n6636), .ZN(n11335) );
  AOI22_X1 U3060 ( .A1(ram[2115]), .A2(n6633), .B1(n11348), .B2(n8936), .ZN(
        n6636) );
  INV_X1 U3061 ( .A(n6637), .ZN(n11336) );
  AOI22_X1 U3062 ( .A1(ram[2116]), .A2(n6633), .B1(n11348), .B2(n8960), .ZN(
        n6637) );
  INV_X1 U3063 ( .A(n6638), .ZN(n11337) );
  AOI22_X1 U3064 ( .A1(ram[2117]), .A2(n6633), .B1(n11348), .B2(n8984), .ZN(
        n6638) );
  INV_X1 U3065 ( .A(n6639), .ZN(n11338) );
  AOI22_X1 U3066 ( .A1(ram[2118]), .A2(n6633), .B1(n11348), .B2(n9008), .ZN(
        n6639) );
  INV_X1 U3067 ( .A(n6640), .ZN(n11339) );
  AOI22_X1 U3068 ( .A1(ram[2119]), .A2(n6633), .B1(n11348), .B2(n9032), .ZN(
        n6640) );
  INV_X1 U3069 ( .A(n6641), .ZN(n11340) );
  AOI22_X1 U3070 ( .A1(ram[2120]), .A2(n6633), .B1(n11348), .B2(n9056), .ZN(
        n6641) );
  INV_X1 U3071 ( .A(n6642), .ZN(n11341) );
  AOI22_X1 U3072 ( .A1(ram[2121]), .A2(n6633), .B1(n11348), .B2(n9080), .ZN(
        n6642) );
  INV_X1 U3073 ( .A(n6643), .ZN(n11342) );
  AOI22_X1 U3074 ( .A1(ram[2122]), .A2(n6633), .B1(n11348), .B2(n9104), .ZN(
        n6643) );
  INV_X1 U3075 ( .A(n6644), .ZN(n11343) );
  AOI22_X1 U3076 ( .A1(ram[2123]), .A2(n6633), .B1(n11348), .B2(n9128), .ZN(
        n6644) );
  INV_X1 U3077 ( .A(n6645), .ZN(n11344) );
  AOI22_X1 U3078 ( .A1(ram[2124]), .A2(n6633), .B1(n11348), .B2(n9152), .ZN(
        n6645) );
  INV_X1 U3079 ( .A(n6646), .ZN(n11345) );
  AOI22_X1 U3080 ( .A1(ram[2125]), .A2(n6633), .B1(n11348), .B2(n9176), .ZN(
        n6646) );
  INV_X1 U3081 ( .A(n6647), .ZN(n11346) );
  AOI22_X1 U3082 ( .A1(ram[2126]), .A2(n6633), .B1(n11348), .B2(n9200), .ZN(
        n6647) );
  INV_X1 U3083 ( .A(n6648), .ZN(n11347) );
  AOI22_X1 U3084 ( .A1(ram[2127]), .A2(n6633), .B1(n11348), .B2(n9224), .ZN(
        n6648) );
  INV_X1 U3085 ( .A(n6666), .ZN(n11298) );
  AOI22_X1 U3086 ( .A1(ram[2144]), .A2(n6667), .B1(n11314), .B2(n8864), .ZN(
        n6666) );
  INV_X1 U3087 ( .A(n6668), .ZN(n11299) );
  AOI22_X1 U3088 ( .A1(ram[2145]), .A2(n6667), .B1(n11314), .B2(n8888), .ZN(
        n6668) );
  INV_X1 U3089 ( .A(n6669), .ZN(n11300) );
  AOI22_X1 U3090 ( .A1(ram[2146]), .A2(n6667), .B1(n11314), .B2(n8912), .ZN(
        n6669) );
  INV_X1 U3091 ( .A(n6670), .ZN(n11301) );
  AOI22_X1 U3092 ( .A1(ram[2147]), .A2(n6667), .B1(n11314), .B2(n8936), .ZN(
        n6670) );
  INV_X1 U3093 ( .A(n6671), .ZN(n11302) );
  AOI22_X1 U3094 ( .A1(ram[2148]), .A2(n6667), .B1(n11314), .B2(n8960), .ZN(
        n6671) );
  INV_X1 U3095 ( .A(n6672), .ZN(n11303) );
  AOI22_X1 U3096 ( .A1(ram[2149]), .A2(n6667), .B1(n11314), .B2(n8984), .ZN(
        n6672) );
  INV_X1 U3097 ( .A(n6673), .ZN(n11304) );
  AOI22_X1 U3098 ( .A1(ram[2150]), .A2(n6667), .B1(n11314), .B2(n9008), .ZN(
        n6673) );
  INV_X1 U3099 ( .A(n6674), .ZN(n11305) );
  AOI22_X1 U3100 ( .A1(ram[2151]), .A2(n6667), .B1(n11314), .B2(n9032), .ZN(
        n6674) );
  INV_X1 U3101 ( .A(n6675), .ZN(n11306) );
  AOI22_X1 U3102 ( .A1(ram[2152]), .A2(n6667), .B1(n11314), .B2(n9056), .ZN(
        n6675) );
  INV_X1 U3103 ( .A(n6676), .ZN(n11307) );
  AOI22_X1 U3104 ( .A1(ram[2153]), .A2(n6667), .B1(n11314), .B2(n9080), .ZN(
        n6676) );
  INV_X1 U3105 ( .A(n6677), .ZN(n11308) );
  AOI22_X1 U3106 ( .A1(ram[2154]), .A2(n6667), .B1(n11314), .B2(n9104), .ZN(
        n6677) );
  INV_X1 U3107 ( .A(n6678), .ZN(n11309) );
  AOI22_X1 U3108 ( .A1(ram[2155]), .A2(n6667), .B1(n11314), .B2(n9128), .ZN(
        n6678) );
  INV_X1 U3109 ( .A(n6679), .ZN(n11310) );
  AOI22_X1 U3110 ( .A1(ram[2156]), .A2(n6667), .B1(n11314), .B2(n9152), .ZN(
        n6679) );
  INV_X1 U3111 ( .A(n6680), .ZN(n11311) );
  AOI22_X1 U3112 ( .A1(ram[2157]), .A2(n6667), .B1(n11314), .B2(n9176), .ZN(
        n6680) );
  INV_X1 U3113 ( .A(n6681), .ZN(n11312) );
  AOI22_X1 U3114 ( .A1(ram[2158]), .A2(n6667), .B1(n11314), .B2(n9200), .ZN(
        n6681) );
  INV_X1 U3115 ( .A(n6682), .ZN(n11313) );
  AOI22_X1 U3116 ( .A1(ram[2159]), .A2(n6667), .B1(n11314), .B2(n9224), .ZN(
        n6682) );
  INV_X1 U3117 ( .A(n6700), .ZN(n11264) );
  AOI22_X1 U3118 ( .A1(ram[2176]), .A2(n6701), .B1(n11280), .B2(n8863), .ZN(
        n6700) );
  INV_X1 U3119 ( .A(n6702), .ZN(n11265) );
  AOI22_X1 U3120 ( .A1(ram[2177]), .A2(n6701), .B1(n11280), .B2(n8887), .ZN(
        n6702) );
  INV_X1 U3121 ( .A(n6703), .ZN(n11266) );
  AOI22_X1 U3122 ( .A1(ram[2178]), .A2(n6701), .B1(n11280), .B2(n8911), .ZN(
        n6703) );
  INV_X1 U3123 ( .A(n6704), .ZN(n11267) );
  AOI22_X1 U3124 ( .A1(ram[2179]), .A2(n6701), .B1(n11280), .B2(n8935), .ZN(
        n6704) );
  INV_X1 U3125 ( .A(n6705), .ZN(n11268) );
  AOI22_X1 U3126 ( .A1(ram[2180]), .A2(n6701), .B1(n11280), .B2(n8959), .ZN(
        n6705) );
  INV_X1 U3127 ( .A(n6706), .ZN(n11269) );
  AOI22_X1 U3128 ( .A1(ram[2181]), .A2(n6701), .B1(n11280), .B2(n8983), .ZN(
        n6706) );
  INV_X1 U3129 ( .A(n6707), .ZN(n11270) );
  AOI22_X1 U3130 ( .A1(ram[2182]), .A2(n6701), .B1(n11280), .B2(n9007), .ZN(
        n6707) );
  INV_X1 U3131 ( .A(n6708), .ZN(n11271) );
  AOI22_X1 U3132 ( .A1(ram[2183]), .A2(n6701), .B1(n11280), .B2(n9031), .ZN(
        n6708) );
  INV_X1 U3133 ( .A(n6709), .ZN(n11272) );
  AOI22_X1 U3134 ( .A1(ram[2184]), .A2(n6701), .B1(n11280), .B2(n9055), .ZN(
        n6709) );
  INV_X1 U3135 ( .A(n6710), .ZN(n11273) );
  AOI22_X1 U3136 ( .A1(ram[2185]), .A2(n6701), .B1(n11280), .B2(n9079), .ZN(
        n6710) );
  INV_X1 U3137 ( .A(n6711), .ZN(n11274) );
  AOI22_X1 U3138 ( .A1(ram[2186]), .A2(n6701), .B1(n11280), .B2(n9103), .ZN(
        n6711) );
  INV_X1 U3139 ( .A(n6712), .ZN(n11275) );
  AOI22_X1 U3140 ( .A1(ram[2187]), .A2(n6701), .B1(n11280), .B2(n9127), .ZN(
        n6712) );
  INV_X1 U3141 ( .A(n6713), .ZN(n11276) );
  AOI22_X1 U3142 ( .A1(ram[2188]), .A2(n6701), .B1(n11280), .B2(n9151), .ZN(
        n6713) );
  INV_X1 U3143 ( .A(n6714), .ZN(n11277) );
  AOI22_X1 U3144 ( .A1(ram[2189]), .A2(n6701), .B1(n11280), .B2(n9175), .ZN(
        n6714) );
  INV_X1 U3145 ( .A(n6715), .ZN(n11278) );
  AOI22_X1 U3146 ( .A1(ram[2190]), .A2(n6701), .B1(n11280), .B2(n9199), .ZN(
        n6715) );
  INV_X1 U3147 ( .A(n6716), .ZN(n11279) );
  AOI22_X1 U3148 ( .A1(ram[2191]), .A2(n6701), .B1(n11280), .B2(n9223), .ZN(
        n6716) );
  INV_X1 U3149 ( .A(n6734), .ZN(n11230) );
  AOI22_X1 U3150 ( .A1(ram[2208]), .A2(n6735), .B1(n11246), .B2(n8863), .ZN(
        n6734) );
  INV_X1 U3151 ( .A(n6736), .ZN(n11231) );
  AOI22_X1 U3152 ( .A1(ram[2209]), .A2(n6735), .B1(n11246), .B2(n8887), .ZN(
        n6736) );
  INV_X1 U3153 ( .A(n6737), .ZN(n11232) );
  AOI22_X1 U3154 ( .A1(ram[2210]), .A2(n6735), .B1(n11246), .B2(n8911), .ZN(
        n6737) );
  INV_X1 U3155 ( .A(n6738), .ZN(n11233) );
  AOI22_X1 U3156 ( .A1(ram[2211]), .A2(n6735), .B1(n11246), .B2(n8935), .ZN(
        n6738) );
  INV_X1 U3157 ( .A(n6739), .ZN(n11234) );
  AOI22_X1 U3158 ( .A1(ram[2212]), .A2(n6735), .B1(n11246), .B2(n8959), .ZN(
        n6739) );
  INV_X1 U3159 ( .A(n6740), .ZN(n11235) );
  AOI22_X1 U3160 ( .A1(ram[2213]), .A2(n6735), .B1(n11246), .B2(n8983), .ZN(
        n6740) );
  INV_X1 U3161 ( .A(n6741), .ZN(n11236) );
  AOI22_X1 U3162 ( .A1(ram[2214]), .A2(n6735), .B1(n11246), .B2(n9007), .ZN(
        n6741) );
  INV_X1 U3163 ( .A(n6742), .ZN(n11237) );
  AOI22_X1 U3164 ( .A1(ram[2215]), .A2(n6735), .B1(n11246), .B2(n9031), .ZN(
        n6742) );
  INV_X1 U3165 ( .A(n6743), .ZN(n11238) );
  AOI22_X1 U3166 ( .A1(ram[2216]), .A2(n6735), .B1(n11246), .B2(n9055), .ZN(
        n6743) );
  INV_X1 U3167 ( .A(n6744), .ZN(n11239) );
  AOI22_X1 U3168 ( .A1(ram[2217]), .A2(n6735), .B1(n11246), .B2(n9079), .ZN(
        n6744) );
  INV_X1 U3169 ( .A(n6745), .ZN(n11240) );
  AOI22_X1 U3170 ( .A1(ram[2218]), .A2(n6735), .B1(n11246), .B2(n9103), .ZN(
        n6745) );
  INV_X1 U3171 ( .A(n6746), .ZN(n11241) );
  AOI22_X1 U3172 ( .A1(ram[2219]), .A2(n6735), .B1(n11246), .B2(n9127), .ZN(
        n6746) );
  INV_X1 U3173 ( .A(n6747), .ZN(n11242) );
  AOI22_X1 U3174 ( .A1(ram[2220]), .A2(n6735), .B1(n11246), .B2(n9151), .ZN(
        n6747) );
  INV_X1 U3175 ( .A(n6748), .ZN(n11243) );
  AOI22_X1 U3176 ( .A1(ram[2221]), .A2(n6735), .B1(n11246), .B2(n9175), .ZN(
        n6748) );
  INV_X1 U3177 ( .A(n6749), .ZN(n11244) );
  AOI22_X1 U3178 ( .A1(ram[2222]), .A2(n6735), .B1(n11246), .B2(n9199), .ZN(
        n6749) );
  INV_X1 U3179 ( .A(n6750), .ZN(n11245) );
  AOI22_X1 U3180 ( .A1(ram[2223]), .A2(n6735), .B1(n11246), .B2(n9223), .ZN(
        n6750) );
  INV_X1 U3181 ( .A(n6768), .ZN(n11196) );
  AOI22_X1 U3182 ( .A1(ram[2240]), .A2(n6769), .B1(n11212), .B2(n8863), .ZN(
        n6768) );
  INV_X1 U3183 ( .A(n6770), .ZN(n11197) );
  AOI22_X1 U3184 ( .A1(ram[2241]), .A2(n6769), .B1(n11212), .B2(n8887), .ZN(
        n6770) );
  INV_X1 U3185 ( .A(n6771), .ZN(n11198) );
  AOI22_X1 U3186 ( .A1(ram[2242]), .A2(n6769), .B1(n11212), .B2(n8911), .ZN(
        n6771) );
  INV_X1 U3187 ( .A(n6772), .ZN(n11199) );
  AOI22_X1 U3188 ( .A1(ram[2243]), .A2(n6769), .B1(n11212), .B2(n8935), .ZN(
        n6772) );
  INV_X1 U3189 ( .A(n6773), .ZN(n11200) );
  AOI22_X1 U3190 ( .A1(ram[2244]), .A2(n6769), .B1(n11212), .B2(n8959), .ZN(
        n6773) );
  INV_X1 U3191 ( .A(n6774), .ZN(n11201) );
  AOI22_X1 U3192 ( .A1(ram[2245]), .A2(n6769), .B1(n11212), .B2(n8983), .ZN(
        n6774) );
  INV_X1 U3193 ( .A(n6775), .ZN(n11202) );
  AOI22_X1 U3194 ( .A1(ram[2246]), .A2(n6769), .B1(n11212), .B2(n9007), .ZN(
        n6775) );
  INV_X1 U3195 ( .A(n6776), .ZN(n11203) );
  AOI22_X1 U3196 ( .A1(ram[2247]), .A2(n6769), .B1(n11212), .B2(n9031), .ZN(
        n6776) );
  INV_X1 U3197 ( .A(n6777), .ZN(n11204) );
  AOI22_X1 U3198 ( .A1(ram[2248]), .A2(n6769), .B1(n11212), .B2(n9055), .ZN(
        n6777) );
  INV_X1 U3199 ( .A(n6778), .ZN(n11205) );
  AOI22_X1 U3200 ( .A1(ram[2249]), .A2(n6769), .B1(n11212), .B2(n9079), .ZN(
        n6778) );
  INV_X1 U3201 ( .A(n6779), .ZN(n11206) );
  AOI22_X1 U3202 ( .A1(ram[2250]), .A2(n6769), .B1(n11212), .B2(n9103), .ZN(
        n6779) );
  INV_X1 U3203 ( .A(n6780), .ZN(n11207) );
  AOI22_X1 U3204 ( .A1(ram[2251]), .A2(n6769), .B1(n11212), .B2(n9127), .ZN(
        n6780) );
  INV_X1 U3205 ( .A(n6781), .ZN(n11208) );
  AOI22_X1 U3206 ( .A1(ram[2252]), .A2(n6769), .B1(n11212), .B2(n9151), .ZN(
        n6781) );
  INV_X1 U3207 ( .A(n6782), .ZN(n11209) );
  AOI22_X1 U3208 ( .A1(ram[2253]), .A2(n6769), .B1(n11212), .B2(n9175), .ZN(
        n6782) );
  INV_X1 U3209 ( .A(n6783), .ZN(n11210) );
  AOI22_X1 U3210 ( .A1(ram[2254]), .A2(n6769), .B1(n11212), .B2(n9199), .ZN(
        n6783) );
  INV_X1 U3211 ( .A(n6784), .ZN(n11211) );
  AOI22_X1 U3212 ( .A1(ram[2255]), .A2(n6769), .B1(n11212), .B2(n9223), .ZN(
        n6784) );
  INV_X1 U3213 ( .A(n6802), .ZN(n11162) );
  AOI22_X1 U3214 ( .A1(ram[2272]), .A2(n6803), .B1(n11178), .B2(n8863), .ZN(
        n6802) );
  INV_X1 U3215 ( .A(n6804), .ZN(n11163) );
  AOI22_X1 U3216 ( .A1(ram[2273]), .A2(n6803), .B1(n11178), .B2(n8887), .ZN(
        n6804) );
  INV_X1 U3217 ( .A(n6805), .ZN(n11164) );
  AOI22_X1 U3218 ( .A1(ram[2274]), .A2(n6803), .B1(n11178), .B2(n8911), .ZN(
        n6805) );
  INV_X1 U3219 ( .A(n6806), .ZN(n11165) );
  AOI22_X1 U3220 ( .A1(ram[2275]), .A2(n6803), .B1(n11178), .B2(n8935), .ZN(
        n6806) );
  INV_X1 U3221 ( .A(n6807), .ZN(n11166) );
  AOI22_X1 U3222 ( .A1(ram[2276]), .A2(n6803), .B1(n11178), .B2(n8959), .ZN(
        n6807) );
  INV_X1 U3223 ( .A(n6808), .ZN(n11167) );
  AOI22_X1 U3224 ( .A1(ram[2277]), .A2(n6803), .B1(n11178), .B2(n8983), .ZN(
        n6808) );
  INV_X1 U3225 ( .A(n6809), .ZN(n11168) );
  AOI22_X1 U3226 ( .A1(ram[2278]), .A2(n6803), .B1(n11178), .B2(n9007), .ZN(
        n6809) );
  INV_X1 U3227 ( .A(n6810), .ZN(n11169) );
  AOI22_X1 U3228 ( .A1(ram[2279]), .A2(n6803), .B1(n11178), .B2(n9031), .ZN(
        n6810) );
  INV_X1 U3229 ( .A(n6811), .ZN(n11170) );
  AOI22_X1 U3230 ( .A1(ram[2280]), .A2(n6803), .B1(n11178), .B2(n9055), .ZN(
        n6811) );
  INV_X1 U3231 ( .A(n6812), .ZN(n11171) );
  AOI22_X1 U3232 ( .A1(ram[2281]), .A2(n6803), .B1(n11178), .B2(n9079), .ZN(
        n6812) );
  INV_X1 U3233 ( .A(n6813), .ZN(n11172) );
  AOI22_X1 U3234 ( .A1(ram[2282]), .A2(n6803), .B1(n11178), .B2(n9103), .ZN(
        n6813) );
  INV_X1 U3235 ( .A(n6814), .ZN(n11173) );
  AOI22_X1 U3236 ( .A1(ram[2283]), .A2(n6803), .B1(n11178), .B2(n9127), .ZN(
        n6814) );
  INV_X1 U3237 ( .A(n6815), .ZN(n11174) );
  AOI22_X1 U3238 ( .A1(ram[2284]), .A2(n6803), .B1(n11178), .B2(n9151), .ZN(
        n6815) );
  INV_X1 U3239 ( .A(n6816), .ZN(n11175) );
  AOI22_X1 U3240 ( .A1(ram[2285]), .A2(n6803), .B1(n11178), .B2(n9175), .ZN(
        n6816) );
  INV_X1 U3241 ( .A(n6817), .ZN(n11176) );
  AOI22_X1 U3242 ( .A1(ram[2286]), .A2(n6803), .B1(n11178), .B2(n9199), .ZN(
        n6817) );
  INV_X1 U3243 ( .A(n6818), .ZN(n11177) );
  AOI22_X1 U3244 ( .A1(ram[2287]), .A2(n6803), .B1(n11178), .B2(n9223), .ZN(
        n6818) );
  INV_X1 U3245 ( .A(n6837), .ZN(n11128) );
  AOI22_X1 U3246 ( .A1(ram[2304]), .A2(n6838), .B1(n11144), .B2(n8863), .ZN(
        n6837) );
  INV_X1 U3247 ( .A(n6839), .ZN(n11129) );
  AOI22_X1 U3248 ( .A1(ram[2305]), .A2(n6838), .B1(n11144), .B2(n8887), .ZN(
        n6839) );
  INV_X1 U3249 ( .A(n6840), .ZN(n11130) );
  AOI22_X1 U3250 ( .A1(ram[2306]), .A2(n6838), .B1(n11144), .B2(n8911), .ZN(
        n6840) );
  INV_X1 U3251 ( .A(n6841), .ZN(n11131) );
  AOI22_X1 U3252 ( .A1(ram[2307]), .A2(n6838), .B1(n11144), .B2(n8935), .ZN(
        n6841) );
  INV_X1 U3253 ( .A(n6842), .ZN(n11132) );
  AOI22_X1 U3254 ( .A1(ram[2308]), .A2(n6838), .B1(n11144), .B2(n8959), .ZN(
        n6842) );
  INV_X1 U3255 ( .A(n6843), .ZN(n11133) );
  AOI22_X1 U3256 ( .A1(ram[2309]), .A2(n6838), .B1(n11144), .B2(n8983), .ZN(
        n6843) );
  INV_X1 U3257 ( .A(n6844), .ZN(n11134) );
  AOI22_X1 U3258 ( .A1(ram[2310]), .A2(n6838), .B1(n11144), .B2(n9007), .ZN(
        n6844) );
  INV_X1 U3259 ( .A(n6845), .ZN(n11135) );
  AOI22_X1 U3260 ( .A1(ram[2311]), .A2(n6838), .B1(n11144), .B2(n9031), .ZN(
        n6845) );
  INV_X1 U3261 ( .A(n6846), .ZN(n11136) );
  AOI22_X1 U3262 ( .A1(ram[2312]), .A2(n6838), .B1(n11144), .B2(n9055), .ZN(
        n6846) );
  INV_X1 U3263 ( .A(n6847), .ZN(n11137) );
  AOI22_X1 U3264 ( .A1(ram[2313]), .A2(n6838), .B1(n11144), .B2(n9079), .ZN(
        n6847) );
  INV_X1 U3265 ( .A(n6848), .ZN(n11138) );
  AOI22_X1 U3266 ( .A1(ram[2314]), .A2(n6838), .B1(n11144), .B2(n9103), .ZN(
        n6848) );
  INV_X1 U3267 ( .A(n6849), .ZN(n11139) );
  AOI22_X1 U3268 ( .A1(ram[2315]), .A2(n6838), .B1(n11144), .B2(n9127), .ZN(
        n6849) );
  INV_X1 U3269 ( .A(n6850), .ZN(n11140) );
  AOI22_X1 U3270 ( .A1(ram[2316]), .A2(n6838), .B1(n11144), .B2(n9151), .ZN(
        n6850) );
  INV_X1 U3271 ( .A(n6851), .ZN(n11141) );
  AOI22_X1 U3272 ( .A1(ram[2317]), .A2(n6838), .B1(n11144), .B2(n9175), .ZN(
        n6851) );
  INV_X1 U3273 ( .A(n6852), .ZN(n11142) );
  AOI22_X1 U3274 ( .A1(ram[2318]), .A2(n6838), .B1(n11144), .B2(n9199), .ZN(
        n6852) );
  INV_X1 U3275 ( .A(n6853), .ZN(n11143) );
  AOI22_X1 U3276 ( .A1(ram[2319]), .A2(n6838), .B1(n11144), .B2(n9223), .ZN(
        n6853) );
  INV_X1 U3277 ( .A(n6872), .ZN(n11094) );
  AOI22_X1 U3278 ( .A1(ram[2336]), .A2(n6873), .B1(n11110), .B2(n8863), .ZN(
        n6872) );
  INV_X1 U3279 ( .A(n6874), .ZN(n11095) );
  AOI22_X1 U3280 ( .A1(ram[2337]), .A2(n6873), .B1(n11110), .B2(n8887), .ZN(
        n6874) );
  INV_X1 U3281 ( .A(n6875), .ZN(n11096) );
  AOI22_X1 U3282 ( .A1(ram[2338]), .A2(n6873), .B1(n11110), .B2(n8911), .ZN(
        n6875) );
  INV_X1 U3283 ( .A(n6876), .ZN(n11097) );
  AOI22_X1 U3284 ( .A1(ram[2339]), .A2(n6873), .B1(n11110), .B2(n8935), .ZN(
        n6876) );
  INV_X1 U3285 ( .A(n6877), .ZN(n11098) );
  AOI22_X1 U3286 ( .A1(ram[2340]), .A2(n6873), .B1(n11110), .B2(n8959), .ZN(
        n6877) );
  INV_X1 U3287 ( .A(n6878), .ZN(n11099) );
  AOI22_X1 U3288 ( .A1(ram[2341]), .A2(n6873), .B1(n11110), .B2(n8983), .ZN(
        n6878) );
  INV_X1 U3289 ( .A(n6879), .ZN(n11100) );
  AOI22_X1 U3290 ( .A1(ram[2342]), .A2(n6873), .B1(n11110), .B2(n9007), .ZN(
        n6879) );
  INV_X1 U3291 ( .A(n6880), .ZN(n11101) );
  AOI22_X1 U3292 ( .A1(ram[2343]), .A2(n6873), .B1(n11110), .B2(n9031), .ZN(
        n6880) );
  INV_X1 U3293 ( .A(n6881), .ZN(n11102) );
  AOI22_X1 U3294 ( .A1(ram[2344]), .A2(n6873), .B1(n11110), .B2(n9055), .ZN(
        n6881) );
  INV_X1 U3295 ( .A(n6882), .ZN(n11103) );
  AOI22_X1 U3296 ( .A1(ram[2345]), .A2(n6873), .B1(n11110), .B2(n9079), .ZN(
        n6882) );
  INV_X1 U3297 ( .A(n6883), .ZN(n11104) );
  AOI22_X1 U3298 ( .A1(ram[2346]), .A2(n6873), .B1(n11110), .B2(n9103), .ZN(
        n6883) );
  INV_X1 U3299 ( .A(n6884), .ZN(n11105) );
  AOI22_X1 U3300 ( .A1(ram[2347]), .A2(n6873), .B1(n11110), .B2(n9127), .ZN(
        n6884) );
  INV_X1 U3301 ( .A(n6885), .ZN(n11106) );
  AOI22_X1 U3302 ( .A1(ram[2348]), .A2(n6873), .B1(n11110), .B2(n9151), .ZN(
        n6885) );
  INV_X1 U3303 ( .A(n6886), .ZN(n11107) );
  AOI22_X1 U3304 ( .A1(ram[2349]), .A2(n6873), .B1(n11110), .B2(n9175), .ZN(
        n6886) );
  INV_X1 U3305 ( .A(n6887), .ZN(n11108) );
  AOI22_X1 U3306 ( .A1(ram[2350]), .A2(n6873), .B1(n11110), .B2(n9199), .ZN(
        n6887) );
  INV_X1 U3307 ( .A(n6888), .ZN(n11109) );
  AOI22_X1 U3308 ( .A1(ram[2351]), .A2(n6873), .B1(n11110), .B2(n9223), .ZN(
        n6888) );
  INV_X1 U3309 ( .A(n6906), .ZN(n11060) );
  AOI22_X1 U3310 ( .A1(ram[2368]), .A2(n6907), .B1(n11076), .B2(n8862), .ZN(
        n6906) );
  INV_X1 U3311 ( .A(n6908), .ZN(n11061) );
  AOI22_X1 U3312 ( .A1(ram[2369]), .A2(n6907), .B1(n11076), .B2(n8886), .ZN(
        n6908) );
  INV_X1 U3313 ( .A(n6909), .ZN(n11062) );
  AOI22_X1 U3314 ( .A1(ram[2370]), .A2(n6907), .B1(n11076), .B2(n8910), .ZN(
        n6909) );
  INV_X1 U3315 ( .A(n6910), .ZN(n11063) );
  AOI22_X1 U3316 ( .A1(ram[2371]), .A2(n6907), .B1(n11076), .B2(n8934), .ZN(
        n6910) );
  INV_X1 U3317 ( .A(n6911), .ZN(n11064) );
  AOI22_X1 U3318 ( .A1(ram[2372]), .A2(n6907), .B1(n11076), .B2(n8958), .ZN(
        n6911) );
  INV_X1 U3319 ( .A(n6912), .ZN(n11065) );
  AOI22_X1 U3320 ( .A1(ram[2373]), .A2(n6907), .B1(n11076), .B2(n8982), .ZN(
        n6912) );
  INV_X1 U3321 ( .A(n6913), .ZN(n11066) );
  AOI22_X1 U3322 ( .A1(ram[2374]), .A2(n6907), .B1(n11076), .B2(n9006), .ZN(
        n6913) );
  INV_X1 U3323 ( .A(n6914), .ZN(n11067) );
  AOI22_X1 U3324 ( .A1(ram[2375]), .A2(n6907), .B1(n11076), .B2(n9030), .ZN(
        n6914) );
  INV_X1 U3325 ( .A(n6915), .ZN(n11068) );
  AOI22_X1 U3326 ( .A1(ram[2376]), .A2(n6907), .B1(n11076), .B2(n9054), .ZN(
        n6915) );
  INV_X1 U3327 ( .A(n6916), .ZN(n11069) );
  AOI22_X1 U3328 ( .A1(ram[2377]), .A2(n6907), .B1(n11076), .B2(n9078), .ZN(
        n6916) );
  INV_X1 U3329 ( .A(n6917), .ZN(n11070) );
  AOI22_X1 U3330 ( .A1(ram[2378]), .A2(n6907), .B1(n11076), .B2(n9102), .ZN(
        n6917) );
  INV_X1 U3331 ( .A(n6918), .ZN(n11071) );
  AOI22_X1 U3332 ( .A1(ram[2379]), .A2(n6907), .B1(n11076), .B2(n9126), .ZN(
        n6918) );
  INV_X1 U3333 ( .A(n6919), .ZN(n11072) );
  AOI22_X1 U3334 ( .A1(ram[2380]), .A2(n6907), .B1(n11076), .B2(n9150), .ZN(
        n6919) );
  INV_X1 U3335 ( .A(n6920), .ZN(n11073) );
  AOI22_X1 U3336 ( .A1(ram[2381]), .A2(n6907), .B1(n11076), .B2(n9174), .ZN(
        n6920) );
  INV_X1 U3337 ( .A(n6921), .ZN(n11074) );
  AOI22_X1 U3338 ( .A1(ram[2382]), .A2(n6907), .B1(n11076), .B2(n9198), .ZN(
        n6921) );
  INV_X1 U3339 ( .A(n6922), .ZN(n11075) );
  AOI22_X1 U3340 ( .A1(ram[2383]), .A2(n6907), .B1(n11076), .B2(n9222), .ZN(
        n6922) );
  INV_X1 U3341 ( .A(n6940), .ZN(n11026) );
  AOI22_X1 U3342 ( .A1(ram[2400]), .A2(n6941), .B1(n11042), .B2(n8862), .ZN(
        n6940) );
  INV_X1 U3343 ( .A(n6942), .ZN(n11027) );
  AOI22_X1 U3344 ( .A1(ram[2401]), .A2(n6941), .B1(n11042), .B2(n8886), .ZN(
        n6942) );
  INV_X1 U3345 ( .A(n6943), .ZN(n11028) );
  AOI22_X1 U3346 ( .A1(ram[2402]), .A2(n6941), .B1(n11042), .B2(n8910), .ZN(
        n6943) );
  INV_X1 U3347 ( .A(n6944), .ZN(n11029) );
  AOI22_X1 U3348 ( .A1(ram[2403]), .A2(n6941), .B1(n11042), .B2(n8934), .ZN(
        n6944) );
  INV_X1 U3349 ( .A(n6945), .ZN(n11030) );
  AOI22_X1 U3350 ( .A1(ram[2404]), .A2(n6941), .B1(n11042), .B2(n8958), .ZN(
        n6945) );
  INV_X1 U3351 ( .A(n6946), .ZN(n11031) );
  AOI22_X1 U3352 ( .A1(ram[2405]), .A2(n6941), .B1(n11042), .B2(n8982), .ZN(
        n6946) );
  INV_X1 U3353 ( .A(n6947), .ZN(n11032) );
  AOI22_X1 U3354 ( .A1(ram[2406]), .A2(n6941), .B1(n11042), .B2(n9006), .ZN(
        n6947) );
  INV_X1 U3355 ( .A(n6948), .ZN(n11033) );
  AOI22_X1 U3356 ( .A1(ram[2407]), .A2(n6941), .B1(n11042), .B2(n9030), .ZN(
        n6948) );
  INV_X1 U3357 ( .A(n6949), .ZN(n11034) );
  AOI22_X1 U3358 ( .A1(ram[2408]), .A2(n6941), .B1(n11042), .B2(n9054), .ZN(
        n6949) );
  INV_X1 U3359 ( .A(n6950), .ZN(n11035) );
  AOI22_X1 U3360 ( .A1(ram[2409]), .A2(n6941), .B1(n11042), .B2(n9078), .ZN(
        n6950) );
  INV_X1 U3361 ( .A(n6951), .ZN(n11036) );
  AOI22_X1 U3362 ( .A1(ram[2410]), .A2(n6941), .B1(n11042), .B2(n9102), .ZN(
        n6951) );
  INV_X1 U3363 ( .A(n6952), .ZN(n11037) );
  AOI22_X1 U3364 ( .A1(ram[2411]), .A2(n6941), .B1(n11042), .B2(n9126), .ZN(
        n6952) );
  INV_X1 U3365 ( .A(n6953), .ZN(n11038) );
  AOI22_X1 U3366 ( .A1(ram[2412]), .A2(n6941), .B1(n11042), .B2(n9150), .ZN(
        n6953) );
  INV_X1 U3367 ( .A(n6954), .ZN(n11039) );
  AOI22_X1 U3368 ( .A1(ram[2413]), .A2(n6941), .B1(n11042), .B2(n9174), .ZN(
        n6954) );
  INV_X1 U3369 ( .A(n6955), .ZN(n11040) );
  AOI22_X1 U3370 ( .A1(ram[2414]), .A2(n6941), .B1(n11042), .B2(n9198), .ZN(
        n6955) );
  INV_X1 U3371 ( .A(n6956), .ZN(n11041) );
  AOI22_X1 U3372 ( .A1(ram[2415]), .A2(n6941), .B1(n11042), .B2(n9222), .ZN(
        n6956) );
  INV_X1 U3373 ( .A(n6974), .ZN(n10992) );
  AOI22_X1 U3374 ( .A1(ram[2432]), .A2(n6975), .B1(n11008), .B2(n8862), .ZN(
        n6974) );
  INV_X1 U3375 ( .A(n6976), .ZN(n10993) );
  AOI22_X1 U3376 ( .A1(ram[2433]), .A2(n6975), .B1(n11008), .B2(n8886), .ZN(
        n6976) );
  INV_X1 U3377 ( .A(n6977), .ZN(n10994) );
  AOI22_X1 U3378 ( .A1(ram[2434]), .A2(n6975), .B1(n11008), .B2(n8910), .ZN(
        n6977) );
  INV_X1 U3379 ( .A(n6978), .ZN(n10995) );
  AOI22_X1 U3380 ( .A1(ram[2435]), .A2(n6975), .B1(n11008), .B2(n8934), .ZN(
        n6978) );
  INV_X1 U3381 ( .A(n6979), .ZN(n10996) );
  AOI22_X1 U3382 ( .A1(ram[2436]), .A2(n6975), .B1(n11008), .B2(n8958), .ZN(
        n6979) );
  INV_X1 U3383 ( .A(n6980), .ZN(n10997) );
  AOI22_X1 U3384 ( .A1(ram[2437]), .A2(n6975), .B1(n11008), .B2(n8982), .ZN(
        n6980) );
  INV_X1 U3385 ( .A(n6981), .ZN(n10998) );
  AOI22_X1 U3386 ( .A1(ram[2438]), .A2(n6975), .B1(n11008), .B2(n9006), .ZN(
        n6981) );
  INV_X1 U3387 ( .A(n6982), .ZN(n10999) );
  AOI22_X1 U3388 ( .A1(ram[2439]), .A2(n6975), .B1(n11008), .B2(n9030), .ZN(
        n6982) );
  INV_X1 U3389 ( .A(n6983), .ZN(n11000) );
  AOI22_X1 U3390 ( .A1(ram[2440]), .A2(n6975), .B1(n11008), .B2(n9054), .ZN(
        n6983) );
  INV_X1 U3391 ( .A(n6984), .ZN(n11001) );
  AOI22_X1 U3392 ( .A1(ram[2441]), .A2(n6975), .B1(n11008), .B2(n9078), .ZN(
        n6984) );
  INV_X1 U3393 ( .A(n6985), .ZN(n11002) );
  AOI22_X1 U3394 ( .A1(ram[2442]), .A2(n6975), .B1(n11008), .B2(n9102), .ZN(
        n6985) );
  INV_X1 U3395 ( .A(n6986), .ZN(n11003) );
  AOI22_X1 U3396 ( .A1(ram[2443]), .A2(n6975), .B1(n11008), .B2(n9126), .ZN(
        n6986) );
  INV_X1 U3397 ( .A(n6987), .ZN(n11004) );
  AOI22_X1 U3398 ( .A1(ram[2444]), .A2(n6975), .B1(n11008), .B2(n9150), .ZN(
        n6987) );
  INV_X1 U3399 ( .A(n6988), .ZN(n11005) );
  AOI22_X1 U3400 ( .A1(ram[2445]), .A2(n6975), .B1(n11008), .B2(n9174), .ZN(
        n6988) );
  INV_X1 U3401 ( .A(n6989), .ZN(n11006) );
  AOI22_X1 U3402 ( .A1(ram[2446]), .A2(n6975), .B1(n11008), .B2(n9198), .ZN(
        n6989) );
  INV_X1 U3403 ( .A(n6990), .ZN(n11007) );
  AOI22_X1 U3404 ( .A1(ram[2447]), .A2(n6975), .B1(n11008), .B2(n9222), .ZN(
        n6990) );
  INV_X1 U3405 ( .A(n7008), .ZN(n10958) );
  AOI22_X1 U3406 ( .A1(ram[2464]), .A2(n7009), .B1(n10974), .B2(n8862), .ZN(
        n7008) );
  INV_X1 U3407 ( .A(n7010), .ZN(n10959) );
  AOI22_X1 U3408 ( .A1(ram[2465]), .A2(n7009), .B1(n10974), .B2(n8886), .ZN(
        n7010) );
  INV_X1 U3409 ( .A(n7011), .ZN(n10960) );
  AOI22_X1 U3410 ( .A1(ram[2466]), .A2(n7009), .B1(n10974), .B2(n8910), .ZN(
        n7011) );
  INV_X1 U3411 ( .A(n7012), .ZN(n10961) );
  AOI22_X1 U3412 ( .A1(ram[2467]), .A2(n7009), .B1(n10974), .B2(n8934), .ZN(
        n7012) );
  INV_X1 U3413 ( .A(n7013), .ZN(n10962) );
  AOI22_X1 U3414 ( .A1(ram[2468]), .A2(n7009), .B1(n10974), .B2(n8958), .ZN(
        n7013) );
  INV_X1 U3415 ( .A(n7014), .ZN(n10963) );
  AOI22_X1 U3416 ( .A1(ram[2469]), .A2(n7009), .B1(n10974), .B2(n8982), .ZN(
        n7014) );
  INV_X1 U3417 ( .A(n7015), .ZN(n10964) );
  AOI22_X1 U3418 ( .A1(ram[2470]), .A2(n7009), .B1(n10974), .B2(n9006), .ZN(
        n7015) );
  INV_X1 U3419 ( .A(n7016), .ZN(n10965) );
  AOI22_X1 U3420 ( .A1(ram[2471]), .A2(n7009), .B1(n10974), .B2(n9030), .ZN(
        n7016) );
  INV_X1 U3421 ( .A(n7017), .ZN(n10966) );
  AOI22_X1 U3422 ( .A1(ram[2472]), .A2(n7009), .B1(n10974), .B2(n9054), .ZN(
        n7017) );
  INV_X1 U3423 ( .A(n7018), .ZN(n10967) );
  AOI22_X1 U3424 ( .A1(ram[2473]), .A2(n7009), .B1(n10974), .B2(n9078), .ZN(
        n7018) );
  INV_X1 U3425 ( .A(n7019), .ZN(n10968) );
  AOI22_X1 U3426 ( .A1(ram[2474]), .A2(n7009), .B1(n10974), .B2(n9102), .ZN(
        n7019) );
  INV_X1 U3427 ( .A(n7020), .ZN(n10969) );
  AOI22_X1 U3428 ( .A1(ram[2475]), .A2(n7009), .B1(n10974), .B2(n9126), .ZN(
        n7020) );
  INV_X1 U3429 ( .A(n7021), .ZN(n10970) );
  AOI22_X1 U3430 ( .A1(ram[2476]), .A2(n7009), .B1(n10974), .B2(n9150), .ZN(
        n7021) );
  INV_X1 U3431 ( .A(n7022), .ZN(n10971) );
  AOI22_X1 U3432 ( .A1(ram[2477]), .A2(n7009), .B1(n10974), .B2(n9174), .ZN(
        n7022) );
  INV_X1 U3433 ( .A(n7023), .ZN(n10972) );
  AOI22_X1 U3434 ( .A1(ram[2478]), .A2(n7009), .B1(n10974), .B2(n9198), .ZN(
        n7023) );
  INV_X1 U3435 ( .A(n7024), .ZN(n10973) );
  AOI22_X1 U3436 ( .A1(ram[2479]), .A2(n7009), .B1(n10974), .B2(n9222), .ZN(
        n7024) );
  INV_X1 U3437 ( .A(n7042), .ZN(n10924) );
  AOI22_X1 U3438 ( .A1(ram[2496]), .A2(n7043), .B1(n10940), .B2(n8862), .ZN(
        n7042) );
  INV_X1 U3439 ( .A(n7044), .ZN(n10925) );
  AOI22_X1 U3440 ( .A1(ram[2497]), .A2(n7043), .B1(n10940), .B2(n8886), .ZN(
        n7044) );
  INV_X1 U3441 ( .A(n7045), .ZN(n10926) );
  AOI22_X1 U3442 ( .A1(ram[2498]), .A2(n7043), .B1(n10940), .B2(n8910), .ZN(
        n7045) );
  INV_X1 U3443 ( .A(n7046), .ZN(n10927) );
  AOI22_X1 U3444 ( .A1(ram[2499]), .A2(n7043), .B1(n10940), .B2(n8934), .ZN(
        n7046) );
  INV_X1 U3445 ( .A(n7047), .ZN(n10928) );
  AOI22_X1 U3446 ( .A1(ram[2500]), .A2(n7043), .B1(n10940), .B2(n8958), .ZN(
        n7047) );
  INV_X1 U3447 ( .A(n7048), .ZN(n10929) );
  AOI22_X1 U3448 ( .A1(ram[2501]), .A2(n7043), .B1(n10940), .B2(n8982), .ZN(
        n7048) );
  INV_X1 U3449 ( .A(n7049), .ZN(n10930) );
  AOI22_X1 U3450 ( .A1(ram[2502]), .A2(n7043), .B1(n10940), .B2(n9006), .ZN(
        n7049) );
  INV_X1 U3451 ( .A(n7050), .ZN(n10931) );
  AOI22_X1 U3452 ( .A1(ram[2503]), .A2(n7043), .B1(n10940), .B2(n9030), .ZN(
        n7050) );
  INV_X1 U3453 ( .A(n7051), .ZN(n10932) );
  AOI22_X1 U3454 ( .A1(ram[2504]), .A2(n7043), .B1(n10940), .B2(n9054), .ZN(
        n7051) );
  INV_X1 U3455 ( .A(n7052), .ZN(n10933) );
  AOI22_X1 U3456 ( .A1(ram[2505]), .A2(n7043), .B1(n10940), .B2(n9078), .ZN(
        n7052) );
  INV_X1 U3457 ( .A(n7053), .ZN(n10934) );
  AOI22_X1 U3458 ( .A1(ram[2506]), .A2(n7043), .B1(n10940), .B2(n9102), .ZN(
        n7053) );
  INV_X1 U3459 ( .A(n7054), .ZN(n10935) );
  AOI22_X1 U3460 ( .A1(ram[2507]), .A2(n7043), .B1(n10940), .B2(n9126), .ZN(
        n7054) );
  INV_X1 U3461 ( .A(n7055), .ZN(n10936) );
  AOI22_X1 U3462 ( .A1(ram[2508]), .A2(n7043), .B1(n10940), .B2(n9150), .ZN(
        n7055) );
  INV_X1 U3463 ( .A(n7056), .ZN(n10937) );
  AOI22_X1 U3464 ( .A1(ram[2509]), .A2(n7043), .B1(n10940), .B2(n9174), .ZN(
        n7056) );
  INV_X1 U3465 ( .A(n7057), .ZN(n10938) );
  AOI22_X1 U3466 ( .A1(ram[2510]), .A2(n7043), .B1(n10940), .B2(n9198), .ZN(
        n7057) );
  INV_X1 U3467 ( .A(n7058), .ZN(n10939) );
  AOI22_X1 U3468 ( .A1(ram[2511]), .A2(n7043), .B1(n10940), .B2(n9222), .ZN(
        n7058) );
  INV_X1 U3469 ( .A(n7076), .ZN(n10890) );
  AOI22_X1 U3470 ( .A1(ram[2528]), .A2(n7077), .B1(n10906), .B2(n8862), .ZN(
        n7076) );
  INV_X1 U3471 ( .A(n7078), .ZN(n10891) );
  AOI22_X1 U3472 ( .A1(ram[2529]), .A2(n7077), .B1(n10906), .B2(n8886), .ZN(
        n7078) );
  INV_X1 U3473 ( .A(n7079), .ZN(n10892) );
  AOI22_X1 U3474 ( .A1(ram[2530]), .A2(n7077), .B1(n10906), .B2(n8910), .ZN(
        n7079) );
  INV_X1 U3475 ( .A(n7080), .ZN(n10893) );
  AOI22_X1 U3476 ( .A1(ram[2531]), .A2(n7077), .B1(n10906), .B2(n8934), .ZN(
        n7080) );
  INV_X1 U3477 ( .A(n7081), .ZN(n10894) );
  AOI22_X1 U3478 ( .A1(ram[2532]), .A2(n7077), .B1(n10906), .B2(n8958), .ZN(
        n7081) );
  INV_X1 U3479 ( .A(n7082), .ZN(n10895) );
  AOI22_X1 U3480 ( .A1(ram[2533]), .A2(n7077), .B1(n10906), .B2(n8982), .ZN(
        n7082) );
  INV_X1 U3481 ( .A(n7083), .ZN(n10896) );
  AOI22_X1 U3482 ( .A1(ram[2534]), .A2(n7077), .B1(n10906), .B2(n9006), .ZN(
        n7083) );
  INV_X1 U3483 ( .A(n7084), .ZN(n10897) );
  AOI22_X1 U3484 ( .A1(ram[2535]), .A2(n7077), .B1(n10906), .B2(n9030), .ZN(
        n7084) );
  INV_X1 U3485 ( .A(n7085), .ZN(n10898) );
  AOI22_X1 U3486 ( .A1(ram[2536]), .A2(n7077), .B1(n10906), .B2(n9054), .ZN(
        n7085) );
  INV_X1 U3487 ( .A(n7086), .ZN(n10899) );
  AOI22_X1 U3488 ( .A1(ram[2537]), .A2(n7077), .B1(n10906), .B2(n9078), .ZN(
        n7086) );
  INV_X1 U3489 ( .A(n7087), .ZN(n10900) );
  AOI22_X1 U3490 ( .A1(ram[2538]), .A2(n7077), .B1(n10906), .B2(n9102), .ZN(
        n7087) );
  INV_X1 U3491 ( .A(n7088), .ZN(n10901) );
  AOI22_X1 U3492 ( .A1(ram[2539]), .A2(n7077), .B1(n10906), .B2(n9126), .ZN(
        n7088) );
  INV_X1 U3493 ( .A(n7089), .ZN(n10902) );
  AOI22_X1 U3494 ( .A1(ram[2540]), .A2(n7077), .B1(n10906), .B2(n9150), .ZN(
        n7089) );
  INV_X1 U3495 ( .A(n7090), .ZN(n10903) );
  AOI22_X1 U3496 ( .A1(ram[2541]), .A2(n7077), .B1(n10906), .B2(n9174), .ZN(
        n7090) );
  INV_X1 U3497 ( .A(n7091), .ZN(n10904) );
  AOI22_X1 U3498 ( .A1(ram[2542]), .A2(n7077), .B1(n10906), .B2(n9198), .ZN(
        n7091) );
  INV_X1 U3499 ( .A(n7092), .ZN(n10905) );
  AOI22_X1 U3500 ( .A1(ram[2543]), .A2(n7077), .B1(n10906), .B2(n9222), .ZN(
        n7092) );
  INV_X1 U3501 ( .A(n7110), .ZN(n10856) );
  AOI22_X1 U3502 ( .A1(ram[2560]), .A2(n7111), .B1(n10872), .B2(n8861), .ZN(
        n7110) );
  INV_X1 U3503 ( .A(n7112), .ZN(n10857) );
  AOI22_X1 U3504 ( .A1(ram[2561]), .A2(n7111), .B1(n10872), .B2(n8885), .ZN(
        n7112) );
  INV_X1 U3505 ( .A(n7113), .ZN(n10858) );
  AOI22_X1 U3506 ( .A1(ram[2562]), .A2(n7111), .B1(n10872), .B2(n8909), .ZN(
        n7113) );
  INV_X1 U3507 ( .A(n7114), .ZN(n10859) );
  AOI22_X1 U3508 ( .A1(ram[2563]), .A2(n7111), .B1(n10872), .B2(n8933), .ZN(
        n7114) );
  INV_X1 U3509 ( .A(n7115), .ZN(n10860) );
  AOI22_X1 U3510 ( .A1(ram[2564]), .A2(n7111), .B1(n10872), .B2(n8957), .ZN(
        n7115) );
  INV_X1 U3511 ( .A(n7116), .ZN(n10861) );
  AOI22_X1 U3512 ( .A1(ram[2565]), .A2(n7111), .B1(n10872), .B2(n8981), .ZN(
        n7116) );
  INV_X1 U3513 ( .A(n7117), .ZN(n10862) );
  AOI22_X1 U3514 ( .A1(ram[2566]), .A2(n7111), .B1(n10872), .B2(n9005), .ZN(
        n7117) );
  INV_X1 U3515 ( .A(n7118), .ZN(n10863) );
  AOI22_X1 U3516 ( .A1(ram[2567]), .A2(n7111), .B1(n10872), .B2(n9029), .ZN(
        n7118) );
  INV_X1 U3517 ( .A(n7119), .ZN(n10864) );
  AOI22_X1 U3518 ( .A1(ram[2568]), .A2(n7111), .B1(n10872), .B2(n9053), .ZN(
        n7119) );
  INV_X1 U3519 ( .A(n7120), .ZN(n10865) );
  AOI22_X1 U3520 ( .A1(ram[2569]), .A2(n7111), .B1(n10872), .B2(n9077), .ZN(
        n7120) );
  INV_X1 U3521 ( .A(n7121), .ZN(n10866) );
  AOI22_X1 U3522 ( .A1(ram[2570]), .A2(n7111), .B1(n10872), .B2(n9101), .ZN(
        n7121) );
  INV_X1 U3523 ( .A(n7122), .ZN(n10867) );
  AOI22_X1 U3524 ( .A1(ram[2571]), .A2(n7111), .B1(n10872), .B2(n9125), .ZN(
        n7122) );
  INV_X1 U3525 ( .A(n7123), .ZN(n10868) );
  AOI22_X1 U3526 ( .A1(ram[2572]), .A2(n7111), .B1(n10872), .B2(n9149), .ZN(
        n7123) );
  INV_X1 U3527 ( .A(n7124), .ZN(n10869) );
  AOI22_X1 U3528 ( .A1(ram[2573]), .A2(n7111), .B1(n10872), .B2(n9173), .ZN(
        n7124) );
  INV_X1 U3529 ( .A(n7125), .ZN(n10870) );
  AOI22_X1 U3530 ( .A1(ram[2574]), .A2(n7111), .B1(n10872), .B2(n9197), .ZN(
        n7125) );
  INV_X1 U3531 ( .A(n7126), .ZN(n10871) );
  AOI22_X1 U3532 ( .A1(ram[2575]), .A2(n7111), .B1(n10872), .B2(n9221), .ZN(
        n7126) );
  INV_X1 U3533 ( .A(n7145), .ZN(n10822) );
  AOI22_X1 U3534 ( .A1(ram[2592]), .A2(n7146), .B1(n10838), .B2(n8861), .ZN(
        n7145) );
  INV_X1 U3535 ( .A(n7147), .ZN(n10823) );
  AOI22_X1 U3536 ( .A1(ram[2593]), .A2(n7146), .B1(n10838), .B2(n8885), .ZN(
        n7147) );
  INV_X1 U3537 ( .A(n7148), .ZN(n10824) );
  AOI22_X1 U3538 ( .A1(ram[2594]), .A2(n7146), .B1(n10838), .B2(n8909), .ZN(
        n7148) );
  INV_X1 U3539 ( .A(n7149), .ZN(n10825) );
  AOI22_X1 U3540 ( .A1(ram[2595]), .A2(n7146), .B1(n10838), .B2(n8933), .ZN(
        n7149) );
  INV_X1 U3541 ( .A(n7150), .ZN(n10826) );
  AOI22_X1 U3542 ( .A1(ram[2596]), .A2(n7146), .B1(n10838), .B2(n8957), .ZN(
        n7150) );
  INV_X1 U3543 ( .A(n7151), .ZN(n10827) );
  AOI22_X1 U3544 ( .A1(ram[2597]), .A2(n7146), .B1(n10838), .B2(n8981), .ZN(
        n7151) );
  INV_X1 U3545 ( .A(n7152), .ZN(n10828) );
  AOI22_X1 U3546 ( .A1(ram[2598]), .A2(n7146), .B1(n10838), .B2(n9005), .ZN(
        n7152) );
  INV_X1 U3547 ( .A(n7153), .ZN(n10829) );
  AOI22_X1 U3548 ( .A1(ram[2599]), .A2(n7146), .B1(n10838), .B2(n9029), .ZN(
        n7153) );
  INV_X1 U3549 ( .A(n7154), .ZN(n10830) );
  AOI22_X1 U3550 ( .A1(ram[2600]), .A2(n7146), .B1(n10838), .B2(n9053), .ZN(
        n7154) );
  INV_X1 U3551 ( .A(n7155), .ZN(n10831) );
  AOI22_X1 U3552 ( .A1(ram[2601]), .A2(n7146), .B1(n10838), .B2(n9077), .ZN(
        n7155) );
  INV_X1 U3553 ( .A(n7156), .ZN(n10832) );
  AOI22_X1 U3554 ( .A1(ram[2602]), .A2(n7146), .B1(n10838), .B2(n9101), .ZN(
        n7156) );
  INV_X1 U3555 ( .A(n7157), .ZN(n10833) );
  AOI22_X1 U3556 ( .A1(ram[2603]), .A2(n7146), .B1(n10838), .B2(n9125), .ZN(
        n7157) );
  INV_X1 U3557 ( .A(n7158), .ZN(n10834) );
  AOI22_X1 U3558 ( .A1(ram[2604]), .A2(n7146), .B1(n10838), .B2(n9149), .ZN(
        n7158) );
  INV_X1 U3559 ( .A(n7159), .ZN(n10835) );
  AOI22_X1 U3560 ( .A1(ram[2605]), .A2(n7146), .B1(n10838), .B2(n9173), .ZN(
        n7159) );
  INV_X1 U3561 ( .A(n7160), .ZN(n10836) );
  AOI22_X1 U3562 ( .A1(ram[2606]), .A2(n7146), .B1(n10838), .B2(n9197), .ZN(
        n7160) );
  INV_X1 U3563 ( .A(n7161), .ZN(n10837) );
  AOI22_X1 U3564 ( .A1(ram[2607]), .A2(n7146), .B1(n10838), .B2(n9221), .ZN(
        n7161) );
  INV_X1 U3565 ( .A(n7179), .ZN(n10788) );
  AOI22_X1 U3566 ( .A1(ram[2624]), .A2(n7180), .B1(n10804), .B2(n8861), .ZN(
        n7179) );
  INV_X1 U3567 ( .A(n7181), .ZN(n10789) );
  AOI22_X1 U3568 ( .A1(ram[2625]), .A2(n7180), .B1(n10804), .B2(n8885), .ZN(
        n7181) );
  INV_X1 U3569 ( .A(n7182), .ZN(n10790) );
  AOI22_X1 U3570 ( .A1(ram[2626]), .A2(n7180), .B1(n10804), .B2(n8909), .ZN(
        n7182) );
  INV_X1 U3571 ( .A(n7183), .ZN(n10791) );
  AOI22_X1 U3572 ( .A1(ram[2627]), .A2(n7180), .B1(n10804), .B2(n8933), .ZN(
        n7183) );
  INV_X1 U3573 ( .A(n7184), .ZN(n10792) );
  AOI22_X1 U3574 ( .A1(ram[2628]), .A2(n7180), .B1(n10804), .B2(n8957), .ZN(
        n7184) );
  INV_X1 U3575 ( .A(n7185), .ZN(n10793) );
  AOI22_X1 U3576 ( .A1(ram[2629]), .A2(n7180), .B1(n10804), .B2(n8981), .ZN(
        n7185) );
  INV_X1 U3577 ( .A(n7186), .ZN(n10794) );
  AOI22_X1 U3578 ( .A1(ram[2630]), .A2(n7180), .B1(n10804), .B2(n9005), .ZN(
        n7186) );
  INV_X1 U3579 ( .A(n7187), .ZN(n10795) );
  AOI22_X1 U3580 ( .A1(ram[2631]), .A2(n7180), .B1(n10804), .B2(n9029), .ZN(
        n7187) );
  INV_X1 U3581 ( .A(n7188), .ZN(n10796) );
  AOI22_X1 U3582 ( .A1(ram[2632]), .A2(n7180), .B1(n10804), .B2(n9053), .ZN(
        n7188) );
  INV_X1 U3583 ( .A(n7189), .ZN(n10797) );
  AOI22_X1 U3584 ( .A1(ram[2633]), .A2(n7180), .B1(n10804), .B2(n9077), .ZN(
        n7189) );
  INV_X1 U3585 ( .A(n7190), .ZN(n10798) );
  AOI22_X1 U3586 ( .A1(ram[2634]), .A2(n7180), .B1(n10804), .B2(n9101), .ZN(
        n7190) );
  INV_X1 U3587 ( .A(n7191), .ZN(n10799) );
  AOI22_X1 U3588 ( .A1(ram[2635]), .A2(n7180), .B1(n10804), .B2(n9125), .ZN(
        n7191) );
  INV_X1 U3589 ( .A(n7192), .ZN(n10800) );
  AOI22_X1 U3590 ( .A1(ram[2636]), .A2(n7180), .B1(n10804), .B2(n9149), .ZN(
        n7192) );
  INV_X1 U3591 ( .A(n7193), .ZN(n10801) );
  AOI22_X1 U3592 ( .A1(ram[2637]), .A2(n7180), .B1(n10804), .B2(n9173), .ZN(
        n7193) );
  INV_X1 U3593 ( .A(n7194), .ZN(n10802) );
  AOI22_X1 U3594 ( .A1(ram[2638]), .A2(n7180), .B1(n10804), .B2(n9197), .ZN(
        n7194) );
  INV_X1 U3595 ( .A(n7195), .ZN(n10803) );
  AOI22_X1 U3596 ( .A1(ram[2639]), .A2(n7180), .B1(n10804), .B2(n9221), .ZN(
        n7195) );
  INV_X1 U3597 ( .A(n7213), .ZN(n10754) );
  AOI22_X1 U3598 ( .A1(ram[2656]), .A2(n7214), .B1(n10770), .B2(n8861), .ZN(
        n7213) );
  INV_X1 U3599 ( .A(n7215), .ZN(n10755) );
  AOI22_X1 U3600 ( .A1(ram[2657]), .A2(n7214), .B1(n10770), .B2(n8885), .ZN(
        n7215) );
  INV_X1 U3601 ( .A(n7216), .ZN(n10756) );
  AOI22_X1 U3602 ( .A1(ram[2658]), .A2(n7214), .B1(n10770), .B2(n8909), .ZN(
        n7216) );
  INV_X1 U3603 ( .A(n7217), .ZN(n10757) );
  AOI22_X1 U3604 ( .A1(ram[2659]), .A2(n7214), .B1(n10770), .B2(n8933), .ZN(
        n7217) );
  INV_X1 U3605 ( .A(n7218), .ZN(n10758) );
  AOI22_X1 U3606 ( .A1(ram[2660]), .A2(n7214), .B1(n10770), .B2(n8957), .ZN(
        n7218) );
  INV_X1 U3607 ( .A(n7219), .ZN(n10759) );
  AOI22_X1 U3608 ( .A1(ram[2661]), .A2(n7214), .B1(n10770), .B2(n8981), .ZN(
        n7219) );
  INV_X1 U3609 ( .A(n7220), .ZN(n10760) );
  AOI22_X1 U3610 ( .A1(ram[2662]), .A2(n7214), .B1(n10770), .B2(n9005), .ZN(
        n7220) );
  INV_X1 U3611 ( .A(n7221), .ZN(n10761) );
  AOI22_X1 U3612 ( .A1(ram[2663]), .A2(n7214), .B1(n10770), .B2(n9029), .ZN(
        n7221) );
  INV_X1 U3613 ( .A(n7222), .ZN(n10762) );
  AOI22_X1 U3614 ( .A1(ram[2664]), .A2(n7214), .B1(n10770), .B2(n9053), .ZN(
        n7222) );
  INV_X1 U3615 ( .A(n7223), .ZN(n10763) );
  AOI22_X1 U3616 ( .A1(ram[2665]), .A2(n7214), .B1(n10770), .B2(n9077), .ZN(
        n7223) );
  INV_X1 U3617 ( .A(n7224), .ZN(n10764) );
  AOI22_X1 U3618 ( .A1(ram[2666]), .A2(n7214), .B1(n10770), .B2(n9101), .ZN(
        n7224) );
  INV_X1 U3619 ( .A(n7225), .ZN(n10765) );
  AOI22_X1 U3620 ( .A1(ram[2667]), .A2(n7214), .B1(n10770), .B2(n9125), .ZN(
        n7225) );
  INV_X1 U3621 ( .A(n7226), .ZN(n10766) );
  AOI22_X1 U3622 ( .A1(ram[2668]), .A2(n7214), .B1(n10770), .B2(n9149), .ZN(
        n7226) );
  INV_X1 U3623 ( .A(n7227), .ZN(n10767) );
  AOI22_X1 U3624 ( .A1(ram[2669]), .A2(n7214), .B1(n10770), .B2(n9173), .ZN(
        n7227) );
  INV_X1 U3625 ( .A(n7228), .ZN(n10768) );
  AOI22_X1 U3626 ( .A1(ram[2670]), .A2(n7214), .B1(n10770), .B2(n9197), .ZN(
        n7228) );
  INV_X1 U3627 ( .A(n7229), .ZN(n10769) );
  AOI22_X1 U3628 ( .A1(ram[2671]), .A2(n7214), .B1(n10770), .B2(n9221), .ZN(
        n7229) );
  INV_X1 U3629 ( .A(n7247), .ZN(n10720) );
  AOI22_X1 U3630 ( .A1(ram[2688]), .A2(n7248), .B1(n10736), .B2(n8861), .ZN(
        n7247) );
  INV_X1 U3631 ( .A(n7249), .ZN(n10721) );
  AOI22_X1 U3632 ( .A1(ram[2689]), .A2(n7248), .B1(n10736), .B2(n8885), .ZN(
        n7249) );
  INV_X1 U3633 ( .A(n7250), .ZN(n10722) );
  AOI22_X1 U3634 ( .A1(ram[2690]), .A2(n7248), .B1(n10736), .B2(n8909), .ZN(
        n7250) );
  INV_X1 U3635 ( .A(n7251), .ZN(n10723) );
  AOI22_X1 U3636 ( .A1(ram[2691]), .A2(n7248), .B1(n10736), .B2(n8933), .ZN(
        n7251) );
  INV_X1 U3637 ( .A(n7252), .ZN(n10724) );
  AOI22_X1 U3638 ( .A1(ram[2692]), .A2(n7248), .B1(n10736), .B2(n8957), .ZN(
        n7252) );
  INV_X1 U3639 ( .A(n7253), .ZN(n10725) );
  AOI22_X1 U3640 ( .A1(ram[2693]), .A2(n7248), .B1(n10736), .B2(n8981), .ZN(
        n7253) );
  INV_X1 U3641 ( .A(n7254), .ZN(n10726) );
  AOI22_X1 U3642 ( .A1(ram[2694]), .A2(n7248), .B1(n10736), .B2(n9005), .ZN(
        n7254) );
  INV_X1 U3643 ( .A(n7255), .ZN(n10727) );
  AOI22_X1 U3644 ( .A1(ram[2695]), .A2(n7248), .B1(n10736), .B2(n9029), .ZN(
        n7255) );
  INV_X1 U3645 ( .A(n7256), .ZN(n10728) );
  AOI22_X1 U3646 ( .A1(ram[2696]), .A2(n7248), .B1(n10736), .B2(n9053), .ZN(
        n7256) );
  INV_X1 U3647 ( .A(n7257), .ZN(n10729) );
  AOI22_X1 U3648 ( .A1(ram[2697]), .A2(n7248), .B1(n10736), .B2(n9077), .ZN(
        n7257) );
  INV_X1 U3649 ( .A(n7258), .ZN(n10730) );
  AOI22_X1 U3650 ( .A1(ram[2698]), .A2(n7248), .B1(n10736), .B2(n9101), .ZN(
        n7258) );
  INV_X1 U3651 ( .A(n7259), .ZN(n10731) );
  AOI22_X1 U3652 ( .A1(ram[2699]), .A2(n7248), .B1(n10736), .B2(n9125), .ZN(
        n7259) );
  INV_X1 U3653 ( .A(n7260), .ZN(n10732) );
  AOI22_X1 U3654 ( .A1(ram[2700]), .A2(n7248), .B1(n10736), .B2(n9149), .ZN(
        n7260) );
  INV_X1 U3655 ( .A(n7261), .ZN(n10733) );
  AOI22_X1 U3656 ( .A1(ram[2701]), .A2(n7248), .B1(n10736), .B2(n9173), .ZN(
        n7261) );
  INV_X1 U3657 ( .A(n7262), .ZN(n10734) );
  AOI22_X1 U3658 ( .A1(ram[2702]), .A2(n7248), .B1(n10736), .B2(n9197), .ZN(
        n7262) );
  INV_X1 U3659 ( .A(n7263), .ZN(n10735) );
  AOI22_X1 U3660 ( .A1(ram[2703]), .A2(n7248), .B1(n10736), .B2(n9221), .ZN(
        n7263) );
  INV_X1 U3661 ( .A(n7281), .ZN(n10686) );
  AOI22_X1 U3662 ( .A1(ram[2720]), .A2(n7282), .B1(n10702), .B2(n8861), .ZN(
        n7281) );
  INV_X1 U3663 ( .A(n7283), .ZN(n10687) );
  AOI22_X1 U3664 ( .A1(ram[2721]), .A2(n7282), .B1(n10702), .B2(n8885), .ZN(
        n7283) );
  INV_X1 U3665 ( .A(n7284), .ZN(n10688) );
  AOI22_X1 U3666 ( .A1(ram[2722]), .A2(n7282), .B1(n10702), .B2(n8909), .ZN(
        n7284) );
  INV_X1 U3667 ( .A(n7285), .ZN(n10689) );
  AOI22_X1 U3668 ( .A1(ram[2723]), .A2(n7282), .B1(n10702), .B2(n8933), .ZN(
        n7285) );
  INV_X1 U3669 ( .A(n7286), .ZN(n10690) );
  AOI22_X1 U3670 ( .A1(ram[2724]), .A2(n7282), .B1(n10702), .B2(n8957), .ZN(
        n7286) );
  INV_X1 U3671 ( .A(n7287), .ZN(n10691) );
  AOI22_X1 U3672 ( .A1(ram[2725]), .A2(n7282), .B1(n10702), .B2(n8981), .ZN(
        n7287) );
  INV_X1 U3673 ( .A(n7288), .ZN(n10692) );
  AOI22_X1 U3674 ( .A1(ram[2726]), .A2(n7282), .B1(n10702), .B2(n9005), .ZN(
        n7288) );
  INV_X1 U3675 ( .A(n7289), .ZN(n10693) );
  AOI22_X1 U3676 ( .A1(ram[2727]), .A2(n7282), .B1(n10702), .B2(n9029), .ZN(
        n7289) );
  INV_X1 U3677 ( .A(n7290), .ZN(n10694) );
  AOI22_X1 U3678 ( .A1(ram[2728]), .A2(n7282), .B1(n10702), .B2(n9053), .ZN(
        n7290) );
  INV_X1 U3679 ( .A(n7291), .ZN(n10695) );
  AOI22_X1 U3680 ( .A1(ram[2729]), .A2(n7282), .B1(n10702), .B2(n9077), .ZN(
        n7291) );
  INV_X1 U3681 ( .A(n7292), .ZN(n10696) );
  AOI22_X1 U3682 ( .A1(ram[2730]), .A2(n7282), .B1(n10702), .B2(n9101), .ZN(
        n7292) );
  INV_X1 U3683 ( .A(n7293), .ZN(n10697) );
  AOI22_X1 U3684 ( .A1(ram[2731]), .A2(n7282), .B1(n10702), .B2(n9125), .ZN(
        n7293) );
  INV_X1 U3685 ( .A(n7294), .ZN(n10698) );
  AOI22_X1 U3686 ( .A1(ram[2732]), .A2(n7282), .B1(n10702), .B2(n9149), .ZN(
        n7294) );
  INV_X1 U3687 ( .A(n7295), .ZN(n10699) );
  AOI22_X1 U3688 ( .A1(ram[2733]), .A2(n7282), .B1(n10702), .B2(n9173), .ZN(
        n7295) );
  INV_X1 U3689 ( .A(n7296), .ZN(n10700) );
  AOI22_X1 U3690 ( .A1(ram[2734]), .A2(n7282), .B1(n10702), .B2(n9197), .ZN(
        n7296) );
  INV_X1 U3691 ( .A(n7297), .ZN(n10701) );
  AOI22_X1 U3692 ( .A1(ram[2735]), .A2(n7282), .B1(n10702), .B2(n9221), .ZN(
        n7297) );
  INV_X1 U3693 ( .A(n7315), .ZN(n10652) );
  AOI22_X1 U3694 ( .A1(ram[2752]), .A2(n7316), .B1(n10668), .B2(n8860), .ZN(
        n7315) );
  INV_X1 U3695 ( .A(n7317), .ZN(n10653) );
  AOI22_X1 U3696 ( .A1(ram[2753]), .A2(n7316), .B1(n10668), .B2(n8884), .ZN(
        n7317) );
  INV_X1 U3697 ( .A(n7318), .ZN(n10654) );
  AOI22_X1 U3698 ( .A1(ram[2754]), .A2(n7316), .B1(n10668), .B2(n8908), .ZN(
        n7318) );
  INV_X1 U3699 ( .A(n7319), .ZN(n10655) );
  AOI22_X1 U3700 ( .A1(ram[2755]), .A2(n7316), .B1(n10668), .B2(n8932), .ZN(
        n7319) );
  INV_X1 U3701 ( .A(n7320), .ZN(n10656) );
  AOI22_X1 U3702 ( .A1(ram[2756]), .A2(n7316), .B1(n10668), .B2(n8956), .ZN(
        n7320) );
  INV_X1 U3703 ( .A(n7321), .ZN(n10657) );
  AOI22_X1 U3704 ( .A1(ram[2757]), .A2(n7316), .B1(n10668), .B2(n8980), .ZN(
        n7321) );
  INV_X1 U3705 ( .A(n7322), .ZN(n10658) );
  AOI22_X1 U3706 ( .A1(ram[2758]), .A2(n7316), .B1(n10668), .B2(n9004), .ZN(
        n7322) );
  INV_X1 U3707 ( .A(n7323), .ZN(n10659) );
  AOI22_X1 U3708 ( .A1(ram[2759]), .A2(n7316), .B1(n10668), .B2(n9028), .ZN(
        n7323) );
  INV_X1 U3709 ( .A(n7324), .ZN(n10660) );
  AOI22_X1 U3710 ( .A1(ram[2760]), .A2(n7316), .B1(n10668), .B2(n9052), .ZN(
        n7324) );
  INV_X1 U3711 ( .A(n7325), .ZN(n10661) );
  AOI22_X1 U3712 ( .A1(ram[2761]), .A2(n7316), .B1(n10668), .B2(n9076), .ZN(
        n7325) );
  INV_X1 U3713 ( .A(n7326), .ZN(n10662) );
  AOI22_X1 U3714 ( .A1(ram[2762]), .A2(n7316), .B1(n10668), .B2(n9100), .ZN(
        n7326) );
  INV_X1 U3715 ( .A(n7327), .ZN(n10663) );
  AOI22_X1 U3716 ( .A1(ram[2763]), .A2(n7316), .B1(n10668), .B2(n9124), .ZN(
        n7327) );
  INV_X1 U3717 ( .A(n7328), .ZN(n10664) );
  AOI22_X1 U3718 ( .A1(ram[2764]), .A2(n7316), .B1(n10668), .B2(n9148), .ZN(
        n7328) );
  INV_X1 U3719 ( .A(n7329), .ZN(n10665) );
  AOI22_X1 U3720 ( .A1(ram[2765]), .A2(n7316), .B1(n10668), .B2(n9172), .ZN(
        n7329) );
  INV_X1 U3721 ( .A(n7330), .ZN(n10666) );
  AOI22_X1 U3722 ( .A1(ram[2766]), .A2(n7316), .B1(n10668), .B2(n9196), .ZN(
        n7330) );
  INV_X1 U3723 ( .A(n7331), .ZN(n10667) );
  AOI22_X1 U3724 ( .A1(ram[2767]), .A2(n7316), .B1(n10668), .B2(n9220), .ZN(
        n7331) );
  INV_X1 U3725 ( .A(n7349), .ZN(n10618) );
  AOI22_X1 U3726 ( .A1(ram[2784]), .A2(n7350), .B1(n10634), .B2(n8860), .ZN(
        n7349) );
  INV_X1 U3727 ( .A(n7351), .ZN(n10619) );
  AOI22_X1 U3728 ( .A1(ram[2785]), .A2(n7350), .B1(n10634), .B2(n8884), .ZN(
        n7351) );
  INV_X1 U3729 ( .A(n7352), .ZN(n10620) );
  AOI22_X1 U3730 ( .A1(ram[2786]), .A2(n7350), .B1(n10634), .B2(n8908), .ZN(
        n7352) );
  INV_X1 U3731 ( .A(n7353), .ZN(n10621) );
  AOI22_X1 U3732 ( .A1(ram[2787]), .A2(n7350), .B1(n10634), .B2(n8932), .ZN(
        n7353) );
  INV_X1 U3733 ( .A(n7354), .ZN(n10622) );
  AOI22_X1 U3734 ( .A1(ram[2788]), .A2(n7350), .B1(n10634), .B2(n8956), .ZN(
        n7354) );
  INV_X1 U3735 ( .A(n7355), .ZN(n10623) );
  AOI22_X1 U3736 ( .A1(ram[2789]), .A2(n7350), .B1(n10634), .B2(n8980), .ZN(
        n7355) );
  INV_X1 U3737 ( .A(n7356), .ZN(n10624) );
  AOI22_X1 U3738 ( .A1(ram[2790]), .A2(n7350), .B1(n10634), .B2(n9004), .ZN(
        n7356) );
  INV_X1 U3739 ( .A(n7357), .ZN(n10625) );
  AOI22_X1 U3740 ( .A1(ram[2791]), .A2(n7350), .B1(n10634), .B2(n9028), .ZN(
        n7357) );
  INV_X1 U3741 ( .A(n7358), .ZN(n10626) );
  AOI22_X1 U3742 ( .A1(ram[2792]), .A2(n7350), .B1(n10634), .B2(n9052), .ZN(
        n7358) );
  INV_X1 U3743 ( .A(n7359), .ZN(n10627) );
  AOI22_X1 U3744 ( .A1(ram[2793]), .A2(n7350), .B1(n10634), .B2(n9076), .ZN(
        n7359) );
  INV_X1 U3745 ( .A(n7360), .ZN(n10628) );
  AOI22_X1 U3746 ( .A1(ram[2794]), .A2(n7350), .B1(n10634), .B2(n9100), .ZN(
        n7360) );
  INV_X1 U3747 ( .A(n7361), .ZN(n10629) );
  AOI22_X1 U3748 ( .A1(ram[2795]), .A2(n7350), .B1(n10634), .B2(n9124), .ZN(
        n7361) );
  INV_X1 U3749 ( .A(n7362), .ZN(n10630) );
  AOI22_X1 U3750 ( .A1(ram[2796]), .A2(n7350), .B1(n10634), .B2(n9148), .ZN(
        n7362) );
  INV_X1 U3751 ( .A(n7363), .ZN(n10631) );
  AOI22_X1 U3752 ( .A1(ram[2797]), .A2(n7350), .B1(n10634), .B2(n9172), .ZN(
        n7363) );
  INV_X1 U3753 ( .A(n7364), .ZN(n10632) );
  AOI22_X1 U3754 ( .A1(ram[2798]), .A2(n7350), .B1(n10634), .B2(n9196), .ZN(
        n7364) );
  INV_X1 U3755 ( .A(n7365), .ZN(n10633) );
  AOI22_X1 U3756 ( .A1(ram[2799]), .A2(n7350), .B1(n10634), .B2(n9220), .ZN(
        n7365) );
  INV_X1 U3757 ( .A(n7383), .ZN(n10584) );
  AOI22_X1 U3758 ( .A1(ram[2816]), .A2(n7384), .B1(n10600), .B2(n8860), .ZN(
        n7383) );
  INV_X1 U3759 ( .A(n7385), .ZN(n10585) );
  AOI22_X1 U3760 ( .A1(ram[2817]), .A2(n7384), .B1(n10600), .B2(n8884), .ZN(
        n7385) );
  INV_X1 U3761 ( .A(n7386), .ZN(n10586) );
  AOI22_X1 U3762 ( .A1(ram[2818]), .A2(n7384), .B1(n10600), .B2(n8908), .ZN(
        n7386) );
  INV_X1 U3763 ( .A(n7387), .ZN(n10587) );
  AOI22_X1 U3764 ( .A1(ram[2819]), .A2(n7384), .B1(n10600), .B2(n8932), .ZN(
        n7387) );
  INV_X1 U3765 ( .A(n7388), .ZN(n10588) );
  AOI22_X1 U3766 ( .A1(ram[2820]), .A2(n7384), .B1(n10600), .B2(n8956), .ZN(
        n7388) );
  INV_X1 U3767 ( .A(n7389), .ZN(n10589) );
  AOI22_X1 U3768 ( .A1(ram[2821]), .A2(n7384), .B1(n10600), .B2(n8980), .ZN(
        n7389) );
  INV_X1 U3769 ( .A(n7390), .ZN(n10590) );
  AOI22_X1 U3770 ( .A1(ram[2822]), .A2(n7384), .B1(n10600), .B2(n9004), .ZN(
        n7390) );
  INV_X1 U3771 ( .A(n7391), .ZN(n10591) );
  AOI22_X1 U3772 ( .A1(ram[2823]), .A2(n7384), .B1(n10600), .B2(n9028), .ZN(
        n7391) );
  INV_X1 U3773 ( .A(n7392), .ZN(n10592) );
  AOI22_X1 U3774 ( .A1(ram[2824]), .A2(n7384), .B1(n10600), .B2(n9052), .ZN(
        n7392) );
  INV_X1 U3775 ( .A(n7393), .ZN(n10593) );
  AOI22_X1 U3776 ( .A1(ram[2825]), .A2(n7384), .B1(n10600), .B2(n9076), .ZN(
        n7393) );
  INV_X1 U3777 ( .A(n7394), .ZN(n10594) );
  AOI22_X1 U3778 ( .A1(ram[2826]), .A2(n7384), .B1(n10600), .B2(n9100), .ZN(
        n7394) );
  INV_X1 U3779 ( .A(n7395), .ZN(n10595) );
  AOI22_X1 U3780 ( .A1(ram[2827]), .A2(n7384), .B1(n10600), .B2(n9124), .ZN(
        n7395) );
  INV_X1 U3781 ( .A(n7396), .ZN(n10596) );
  AOI22_X1 U3782 ( .A1(ram[2828]), .A2(n7384), .B1(n10600), .B2(n9148), .ZN(
        n7396) );
  INV_X1 U3783 ( .A(n7397), .ZN(n10597) );
  AOI22_X1 U3784 ( .A1(ram[2829]), .A2(n7384), .B1(n10600), .B2(n9172), .ZN(
        n7397) );
  INV_X1 U3785 ( .A(n7398), .ZN(n10598) );
  AOI22_X1 U3786 ( .A1(ram[2830]), .A2(n7384), .B1(n10600), .B2(n9196), .ZN(
        n7398) );
  INV_X1 U3787 ( .A(n7399), .ZN(n10599) );
  AOI22_X1 U3788 ( .A1(ram[2831]), .A2(n7384), .B1(n10600), .B2(n9220), .ZN(
        n7399) );
  INV_X1 U3789 ( .A(n7418), .ZN(n10550) );
  AOI22_X1 U3790 ( .A1(ram[2848]), .A2(n7419), .B1(n10566), .B2(n8860), .ZN(
        n7418) );
  INV_X1 U3791 ( .A(n7420), .ZN(n10551) );
  AOI22_X1 U3792 ( .A1(ram[2849]), .A2(n7419), .B1(n10566), .B2(n8884), .ZN(
        n7420) );
  INV_X1 U3793 ( .A(n7421), .ZN(n10552) );
  AOI22_X1 U3794 ( .A1(ram[2850]), .A2(n7419), .B1(n10566), .B2(n8908), .ZN(
        n7421) );
  INV_X1 U3795 ( .A(n7422), .ZN(n10553) );
  AOI22_X1 U3796 ( .A1(ram[2851]), .A2(n7419), .B1(n10566), .B2(n8932), .ZN(
        n7422) );
  INV_X1 U3797 ( .A(n7423), .ZN(n10554) );
  AOI22_X1 U3798 ( .A1(ram[2852]), .A2(n7419), .B1(n10566), .B2(n8956), .ZN(
        n7423) );
  INV_X1 U3799 ( .A(n7424), .ZN(n10555) );
  AOI22_X1 U3800 ( .A1(ram[2853]), .A2(n7419), .B1(n10566), .B2(n8980), .ZN(
        n7424) );
  INV_X1 U3801 ( .A(n7425), .ZN(n10556) );
  AOI22_X1 U3802 ( .A1(ram[2854]), .A2(n7419), .B1(n10566), .B2(n9004), .ZN(
        n7425) );
  INV_X1 U3803 ( .A(n7426), .ZN(n10557) );
  AOI22_X1 U3804 ( .A1(ram[2855]), .A2(n7419), .B1(n10566), .B2(n9028), .ZN(
        n7426) );
  INV_X1 U3805 ( .A(n7427), .ZN(n10558) );
  AOI22_X1 U3806 ( .A1(ram[2856]), .A2(n7419), .B1(n10566), .B2(n9052), .ZN(
        n7427) );
  INV_X1 U3807 ( .A(n7428), .ZN(n10559) );
  AOI22_X1 U3808 ( .A1(ram[2857]), .A2(n7419), .B1(n10566), .B2(n9076), .ZN(
        n7428) );
  INV_X1 U3809 ( .A(n7429), .ZN(n10560) );
  AOI22_X1 U3810 ( .A1(ram[2858]), .A2(n7419), .B1(n10566), .B2(n9100), .ZN(
        n7429) );
  INV_X1 U3811 ( .A(n7430), .ZN(n10561) );
  AOI22_X1 U3812 ( .A1(ram[2859]), .A2(n7419), .B1(n10566), .B2(n9124), .ZN(
        n7430) );
  INV_X1 U3813 ( .A(n7431), .ZN(n10562) );
  AOI22_X1 U3814 ( .A1(ram[2860]), .A2(n7419), .B1(n10566), .B2(n9148), .ZN(
        n7431) );
  INV_X1 U3815 ( .A(n7432), .ZN(n10563) );
  AOI22_X1 U3816 ( .A1(ram[2861]), .A2(n7419), .B1(n10566), .B2(n9172), .ZN(
        n7432) );
  INV_X1 U3817 ( .A(n7433), .ZN(n10564) );
  AOI22_X1 U3818 ( .A1(ram[2862]), .A2(n7419), .B1(n10566), .B2(n9196), .ZN(
        n7433) );
  INV_X1 U3819 ( .A(n7434), .ZN(n10565) );
  AOI22_X1 U3820 ( .A1(ram[2863]), .A2(n7419), .B1(n10566), .B2(n9220), .ZN(
        n7434) );
  INV_X1 U3821 ( .A(n7452), .ZN(n10516) );
  AOI22_X1 U3822 ( .A1(ram[2880]), .A2(n7453), .B1(n10532), .B2(n8860), .ZN(
        n7452) );
  INV_X1 U3823 ( .A(n7454), .ZN(n10517) );
  AOI22_X1 U3824 ( .A1(ram[2881]), .A2(n7453), .B1(n10532), .B2(n8884), .ZN(
        n7454) );
  INV_X1 U3825 ( .A(n7455), .ZN(n10518) );
  AOI22_X1 U3826 ( .A1(ram[2882]), .A2(n7453), .B1(n10532), .B2(n8908), .ZN(
        n7455) );
  INV_X1 U3827 ( .A(n7456), .ZN(n10519) );
  AOI22_X1 U3828 ( .A1(ram[2883]), .A2(n7453), .B1(n10532), .B2(n8932), .ZN(
        n7456) );
  INV_X1 U3829 ( .A(n7457), .ZN(n10520) );
  AOI22_X1 U3830 ( .A1(ram[2884]), .A2(n7453), .B1(n10532), .B2(n8956), .ZN(
        n7457) );
  INV_X1 U3831 ( .A(n7458), .ZN(n10521) );
  AOI22_X1 U3832 ( .A1(ram[2885]), .A2(n7453), .B1(n10532), .B2(n8980), .ZN(
        n7458) );
  INV_X1 U3833 ( .A(n7459), .ZN(n10522) );
  AOI22_X1 U3834 ( .A1(ram[2886]), .A2(n7453), .B1(n10532), .B2(n9004), .ZN(
        n7459) );
  INV_X1 U3835 ( .A(n7460), .ZN(n10523) );
  AOI22_X1 U3836 ( .A1(ram[2887]), .A2(n7453), .B1(n10532), .B2(n9028), .ZN(
        n7460) );
  INV_X1 U3837 ( .A(n7461), .ZN(n10524) );
  AOI22_X1 U3838 ( .A1(ram[2888]), .A2(n7453), .B1(n10532), .B2(n9052), .ZN(
        n7461) );
  INV_X1 U3839 ( .A(n7462), .ZN(n10525) );
  AOI22_X1 U3840 ( .A1(ram[2889]), .A2(n7453), .B1(n10532), .B2(n9076), .ZN(
        n7462) );
  INV_X1 U3841 ( .A(n7463), .ZN(n10526) );
  AOI22_X1 U3842 ( .A1(ram[2890]), .A2(n7453), .B1(n10532), .B2(n9100), .ZN(
        n7463) );
  INV_X1 U3843 ( .A(n7464), .ZN(n10527) );
  AOI22_X1 U3844 ( .A1(ram[2891]), .A2(n7453), .B1(n10532), .B2(n9124), .ZN(
        n7464) );
  INV_X1 U3845 ( .A(n7465), .ZN(n10528) );
  AOI22_X1 U3846 ( .A1(ram[2892]), .A2(n7453), .B1(n10532), .B2(n9148), .ZN(
        n7465) );
  INV_X1 U3847 ( .A(n7466), .ZN(n10529) );
  AOI22_X1 U3848 ( .A1(ram[2893]), .A2(n7453), .B1(n10532), .B2(n9172), .ZN(
        n7466) );
  INV_X1 U3849 ( .A(n7467), .ZN(n10530) );
  AOI22_X1 U3850 ( .A1(ram[2894]), .A2(n7453), .B1(n10532), .B2(n9196), .ZN(
        n7467) );
  INV_X1 U3851 ( .A(n7468), .ZN(n10531) );
  AOI22_X1 U3852 ( .A1(ram[2895]), .A2(n7453), .B1(n10532), .B2(n9220), .ZN(
        n7468) );
  INV_X1 U3853 ( .A(n7486), .ZN(n10482) );
  AOI22_X1 U3854 ( .A1(ram[2912]), .A2(n7487), .B1(n10498), .B2(n8860), .ZN(
        n7486) );
  INV_X1 U3855 ( .A(n7488), .ZN(n10483) );
  AOI22_X1 U3856 ( .A1(ram[2913]), .A2(n7487), .B1(n10498), .B2(n8884), .ZN(
        n7488) );
  INV_X1 U3857 ( .A(n7489), .ZN(n10484) );
  AOI22_X1 U3858 ( .A1(ram[2914]), .A2(n7487), .B1(n10498), .B2(n8908), .ZN(
        n7489) );
  INV_X1 U3859 ( .A(n7490), .ZN(n10485) );
  AOI22_X1 U3860 ( .A1(ram[2915]), .A2(n7487), .B1(n10498), .B2(n8932), .ZN(
        n7490) );
  INV_X1 U3861 ( .A(n7491), .ZN(n10486) );
  AOI22_X1 U3862 ( .A1(ram[2916]), .A2(n7487), .B1(n10498), .B2(n8956), .ZN(
        n7491) );
  INV_X1 U3863 ( .A(n7492), .ZN(n10487) );
  AOI22_X1 U3864 ( .A1(ram[2917]), .A2(n7487), .B1(n10498), .B2(n8980), .ZN(
        n7492) );
  INV_X1 U3865 ( .A(n7493), .ZN(n10488) );
  AOI22_X1 U3866 ( .A1(ram[2918]), .A2(n7487), .B1(n10498), .B2(n9004), .ZN(
        n7493) );
  INV_X1 U3867 ( .A(n7494), .ZN(n10489) );
  AOI22_X1 U3868 ( .A1(ram[2919]), .A2(n7487), .B1(n10498), .B2(n9028), .ZN(
        n7494) );
  INV_X1 U3869 ( .A(n7495), .ZN(n10490) );
  AOI22_X1 U3870 ( .A1(ram[2920]), .A2(n7487), .B1(n10498), .B2(n9052), .ZN(
        n7495) );
  INV_X1 U3871 ( .A(n7496), .ZN(n10491) );
  AOI22_X1 U3872 ( .A1(ram[2921]), .A2(n7487), .B1(n10498), .B2(n9076), .ZN(
        n7496) );
  INV_X1 U3873 ( .A(n7497), .ZN(n10492) );
  AOI22_X1 U3874 ( .A1(ram[2922]), .A2(n7487), .B1(n10498), .B2(n9100), .ZN(
        n7497) );
  INV_X1 U3875 ( .A(n7498), .ZN(n10493) );
  AOI22_X1 U3876 ( .A1(ram[2923]), .A2(n7487), .B1(n10498), .B2(n9124), .ZN(
        n7498) );
  INV_X1 U3877 ( .A(n7499), .ZN(n10494) );
  AOI22_X1 U3878 ( .A1(ram[2924]), .A2(n7487), .B1(n10498), .B2(n9148), .ZN(
        n7499) );
  INV_X1 U3879 ( .A(n7500), .ZN(n10495) );
  AOI22_X1 U3880 ( .A1(ram[2925]), .A2(n7487), .B1(n10498), .B2(n9172), .ZN(
        n7500) );
  INV_X1 U3881 ( .A(n7501), .ZN(n10496) );
  AOI22_X1 U3882 ( .A1(ram[2926]), .A2(n7487), .B1(n10498), .B2(n9196), .ZN(
        n7501) );
  INV_X1 U3883 ( .A(n7502), .ZN(n10497) );
  AOI22_X1 U3884 ( .A1(ram[2927]), .A2(n7487), .B1(n10498), .B2(n9220), .ZN(
        n7502) );
  INV_X1 U3885 ( .A(n7520), .ZN(n10448) );
  AOI22_X1 U3886 ( .A1(ram[2944]), .A2(n7521), .B1(n10464), .B2(n8859), .ZN(
        n7520) );
  INV_X1 U3887 ( .A(n7522), .ZN(n10449) );
  AOI22_X1 U3888 ( .A1(ram[2945]), .A2(n7521), .B1(n10464), .B2(n8883), .ZN(
        n7522) );
  INV_X1 U3889 ( .A(n7523), .ZN(n10450) );
  AOI22_X1 U3890 ( .A1(ram[2946]), .A2(n7521), .B1(n10464), .B2(n8907), .ZN(
        n7523) );
  INV_X1 U3891 ( .A(n7524), .ZN(n10451) );
  AOI22_X1 U3892 ( .A1(ram[2947]), .A2(n7521), .B1(n10464), .B2(n8931), .ZN(
        n7524) );
  INV_X1 U3893 ( .A(n7525), .ZN(n10452) );
  AOI22_X1 U3894 ( .A1(ram[2948]), .A2(n7521), .B1(n10464), .B2(n8955), .ZN(
        n7525) );
  INV_X1 U3895 ( .A(n7526), .ZN(n10453) );
  AOI22_X1 U3896 ( .A1(ram[2949]), .A2(n7521), .B1(n10464), .B2(n8979), .ZN(
        n7526) );
  INV_X1 U3897 ( .A(n7527), .ZN(n10454) );
  AOI22_X1 U3898 ( .A1(ram[2950]), .A2(n7521), .B1(n10464), .B2(n9003), .ZN(
        n7527) );
  INV_X1 U3899 ( .A(n7528), .ZN(n10455) );
  AOI22_X1 U3900 ( .A1(ram[2951]), .A2(n7521), .B1(n10464), .B2(n9027), .ZN(
        n7528) );
  INV_X1 U3901 ( .A(n7529), .ZN(n10456) );
  AOI22_X1 U3902 ( .A1(ram[2952]), .A2(n7521), .B1(n10464), .B2(n9051), .ZN(
        n7529) );
  INV_X1 U3903 ( .A(n7530), .ZN(n10457) );
  AOI22_X1 U3904 ( .A1(ram[2953]), .A2(n7521), .B1(n10464), .B2(n9075), .ZN(
        n7530) );
  INV_X1 U3905 ( .A(n7531), .ZN(n10458) );
  AOI22_X1 U3906 ( .A1(ram[2954]), .A2(n7521), .B1(n10464), .B2(n9099), .ZN(
        n7531) );
  INV_X1 U3907 ( .A(n7532), .ZN(n10459) );
  AOI22_X1 U3908 ( .A1(ram[2955]), .A2(n7521), .B1(n10464), .B2(n9123), .ZN(
        n7532) );
  INV_X1 U3909 ( .A(n7533), .ZN(n10460) );
  AOI22_X1 U3910 ( .A1(ram[2956]), .A2(n7521), .B1(n10464), .B2(n9147), .ZN(
        n7533) );
  INV_X1 U3911 ( .A(n7534), .ZN(n10461) );
  AOI22_X1 U3912 ( .A1(ram[2957]), .A2(n7521), .B1(n10464), .B2(n9171), .ZN(
        n7534) );
  INV_X1 U3913 ( .A(n7535), .ZN(n10462) );
  AOI22_X1 U3914 ( .A1(ram[2958]), .A2(n7521), .B1(n10464), .B2(n9195), .ZN(
        n7535) );
  INV_X1 U3915 ( .A(n7536), .ZN(n10463) );
  AOI22_X1 U3916 ( .A1(ram[2959]), .A2(n7521), .B1(n10464), .B2(n9219), .ZN(
        n7536) );
  INV_X1 U3917 ( .A(n7554), .ZN(n10414) );
  AOI22_X1 U3918 ( .A1(ram[2976]), .A2(n7555), .B1(n10430), .B2(n8859), .ZN(
        n7554) );
  INV_X1 U3919 ( .A(n7556), .ZN(n10415) );
  AOI22_X1 U3920 ( .A1(ram[2977]), .A2(n7555), .B1(n10430), .B2(n8883), .ZN(
        n7556) );
  INV_X1 U3921 ( .A(n7557), .ZN(n10416) );
  AOI22_X1 U3922 ( .A1(ram[2978]), .A2(n7555), .B1(n10430), .B2(n8907), .ZN(
        n7557) );
  INV_X1 U3923 ( .A(n7558), .ZN(n10417) );
  AOI22_X1 U3924 ( .A1(ram[2979]), .A2(n7555), .B1(n10430), .B2(n8931), .ZN(
        n7558) );
  INV_X1 U3925 ( .A(n7559), .ZN(n10418) );
  AOI22_X1 U3926 ( .A1(ram[2980]), .A2(n7555), .B1(n10430), .B2(n8955), .ZN(
        n7559) );
  INV_X1 U3927 ( .A(n7560), .ZN(n10419) );
  AOI22_X1 U3928 ( .A1(ram[2981]), .A2(n7555), .B1(n10430), .B2(n8979), .ZN(
        n7560) );
  INV_X1 U3929 ( .A(n7561), .ZN(n10420) );
  AOI22_X1 U3930 ( .A1(ram[2982]), .A2(n7555), .B1(n10430), .B2(n9003), .ZN(
        n7561) );
  INV_X1 U3931 ( .A(n7562), .ZN(n10421) );
  AOI22_X1 U3932 ( .A1(ram[2983]), .A2(n7555), .B1(n10430), .B2(n9027), .ZN(
        n7562) );
  INV_X1 U3933 ( .A(n7563), .ZN(n10422) );
  AOI22_X1 U3934 ( .A1(ram[2984]), .A2(n7555), .B1(n10430), .B2(n9051), .ZN(
        n7563) );
  INV_X1 U3935 ( .A(n7564), .ZN(n10423) );
  AOI22_X1 U3936 ( .A1(ram[2985]), .A2(n7555), .B1(n10430), .B2(n9075), .ZN(
        n7564) );
  INV_X1 U3937 ( .A(n7565), .ZN(n10424) );
  AOI22_X1 U3938 ( .A1(ram[2986]), .A2(n7555), .B1(n10430), .B2(n9099), .ZN(
        n7565) );
  INV_X1 U3939 ( .A(n7566), .ZN(n10425) );
  AOI22_X1 U3940 ( .A1(ram[2987]), .A2(n7555), .B1(n10430), .B2(n9123), .ZN(
        n7566) );
  INV_X1 U3941 ( .A(n7567), .ZN(n10426) );
  AOI22_X1 U3942 ( .A1(ram[2988]), .A2(n7555), .B1(n10430), .B2(n9147), .ZN(
        n7567) );
  INV_X1 U3943 ( .A(n7568), .ZN(n10427) );
  AOI22_X1 U3944 ( .A1(ram[2989]), .A2(n7555), .B1(n10430), .B2(n9171), .ZN(
        n7568) );
  INV_X1 U3945 ( .A(n7569), .ZN(n10428) );
  AOI22_X1 U3946 ( .A1(ram[2990]), .A2(n7555), .B1(n10430), .B2(n9195), .ZN(
        n7569) );
  INV_X1 U3947 ( .A(n7570), .ZN(n10429) );
  AOI22_X1 U3948 ( .A1(ram[2991]), .A2(n7555), .B1(n10430), .B2(n9219), .ZN(
        n7570) );
  INV_X1 U3949 ( .A(n7588), .ZN(n10380) );
  AOI22_X1 U3950 ( .A1(ram[3008]), .A2(n7589), .B1(n10396), .B2(n8859), .ZN(
        n7588) );
  INV_X1 U3951 ( .A(n7590), .ZN(n10381) );
  AOI22_X1 U3952 ( .A1(ram[3009]), .A2(n7589), .B1(n10396), .B2(n8883), .ZN(
        n7590) );
  INV_X1 U3953 ( .A(n7591), .ZN(n10382) );
  AOI22_X1 U3954 ( .A1(ram[3010]), .A2(n7589), .B1(n10396), .B2(n8907), .ZN(
        n7591) );
  INV_X1 U3955 ( .A(n7592), .ZN(n10383) );
  AOI22_X1 U3956 ( .A1(ram[3011]), .A2(n7589), .B1(n10396), .B2(n8931), .ZN(
        n7592) );
  INV_X1 U3957 ( .A(n7593), .ZN(n10384) );
  AOI22_X1 U3958 ( .A1(ram[3012]), .A2(n7589), .B1(n10396), .B2(n8955), .ZN(
        n7593) );
  INV_X1 U3959 ( .A(n7594), .ZN(n10385) );
  AOI22_X1 U3960 ( .A1(ram[3013]), .A2(n7589), .B1(n10396), .B2(n8979), .ZN(
        n7594) );
  INV_X1 U3961 ( .A(n7595), .ZN(n10386) );
  AOI22_X1 U3962 ( .A1(ram[3014]), .A2(n7589), .B1(n10396), .B2(n9003), .ZN(
        n7595) );
  INV_X1 U3963 ( .A(n7596), .ZN(n10387) );
  AOI22_X1 U3964 ( .A1(ram[3015]), .A2(n7589), .B1(n10396), .B2(n9027), .ZN(
        n7596) );
  INV_X1 U3965 ( .A(n7597), .ZN(n10388) );
  AOI22_X1 U3966 ( .A1(ram[3016]), .A2(n7589), .B1(n10396), .B2(n9051), .ZN(
        n7597) );
  INV_X1 U3967 ( .A(n7598), .ZN(n10389) );
  AOI22_X1 U3968 ( .A1(ram[3017]), .A2(n7589), .B1(n10396), .B2(n9075), .ZN(
        n7598) );
  INV_X1 U3969 ( .A(n7599), .ZN(n10390) );
  AOI22_X1 U3970 ( .A1(ram[3018]), .A2(n7589), .B1(n10396), .B2(n9099), .ZN(
        n7599) );
  INV_X1 U3971 ( .A(n7600), .ZN(n10391) );
  AOI22_X1 U3972 ( .A1(ram[3019]), .A2(n7589), .B1(n10396), .B2(n9123), .ZN(
        n7600) );
  INV_X1 U3973 ( .A(n7601), .ZN(n10392) );
  AOI22_X1 U3974 ( .A1(ram[3020]), .A2(n7589), .B1(n10396), .B2(n9147), .ZN(
        n7601) );
  INV_X1 U3975 ( .A(n7602), .ZN(n10393) );
  AOI22_X1 U3976 ( .A1(ram[3021]), .A2(n7589), .B1(n10396), .B2(n9171), .ZN(
        n7602) );
  INV_X1 U3977 ( .A(n7603), .ZN(n10394) );
  AOI22_X1 U3978 ( .A1(ram[3022]), .A2(n7589), .B1(n10396), .B2(n9195), .ZN(
        n7603) );
  INV_X1 U3979 ( .A(n7604), .ZN(n10395) );
  AOI22_X1 U3980 ( .A1(ram[3023]), .A2(n7589), .B1(n10396), .B2(n9219), .ZN(
        n7604) );
  INV_X1 U3981 ( .A(n7622), .ZN(n10346) );
  AOI22_X1 U3982 ( .A1(ram[3040]), .A2(n7623), .B1(n10362), .B2(n8859), .ZN(
        n7622) );
  INV_X1 U3983 ( .A(n7624), .ZN(n10347) );
  AOI22_X1 U3984 ( .A1(ram[3041]), .A2(n7623), .B1(n10362), .B2(n8883), .ZN(
        n7624) );
  INV_X1 U3985 ( .A(n7625), .ZN(n10348) );
  AOI22_X1 U3986 ( .A1(ram[3042]), .A2(n7623), .B1(n10362), .B2(n8907), .ZN(
        n7625) );
  INV_X1 U3987 ( .A(n7626), .ZN(n10349) );
  AOI22_X1 U3988 ( .A1(ram[3043]), .A2(n7623), .B1(n10362), .B2(n8931), .ZN(
        n7626) );
  INV_X1 U3989 ( .A(n7627), .ZN(n10350) );
  AOI22_X1 U3990 ( .A1(ram[3044]), .A2(n7623), .B1(n10362), .B2(n8955), .ZN(
        n7627) );
  INV_X1 U3991 ( .A(n7628), .ZN(n10351) );
  AOI22_X1 U3992 ( .A1(ram[3045]), .A2(n7623), .B1(n10362), .B2(n8979), .ZN(
        n7628) );
  INV_X1 U3993 ( .A(n7629), .ZN(n10352) );
  AOI22_X1 U3994 ( .A1(ram[3046]), .A2(n7623), .B1(n10362), .B2(n9003), .ZN(
        n7629) );
  INV_X1 U3995 ( .A(n7630), .ZN(n10353) );
  AOI22_X1 U3996 ( .A1(ram[3047]), .A2(n7623), .B1(n10362), .B2(n9027), .ZN(
        n7630) );
  INV_X1 U3997 ( .A(n7631), .ZN(n10354) );
  AOI22_X1 U3998 ( .A1(ram[3048]), .A2(n7623), .B1(n10362), .B2(n9051), .ZN(
        n7631) );
  INV_X1 U3999 ( .A(n7632), .ZN(n10355) );
  AOI22_X1 U4000 ( .A1(ram[3049]), .A2(n7623), .B1(n10362), .B2(n9075), .ZN(
        n7632) );
  INV_X1 U4001 ( .A(n7633), .ZN(n10356) );
  AOI22_X1 U4002 ( .A1(ram[3050]), .A2(n7623), .B1(n10362), .B2(n9099), .ZN(
        n7633) );
  INV_X1 U4003 ( .A(n7634), .ZN(n10357) );
  AOI22_X1 U4004 ( .A1(ram[3051]), .A2(n7623), .B1(n10362), .B2(n9123), .ZN(
        n7634) );
  INV_X1 U4005 ( .A(n7635), .ZN(n10358) );
  AOI22_X1 U4006 ( .A1(ram[3052]), .A2(n7623), .B1(n10362), .B2(n9147), .ZN(
        n7635) );
  INV_X1 U4007 ( .A(n7636), .ZN(n10359) );
  AOI22_X1 U4008 ( .A1(ram[3053]), .A2(n7623), .B1(n10362), .B2(n9171), .ZN(
        n7636) );
  INV_X1 U4009 ( .A(n7637), .ZN(n10360) );
  AOI22_X1 U4010 ( .A1(ram[3054]), .A2(n7623), .B1(n10362), .B2(n9195), .ZN(
        n7637) );
  INV_X1 U4011 ( .A(n7638), .ZN(n10361) );
  AOI22_X1 U4012 ( .A1(ram[3055]), .A2(n7623), .B1(n10362), .B2(n9219), .ZN(
        n7638) );
  INV_X1 U4013 ( .A(n7656), .ZN(n10312) );
  AOI22_X1 U4014 ( .A1(ram[3072]), .A2(n7657), .B1(n10328), .B2(n8859), .ZN(
        n7656) );
  INV_X1 U4015 ( .A(n7658), .ZN(n10313) );
  AOI22_X1 U4016 ( .A1(ram[3073]), .A2(n7657), .B1(n10328), .B2(n8883), .ZN(
        n7658) );
  INV_X1 U4017 ( .A(n7659), .ZN(n10314) );
  AOI22_X1 U4018 ( .A1(ram[3074]), .A2(n7657), .B1(n10328), .B2(n8907), .ZN(
        n7659) );
  INV_X1 U4019 ( .A(n7660), .ZN(n10315) );
  AOI22_X1 U4020 ( .A1(ram[3075]), .A2(n7657), .B1(n10328), .B2(n8931), .ZN(
        n7660) );
  INV_X1 U4021 ( .A(n7661), .ZN(n10316) );
  AOI22_X1 U4022 ( .A1(ram[3076]), .A2(n7657), .B1(n10328), .B2(n8955), .ZN(
        n7661) );
  INV_X1 U4023 ( .A(n7662), .ZN(n10317) );
  AOI22_X1 U4024 ( .A1(ram[3077]), .A2(n7657), .B1(n10328), .B2(n8979), .ZN(
        n7662) );
  INV_X1 U4025 ( .A(n7663), .ZN(n10318) );
  AOI22_X1 U4026 ( .A1(ram[3078]), .A2(n7657), .B1(n10328), .B2(n9003), .ZN(
        n7663) );
  INV_X1 U4027 ( .A(n7664), .ZN(n10319) );
  AOI22_X1 U4028 ( .A1(ram[3079]), .A2(n7657), .B1(n10328), .B2(n9027), .ZN(
        n7664) );
  INV_X1 U4029 ( .A(n7665), .ZN(n10320) );
  AOI22_X1 U4030 ( .A1(ram[3080]), .A2(n7657), .B1(n10328), .B2(n9051), .ZN(
        n7665) );
  INV_X1 U4031 ( .A(n7666), .ZN(n10321) );
  AOI22_X1 U4032 ( .A1(ram[3081]), .A2(n7657), .B1(n10328), .B2(n9075), .ZN(
        n7666) );
  INV_X1 U4033 ( .A(n7667), .ZN(n10322) );
  AOI22_X1 U4034 ( .A1(ram[3082]), .A2(n7657), .B1(n10328), .B2(n9099), .ZN(
        n7667) );
  INV_X1 U4035 ( .A(n7668), .ZN(n10323) );
  AOI22_X1 U4036 ( .A1(ram[3083]), .A2(n7657), .B1(n10328), .B2(n9123), .ZN(
        n7668) );
  INV_X1 U4037 ( .A(n7669), .ZN(n10324) );
  AOI22_X1 U4038 ( .A1(ram[3084]), .A2(n7657), .B1(n10328), .B2(n9147), .ZN(
        n7669) );
  INV_X1 U4039 ( .A(n7670), .ZN(n10325) );
  AOI22_X1 U4040 ( .A1(ram[3085]), .A2(n7657), .B1(n10328), .B2(n9171), .ZN(
        n7670) );
  INV_X1 U4041 ( .A(n7671), .ZN(n10326) );
  AOI22_X1 U4042 ( .A1(ram[3086]), .A2(n7657), .B1(n10328), .B2(n9195), .ZN(
        n7671) );
  INV_X1 U4043 ( .A(n7672), .ZN(n10327) );
  AOI22_X1 U4044 ( .A1(ram[3087]), .A2(n7657), .B1(n10328), .B2(n9219), .ZN(
        n7672) );
  INV_X1 U4045 ( .A(n7691), .ZN(n10278) );
  AOI22_X1 U4046 ( .A1(ram[3104]), .A2(n7692), .B1(n10294), .B2(n8859), .ZN(
        n7691) );
  INV_X1 U4047 ( .A(n7693), .ZN(n10279) );
  AOI22_X1 U4048 ( .A1(ram[3105]), .A2(n7692), .B1(n10294), .B2(n8883), .ZN(
        n7693) );
  INV_X1 U4049 ( .A(n7694), .ZN(n10280) );
  AOI22_X1 U4050 ( .A1(ram[3106]), .A2(n7692), .B1(n10294), .B2(n8907), .ZN(
        n7694) );
  INV_X1 U4051 ( .A(n7695), .ZN(n10281) );
  AOI22_X1 U4052 ( .A1(ram[3107]), .A2(n7692), .B1(n10294), .B2(n8931), .ZN(
        n7695) );
  INV_X1 U4053 ( .A(n7696), .ZN(n10282) );
  AOI22_X1 U4054 ( .A1(ram[3108]), .A2(n7692), .B1(n10294), .B2(n8955), .ZN(
        n7696) );
  INV_X1 U4055 ( .A(n7697), .ZN(n10283) );
  AOI22_X1 U4056 ( .A1(ram[3109]), .A2(n7692), .B1(n10294), .B2(n8979), .ZN(
        n7697) );
  INV_X1 U4057 ( .A(n7698), .ZN(n10284) );
  AOI22_X1 U4058 ( .A1(ram[3110]), .A2(n7692), .B1(n10294), .B2(n9003), .ZN(
        n7698) );
  INV_X1 U4059 ( .A(n7699), .ZN(n10285) );
  AOI22_X1 U4060 ( .A1(ram[3111]), .A2(n7692), .B1(n10294), .B2(n9027), .ZN(
        n7699) );
  INV_X1 U4061 ( .A(n7700), .ZN(n10286) );
  AOI22_X1 U4062 ( .A1(ram[3112]), .A2(n7692), .B1(n10294), .B2(n9051), .ZN(
        n7700) );
  INV_X1 U4063 ( .A(n7701), .ZN(n10287) );
  AOI22_X1 U4064 ( .A1(ram[3113]), .A2(n7692), .B1(n10294), .B2(n9075), .ZN(
        n7701) );
  INV_X1 U4065 ( .A(n7702), .ZN(n10288) );
  AOI22_X1 U4066 ( .A1(ram[3114]), .A2(n7692), .B1(n10294), .B2(n9099), .ZN(
        n7702) );
  INV_X1 U4067 ( .A(n7703), .ZN(n10289) );
  AOI22_X1 U4068 ( .A1(ram[3115]), .A2(n7692), .B1(n10294), .B2(n9123), .ZN(
        n7703) );
  INV_X1 U4069 ( .A(n7704), .ZN(n10290) );
  AOI22_X1 U4070 ( .A1(ram[3116]), .A2(n7692), .B1(n10294), .B2(n9147), .ZN(
        n7704) );
  INV_X1 U4071 ( .A(n7705), .ZN(n10291) );
  AOI22_X1 U4072 ( .A1(ram[3117]), .A2(n7692), .B1(n10294), .B2(n9171), .ZN(
        n7705) );
  INV_X1 U4073 ( .A(n7706), .ZN(n10292) );
  AOI22_X1 U4074 ( .A1(ram[3118]), .A2(n7692), .B1(n10294), .B2(n9195), .ZN(
        n7706) );
  INV_X1 U4075 ( .A(n7707), .ZN(n10293) );
  AOI22_X1 U4076 ( .A1(ram[3119]), .A2(n7692), .B1(n10294), .B2(n9219), .ZN(
        n7707) );
  INV_X1 U4077 ( .A(n7725), .ZN(n10244) );
  AOI22_X1 U4078 ( .A1(ram[3136]), .A2(n7726), .B1(n10260), .B2(n8858), .ZN(
        n7725) );
  INV_X1 U4079 ( .A(n7727), .ZN(n10245) );
  AOI22_X1 U4080 ( .A1(ram[3137]), .A2(n7726), .B1(n10260), .B2(n8882), .ZN(
        n7727) );
  INV_X1 U4081 ( .A(n7728), .ZN(n10246) );
  AOI22_X1 U4082 ( .A1(ram[3138]), .A2(n7726), .B1(n10260), .B2(n8906), .ZN(
        n7728) );
  INV_X1 U4083 ( .A(n7729), .ZN(n10247) );
  AOI22_X1 U4084 ( .A1(ram[3139]), .A2(n7726), .B1(n10260), .B2(n8930), .ZN(
        n7729) );
  INV_X1 U4085 ( .A(n7730), .ZN(n10248) );
  AOI22_X1 U4086 ( .A1(ram[3140]), .A2(n7726), .B1(n10260), .B2(n8954), .ZN(
        n7730) );
  INV_X1 U4087 ( .A(n7731), .ZN(n10249) );
  AOI22_X1 U4088 ( .A1(ram[3141]), .A2(n7726), .B1(n10260), .B2(n8978), .ZN(
        n7731) );
  INV_X1 U4089 ( .A(n7732), .ZN(n10250) );
  AOI22_X1 U4090 ( .A1(ram[3142]), .A2(n7726), .B1(n10260), .B2(n9002), .ZN(
        n7732) );
  INV_X1 U4091 ( .A(n7733), .ZN(n10251) );
  AOI22_X1 U4092 ( .A1(ram[3143]), .A2(n7726), .B1(n10260), .B2(n9026), .ZN(
        n7733) );
  INV_X1 U4093 ( .A(n7734), .ZN(n10252) );
  AOI22_X1 U4094 ( .A1(ram[3144]), .A2(n7726), .B1(n10260), .B2(n9050), .ZN(
        n7734) );
  INV_X1 U4095 ( .A(n7735), .ZN(n10253) );
  AOI22_X1 U4096 ( .A1(ram[3145]), .A2(n7726), .B1(n10260), .B2(n9074), .ZN(
        n7735) );
  INV_X1 U4097 ( .A(n7736), .ZN(n10254) );
  AOI22_X1 U4098 ( .A1(ram[3146]), .A2(n7726), .B1(n10260), .B2(n9098), .ZN(
        n7736) );
  INV_X1 U4099 ( .A(n7737), .ZN(n10255) );
  AOI22_X1 U4100 ( .A1(ram[3147]), .A2(n7726), .B1(n10260), .B2(n9122), .ZN(
        n7737) );
  INV_X1 U4101 ( .A(n7738), .ZN(n10256) );
  AOI22_X1 U4102 ( .A1(ram[3148]), .A2(n7726), .B1(n10260), .B2(n9146), .ZN(
        n7738) );
  INV_X1 U4103 ( .A(n7739), .ZN(n10257) );
  AOI22_X1 U4104 ( .A1(ram[3149]), .A2(n7726), .B1(n10260), .B2(n9170), .ZN(
        n7739) );
  INV_X1 U4105 ( .A(n7740), .ZN(n10258) );
  AOI22_X1 U4106 ( .A1(ram[3150]), .A2(n7726), .B1(n10260), .B2(n9194), .ZN(
        n7740) );
  INV_X1 U4107 ( .A(n7741), .ZN(n10259) );
  AOI22_X1 U4108 ( .A1(ram[3151]), .A2(n7726), .B1(n10260), .B2(n9218), .ZN(
        n7741) );
  INV_X1 U4109 ( .A(n7759), .ZN(n10210) );
  AOI22_X1 U4110 ( .A1(ram[3168]), .A2(n7760), .B1(n10226), .B2(n8858), .ZN(
        n7759) );
  INV_X1 U4111 ( .A(n7761), .ZN(n10211) );
  AOI22_X1 U4112 ( .A1(ram[3169]), .A2(n7760), .B1(n10226), .B2(n8882), .ZN(
        n7761) );
  INV_X1 U4113 ( .A(n7762), .ZN(n10212) );
  AOI22_X1 U4114 ( .A1(ram[3170]), .A2(n7760), .B1(n10226), .B2(n8906), .ZN(
        n7762) );
  INV_X1 U4115 ( .A(n7763), .ZN(n10213) );
  AOI22_X1 U4116 ( .A1(ram[3171]), .A2(n7760), .B1(n10226), .B2(n8930), .ZN(
        n7763) );
  INV_X1 U4117 ( .A(n7764), .ZN(n10214) );
  AOI22_X1 U4118 ( .A1(ram[3172]), .A2(n7760), .B1(n10226), .B2(n8954), .ZN(
        n7764) );
  INV_X1 U4119 ( .A(n7765), .ZN(n10215) );
  AOI22_X1 U4120 ( .A1(ram[3173]), .A2(n7760), .B1(n10226), .B2(n8978), .ZN(
        n7765) );
  INV_X1 U4121 ( .A(n7766), .ZN(n10216) );
  AOI22_X1 U4122 ( .A1(ram[3174]), .A2(n7760), .B1(n10226), .B2(n9002), .ZN(
        n7766) );
  INV_X1 U4123 ( .A(n7767), .ZN(n10217) );
  AOI22_X1 U4124 ( .A1(ram[3175]), .A2(n7760), .B1(n10226), .B2(n9026), .ZN(
        n7767) );
  INV_X1 U4125 ( .A(n7768), .ZN(n10218) );
  AOI22_X1 U4126 ( .A1(ram[3176]), .A2(n7760), .B1(n10226), .B2(n9050), .ZN(
        n7768) );
  INV_X1 U4127 ( .A(n7769), .ZN(n10219) );
  AOI22_X1 U4128 ( .A1(ram[3177]), .A2(n7760), .B1(n10226), .B2(n9074), .ZN(
        n7769) );
  INV_X1 U4129 ( .A(n7770), .ZN(n10220) );
  AOI22_X1 U4130 ( .A1(ram[3178]), .A2(n7760), .B1(n10226), .B2(n9098), .ZN(
        n7770) );
  INV_X1 U4131 ( .A(n7771), .ZN(n10221) );
  AOI22_X1 U4132 ( .A1(ram[3179]), .A2(n7760), .B1(n10226), .B2(n9122), .ZN(
        n7771) );
  INV_X1 U4133 ( .A(n7772), .ZN(n10222) );
  AOI22_X1 U4134 ( .A1(ram[3180]), .A2(n7760), .B1(n10226), .B2(n9146), .ZN(
        n7772) );
  INV_X1 U4135 ( .A(n7773), .ZN(n10223) );
  AOI22_X1 U4136 ( .A1(ram[3181]), .A2(n7760), .B1(n10226), .B2(n9170), .ZN(
        n7773) );
  INV_X1 U4137 ( .A(n7774), .ZN(n10224) );
  AOI22_X1 U4138 ( .A1(ram[3182]), .A2(n7760), .B1(n10226), .B2(n9194), .ZN(
        n7774) );
  INV_X1 U4139 ( .A(n7775), .ZN(n10225) );
  AOI22_X1 U4140 ( .A1(ram[3183]), .A2(n7760), .B1(n10226), .B2(n9218), .ZN(
        n7775) );
  INV_X1 U4141 ( .A(n7793), .ZN(n10176) );
  AOI22_X1 U4142 ( .A1(ram[3200]), .A2(n7794), .B1(n10192), .B2(n8858), .ZN(
        n7793) );
  INV_X1 U4143 ( .A(n7795), .ZN(n10177) );
  AOI22_X1 U4144 ( .A1(ram[3201]), .A2(n7794), .B1(n10192), .B2(n8882), .ZN(
        n7795) );
  INV_X1 U4145 ( .A(n7796), .ZN(n10178) );
  AOI22_X1 U4146 ( .A1(ram[3202]), .A2(n7794), .B1(n10192), .B2(n8906), .ZN(
        n7796) );
  INV_X1 U4147 ( .A(n7797), .ZN(n10179) );
  AOI22_X1 U4148 ( .A1(ram[3203]), .A2(n7794), .B1(n10192), .B2(n8930), .ZN(
        n7797) );
  INV_X1 U4149 ( .A(n7798), .ZN(n10180) );
  AOI22_X1 U4150 ( .A1(ram[3204]), .A2(n7794), .B1(n10192), .B2(n8954), .ZN(
        n7798) );
  INV_X1 U4151 ( .A(n7799), .ZN(n10181) );
  AOI22_X1 U4152 ( .A1(ram[3205]), .A2(n7794), .B1(n10192), .B2(n8978), .ZN(
        n7799) );
  INV_X1 U4153 ( .A(n7800), .ZN(n10182) );
  AOI22_X1 U4154 ( .A1(ram[3206]), .A2(n7794), .B1(n10192), .B2(n9002), .ZN(
        n7800) );
  INV_X1 U4155 ( .A(n7801), .ZN(n10183) );
  AOI22_X1 U4156 ( .A1(ram[3207]), .A2(n7794), .B1(n10192), .B2(n9026), .ZN(
        n7801) );
  INV_X1 U4157 ( .A(n7802), .ZN(n10184) );
  AOI22_X1 U4158 ( .A1(ram[3208]), .A2(n7794), .B1(n10192), .B2(n9050), .ZN(
        n7802) );
  INV_X1 U4159 ( .A(n7803), .ZN(n10185) );
  AOI22_X1 U4160 ( .A1(ram[3209]), .A2(n7794), .B1(n10192), .B2(n9074), .ZN(
        n7803) );
  INV_X1 U4161 ( .A(n7804), .ZN(n10186) );
  AOI22_X1 U4162 ( .A1(ram[3210]), .A2(n7794), .B1(n10192), .B2(n9098), .ZN(
        n7804) );
  INV_X1 U4163 ( .A(n7805), .ZN(n10187) );
  AOI22_X1 U4164 ( .A1(ram[3211]), .A2(n7794), .B1(n10192), .B2(n9122), .ZN(
        n7805) );
  INV_X1 U4165 ( .A(n7806), .ZN(n10188) );
  AOI22_X1 U4166 ( .A1(ram[3212]), .A2(n7794), .B1(n10192), .B2(n9146), .ZN(
        n7806) );
  INV_X1 U4167 ( .A(n7807), .ZN(n10189) );
  AOI22_X1 U4168 ( .A1(ram[3213]), .A2(n7794), .B1(n10192), .B2(n9170), .ZN(
        n7807) );
  INV_X1 U4169 ( .A(n7808), .ZN(n10190) );
  AOI22_X1 U4170 ( .A1(ram[3214]), .A2(n7794), .B1(n10192), .B2(n9194), .ZN(
        n7808) );
  INV_X1 U4171 ( .A(n7809), .ZN(n10191) );
  AOI22_X1 U4172 ( .A1(ram[3215]), .A2(n7794), .B1(n10192), .B2(n9218), .ZN(
        n7809) );
  INV_X1 U4173 ( .A(n7827), .ZN(n10142) );
  AOI22_X1 U4174 ( .A1(ram[3232]), .A2(n7828), .B1(n10158), .B2(n8858), .ZN(
        n7827) );
  INV_X1 U4175 ( .A(n7829), .ZN(n10143) );
  AOI22_X1 U4176 ( .A1(ram[3233]), .A2(n7828), .B1(n10158), .B2(n8882), .ZN(
        n7829) );
  INV_X1 U4177 ( .A(n7830), .ZN(n10144) );
  AOI22_X1 U4178 ( .A1(ram[3234]), .A2(n7828), .B1(n10158), .B2(n8906), .ZN(
        n7830) );
  INV_X1 U4179 ( .A(n7831), .ZN(n10145) );
  AOI22_X1 U4180 ( .A1(ram[3235]), .A2(n7828), .B1(n10158), .B2(n8930), .ZN(
        n7831) );
  INV_X1 U4181 ( .A(n7832), .ZN(n10146) );
  AOI22_X1 U4182 ( .A1(ram[3236]), .A2(n7828), .B1(n10158), .B2(n8954), .ZN(
        n7832) );
  INV_X1 U4183 ( .A(n7833), .ZN(n10147) );
  AOI22_X1 U4184 ( .A1(ram[3237]), .A2(n7828), .B1(n10158), .B2(n8978), .ZN(
        n7833) );
  INV_X1 U4185 ( .A(n7834), .ZN(n10148) );
  AOI22_X1 U4186 ( .A1(ram[3238]), .A2(n7828), .B1(n10158), .B2(n9002), .ZN(
        n7834) );
  INV_X1 U4187 ( .A(n7835), .ZN(n10149) );
  AOI22_X1 U4188 ( .A1(ram[3239]), .A2(n7828), .B1(n10158), .B2(n9026), .ZN(
        n7835) );
  INV_X1 U4189 ( .A(n7836), .ZN(n10150) );
  AOI22_X1 U4190 ( .A1(ram[3240]), .A2(n7828), .B1(n10158), .B2(n9050), .ZN(
        n7836) );
  INV_X1 U4191 ( .A(n7837), .ZN(n10151) );
  AOI22_X1 U4192 ( .A1(ram[3241]), .A2(n7828), .B1(n10158), .B2(n9074), .ZN(
        n7837) );
  INV_X1 U4193 ( .A(n7838), .ZN(n10152) );
  AOI22_X1 U4194 ( .A1(ram[3242]), .A2(n7828), .B1(n10158), .B2(n9098), .ZN(
        n7838) );
  INV_X1 U4195 ( .A(n7839), .ZN(n10153) );
  AOI22_X1 U4196 ( .A1(ram[3243]), .A2(n7828), .B1(n10158), .B2(n9122), .ZN(
        n7839) );
  INV_X1 U4197 ( .A(n7840), .ZN(n10154) );
  AOI22_X1 U4198 ( .A1(ram[3244]), .A2(n7828), .B1(n10158), .B2(n9146), .ZN(
        n7840) );
  INV_X1 U4199 ( .A(n7841), .ZN(n10155) );
  AOI22_X1 U4200 ( .A1(ram[3245]), .A2(n7828), .B1(n10158), .B2(n9170), .ZN(
        n7841) );
  INV_X1 U4201 ( .A(n7842), .ZN(n10156) );
  AOI22_X1 U4202 ( .A1(ram[3246]), .A2(n7828), .B1(n10158), .B2(n9194), .ZN(
        n7842) );
  INV_X1 U4203 ( .A(n7843), .ZN(n10157) );
  AOI22_X1 U4204 ( .A1(ram[3247]), .A2(n7828), .B1(n10158), .B2(n9218), .ZN(
        n7843) );
  INV_X1 U4205 ( .A(n7861), .ZN(n10108) );
  AOI22_X1 U4206 ( .A1(ram[3264]), .A2(n7862), .B1(n10124), .B2(n8858), .ZN(
        n7861) );
  INV_X1 U4207 ( .A(n7863), .ZN(n10109) );
  AOI22_X1 U4208 ( .A1(ram[3265]), .A2(n7862), .B1(n10124), .B2(n8882), .ZN(
        n7863) );
  INV_X1 U4209 ( .A(n7864), .ZN(n10110) );
  AOI22_X1 U4210 ( .A1(ram[3266]), .A2(n7862), .B1(n10124), .B2(n8906), .ZN(
        n7864) );
  INV_X1 U4211 ( .A(n7865), .ZN(n10111) );
  AOI22_X1 U4212 ( .A1(ram[3267]), .A2(n7862), .B1(n10124), .B2(n8930), .ZN(
        n7865) );
  INV_X1 U4213 ( .A(n7866), .ZN(n10112) );
  AOI22_X1 U4214 ( .A1(ram[3268]), .A2(n7862), .B1(n10124), .B2(n8954), .ZN(
        n7866) );
  INV_X1 U4215 ( .A(n7867), .ZN(n10113) );
  AOI22_X1 U4216 ( .A1(ram[3269]), .A2(n7862), .B1(n10124), .B2(n8978), .ZN(
        n7867) );
  INV_X1 U4217 ( .A(n7868), .ZN(n10114) );
  AOI22_X1 U4218 ( .A1(ram[3270]), .A2(n7862), .B1(n10124), .B2(n9002), .ZN(
        n7868) );
  INV_X1 U4219 ( .A(n7869), .ZN(n10115) );
  AOI22_X1 U4220 ( .A1(ram[3271]), .A2(n7862), .B1(n10124), .B2(n9026), .ZN(
        n7869) );
  INV_X1 U4221 ( .A(n7870), .ZN(n10116) );
  AOI22_X1 U4222 ( .A1(ram[3272]), .A2(n7862), .B1(n10124), .B2(n9050), .ZN(
        n7870) );
  INV_X1 U4223 ( .A(n7871), .ZN(n10117) );
  AOI22_X1 U4224 ( .A1(ram[3273]), .A2(n7862), .B1(n10124), .B2(n9074), .ZN(
        n7871) );
  INV_X1 U4225 ( .A(n7872), .ZN(n10118) );
  AOI22_X1 U4226 ( .A1(ram[3274]), .A2(n7862), .B1(n10124), .B2(n9098), .ZN(
        n7872) );
  INV_X1 U4227 ( .A(n7873), .ZN(n10119) );
  AOI22_X1 U4228 ( .A1(ram[3275]), .A2(n7862), .B1(n10124), .B2(n9122), .ZN(
        n7873) );
  INV_X1 U4229 ( .A(n7874), .ZN(n10120) );
  AOI22_X1 U4230 ( .A1(ram[3276]), .A2(n7862), .B1(n10124), .B2(n9146), .ZN(
        n7874) );
  INV_X1 U4231 ( .A(n7875), .ZN(n10121) );
  AOI22_X1 U4232 ( .A1(ram[3277]), .A2(n7862), .B1(n10124), .B2(n9170), .ZN(
        n7875) );
  INV_X1 U4233 ( .A(n7876), .ZN(n10122) );
  AOI22_X1 U4234 ( .A1(ram[3278]), .A2(n7862), .B1(n10124), .B2(n9194), .ZN(
        n7876) );
  INV_X1 U4235 ( .A(n7877), .ZN(n10123) );
  AOI22_X1 U4236 ( .A1(ram[3279]), .A2(n7862), .B1(n10124), .B2(n9218), .ZN(
        n7877) );
  INV_X1 U4237 ( .A(n7895), .ZN(n10074) );
  AOI22_X1 U4238 ( .A1(ram[3296]), .A2(n7896), .B1(n10090), .B2(n8858), .ZN(
        n7895) );
  INV_X1 U4239 ( .A(n7897), .ZN(n10075) );
  AOI22_X1 U4240 ( .A1(ram[3297]), .A2(n7896), .B1(n10090), .B2(n8882), .ZN(
        n7897) );
  INV_X1 U4241 ( .A(n7898), .ZN(n10076) );
  AOI22_X1 U4242 ( .A1(ram[3298]), .A2(n7896), .B1(n10090), .B2(n8906), .ZN(
        n7898) );
  INV_X1 U4243 ( .A(n7899), .ZN(n10077) );
  AOI22_X1 U4244 ( .A1(ram[3299]), .A2(n7896), .B1(n10090), .B2(n8930), .ZN(
        n7899) );
  INV_X1 U4245 ( .A(n7900), .ZN(n10078) );
  AOI22_X1 U4246 ( .A1(ram[3300]), .A2(n7896), .B1(n10090), .B2(n8954), .ZN(
        n7900) );
  INV_X1 U4247 ( .A(n7901), .ZN(n10079) );
  AOI22_X1 U4248 ( .A1(ram[3301]), .A2(n7896), .B1(n10090), .B2(n8978), .ZN(
        n7901) );
  INV_X1 U4249 ( .A(n7902), .ZN(n10080) );
  AOI22_X1 U4250 ( .A1(ram[3302]), .A2(n7896), .B1(n10090), .B2(n9002), .ZN(
        n7902) );
  INV_X1 U4251 ( .A(n7903), .ZN(n10081) );
  AOI22_X1 U4252 ( .A1(ram[3303]), .A2(n7896), .B1(n10090), .B2(n9026), .ZN(
        n7903) );
  INV_X1 U4253 ( .A(n7904), .ZN(n10082) );
  AOI22_X1 U4254 ( .A1(ram[3304]), .A2(n7896), .B1(n10090), .B2(n9050), .ZN(
        n7904) );
  INV_X1 U4255 ( .A(n7905), .ZN(n10083) );
  AOI22_X1 U4256 ( .A1(ram[3305]), .A2(n7896), .B1(n10090), .B2(n9074), .ZN(
        n7905) );
  INV_X1 U4257 ( .A(n7906), .ZN(n10084) );
  AOI22_X1 U4258 ( .A1(ram[3306]), .A2(n7896), .B1(n10090), .B2(n9098), .ZN(
        n7906) );
  INV_X1 U4259 ( .A(n7907), .ZN(n10085) );
  AOI22_X1 U4260 ( .A1(ram[3307]), .A2(n7896), .B1(n10090), .B2(n9122), .ZN(
        n7907) );
  INV_X1 U4261 ( .A(n7908), .ZN(n10086) );
  AOI22_X1 U4262 ( .A1(ram[3308]), .A2(n7896), .B1(n10090), .B2(n9146), .ZN(
        n7908) );
  INV_X1 U4263 ( .A(n7909), .ZN(n10087) );
  AOI22_X1 U4264 ( .A1(ram[3309]), .A2(n7896), .B1(n10090), .B2(n9170), .ZN(
        n7909) );
  INV_X1 U4265 ( .A(n7910), .ZN(n10088) );
  AOI22_X1 U4266 ( .A1(ram[3310]), .A2(n7896), .B1(n10090), .B2(n9194), .ZN(
        n7910) );
  INV_X1 U4267 ( .A(n7911), .ZN(n10089) );
  AOI22_X1 U4268 ( .A1(ram[3311]), .A2(n7896), .B1(n10090), .B2(n9218), .ZN(
        n7911) );
  INV_X1 U4269 ( .A(n7930), .ZN(n10040) );
  AOI22_X1 U4270 ( .A1(ram[3328]), .A2(n7931), .B1(n10056), .B2(n8857), .ZN(
        n7930) );
  INV_X1 U4271 ( .A(n7932), .ZN(n10041) );
  AOI22_X1 U4272 ( .A1(ram[3329]), .A2(n7931), .B1(n10056), .B2(n8881), .ZN(
        n7932) );
  INV_X1 U4273 ( .A(n7933), .ZN(n10042) );
  AOI22_X1 U4274 ( .A1(ram[3330]), .A2(n7931), .B1(n10056), .B2(n8905), .ZN(
        n7933) );
  INV_X1 U4275 ( .A(n7934), .ZN(n10043) );
  AOI22_X1 U4276 ( .A1(ram[3331]), .A2(n7931), .B1(n10056), .B2(n8929), .ZN(
        n7934) );
  INV_X1 U4277 ( .A(n7935), .ZN(n10044) );
  AOI22_X1 U4278 ( .A1(ram[3332]), .A2(n7931), .B1(n10056), .B2(n8953), .ZN(
        n7935) );
  INV_X1 U4279 ( .A(n7936), .ZN(n10045) );
  AOI22_X1 U4280 ( .A1(ram[3333]), .A2(n7931), .B1(n10056), .B2(n8977), .ZN(
        n7936) );
  INV_X1 U4281 ( .A(n7937), .ZN(n10046) );
  AOI22_X1 U4282 ( .A1(ram[3334]), .A2(n7931), .B1(n10056), .B2(n9001), .ZN(
        n7937) );
  INV_X1 U4283 ( .A(n7938), .ZN(n10047) );
  AOI22_X1 U4284 ( .A1(ram[3335]), .A2(n7931), .B1(n10056), .B2(n9025), .ZN(
        n7938) );
  INV_X1 U4285 ( .A(n7939), .ZN(n10048) );
  AOI22_X1 U4286 ( .A1(ram[3336]), .A2(n7931), .B1(n10056), .B2(n9049), .ZN(
        n7939) );
  INV_X1 U4287 ( .A(n7940), .ZN(n10049) );
  AOI22_X1 U4288 ( .A1(ram[3337]), .A2(n7931), .B1(n10056), .B2(n9073), .ZN(
        n7940) );
  INV_X1 U4289 ( .A(n7941), .ZN(n10050) );
  AOI22_X1 U4290 ( .A1(ram[3338]), .A2(n7931), .B1(n10056), .B2(n9097), .ZN(
        n7941) );
  INV_X1 U4291 ( .A(n7942), .ZN(n10051) );
  AOI22_X1 U4292 ( .A1(ram[3339]), .A2(n7931), .B1(n10056), .B2(n9121), .ZN(
        n7942) );
  INV_X1 U4293 ( .A(n7943), .ZN(n10052) );
  AOI22_X1 U4294 ( .A1(ram[3340]), .A2(n7931), .B1(n10056), .B2(n9145), .ZN(
        n7943) );
  INV_X1 U4295 ( .A(n7944), .ZN(n10053) );
  AOI22_X1 U4296 ( .A1(ram[3341]), .A2(n7931), .B1(n10056), .B2(n9169), .ZN(
        n7944) );
  INV_X1 U4297 ( .A(n7945), .ZN(n10054) );
  AOI22_X1 U4298 ( .A1(ram[3342]), .A2(n7931), .B1(n10056), .B2(n9193), .ZN(
        n7945) );
  INV_X1 U4299 ( .A(n7946), .ZN(n10055) );
  AOI22_X1 U4300 ( .A1(ram[3343]), .A2(n7931), .B1(n10056), .B2(n9217), .ZN(
        n7946) );
  INV_X1 U4301 ( .A(n7965), .ZN(n10006) );
  AOI22_X1 U4302 ( .A1(ram[3360]), .A2(n7966), .B1(n10022), .B2(n8857), .ZN(
        n7965) );
  INV_X1 U4303 ( .A(n7967), .ZN(n10007) );
  AOI22_X1 U4304 ( .A1(ram[3361]), .A2(n7966), .B1(n10022), .B2(n8881), .ZN(
        n7967) );
  INV_X1 U4305 ( .A(n7968), .ZN(n10008) );
  AOI22_X1 U4306 ( .A1(ram[3362]), .A2(n7966), .B1(n10022), .B2(n8905), .ZN(
        n7968) );
  INV_X1 U4307 ( .A(n7969), .ZN(n10009) );
  AOI22_X1 U4308 ( .A1(ram[3363]), .A2(n7966), .B1(n10022), .B2(n8929), .ZN(
        n7969) );
  INV_X1 U4309 ( .A(n7970), .ZN(n10010) );
  AOI22_X1 U4310 ( .A1(ram[3364]), .A2(n7966), .B1(n10022), .B2(n8953), .ZN(
        n7970) );
  INV_X1 U4311 ( .A(n7971), .ZN(n10011) );
  AOI22_X1 U4312 ( .A1(ram[3365]), .A2(n7966), .B1(n10022), .B2(n8977), .ZN(
        n7971) );
  INV_X1 U4313 ( .A(n7972), .ZN(n10012) );
  AOI22_X1 U4314 ( .A1(ram[3366]), .A2(n7966), .B1(n10022), .B2(n9001), .ZN(
        n7972) );
  INV_X1 U4315 ( .A(n7973), .ZN(n10013) );
  AOI22_X1 U4316 ( .A1(ram[3367]), .A2(n7966), .B1(n10022), .B2(n9025), .ZN(
        n7973) );
  INV_X1 U4317 ( .A(n7974), .ZN(n10014) );
  AOI22_X1 U4318 ( .A1(ram[3368]), .A2(n7966), .B1(n10022), .B2(n9049), .ZN(
        n7974) );
  INV_X1 U4319 ( .A(n7975), .ZN(n10015) );
  AOI22_X1 U4320 ( .A1(ram[3369]), .A2(n7966), .B1(n10022), .B2(n9073), .ZN(
        n7975) );
  INV_X1 U4321 ( .A(n7976), .ZN(n10016) );
  AOI22_X1 U4322 ( .A1(ram[3370]), .A2(n7966), .B1(n10022), .B2(n9097), .ZN(
        n7976) );
  INV_X1 U4323 ( .A(n7977), .ZN(n10017) );
  AOI22_X1 U4324 ( .A1(ram[3371]), .A2(n7966), .B1(n10022), .B2(n9121), .ZN(
        n7977) );
  INV_X1 U4325 ( .A(n7978), .ZN(n10018) );
  AOI22_X1 U4326 ( .A1(ram[3372]), .A2(n7966), .B1(n10022), .B2(n9145), .ZN(
        n7978) );
  INV_X1 U4327 ( .A(n7979), .ZN(n10019) );
  AOI22_X1 U4328 ( .A1(ram[3373]), .A2(n7966), .B1(n10022), .B2(n9169), .ZN(
        n7979) );
  INV_X1 U4329 ( .A(n7980), .ZN(n10020) );
  AOI22_X1 U4330 ( .A1(ram[3374]), .A2(n7966), .B1(n10022), .B2(n9193), .ZN(
        n7980) );
  INV_X1 U4331 ( .A(n7981), .ZN(n10021) );
  AOI22_X1 U4332 ( .A1(ram[3375]), .A2(n7966), .B1(n10022), .B2(n9217), .ZN(
        n7981) );
  INV_X1 U4333 ( .A(n7999), .ZN(n9972) );
  AOI22_X1 U4334 ( .A1(ram[3392]), .A2(n8000), .B1(n9988), .B2(n8857), .ZN(
        n7999) );
  INV_X1 U4335 ( .A(n8001), .ZN(n9973) );
  AOI22_X1 U4336 ( .A1(ram[3393]), .A2(n8000), .B1(n9988), .B2(n8881), .ZN(
        n8001) );
  INV_X1 U4337 ( .A(n8002), .ZN(n9974) );
  AOI22_X1 U4338 ( .A1(ram[3394]), .A2(n8000), .B1(n9988), .B2(n8905), .ZN(
        n8002) );
  INV_X1 U4339 ( .A(n8003), .ZN(n9975) );
  AOI22_X1 U4340 ( .A1(ram[3395]), .A2(n8000), .B1(n9988), .B2(n8929), .ZN(
        n8003) );
  INV_X1 U4341 ( .A(n8004), .ZN(n9976) );
  AOI22_X1 U4342 ( .A1(ram[3396]), .A2(n8000), .B1(n9988), .B2(n8953), .ZN(
        n8004) );
  INV_X1 U4343 ( .A(n8005), .ZN(n9977) );
  AOI22_X1 U4344 ( .A1(ram[3397]), .A2(n8000), .B1(n9988), .B2(n8977), .ZN(
        n8005) );
  INV_X1 U4345 ( .A(n8006), .ZN(n9978) );
  AOI22_X1 U4346 ( .A1(ram[3398]), .A2(n8000), .B1(n9988), .B2(n9001), .ZN(
        n8006) );
  INV_X1 U4347 ( .A(n8007), .ZN(n9979) );
  AOI22_X1 U4348 ( .A1(ram[3399]), .A2(n8000), .B1(n9988), .B2(n9025), .ZN(
        n8007) );
  INV_X1 U4349 ( .A(n8008), .ZN(n9980) );
  AOI22_X1 U4350 ( .A1(ram[3400]), .A2(n8000), .B1(n9988), .B2(n9049), .ZN(
        n8008) );
  INV_X1 U4351 ( .A(n8009), .ZN(n9981) );
  AOI22_X1 U4352 ( .A1(ram[3401]), .A2(n8000), .B1(n9988), .B2(n9073), .ZN(
        n8009) );
  INV_X1 U4353 ( .A(n8010), .ZN(n9982) );
  AOI22_X1 U4354 ( .A1(ram[3402]), .A2(n8000), .B1(n9988), .B2(n9097), .ZN(
        n8010) );
  INV_X1 U4355 ( .A(n8011), .ZN(n9983) );
  AOI22_X1 U4356 ( .A1(ram[3403]), .A2(n8000), .B1(n9988), .B2(n9121), .ZN(
        n8011) );
  INV_X1 U4357 ( .A(n8012), .ZN(n9984) );
  AOI22_X1 U4358 ( .A1(ram[3404]), .A2(n8000), .B1(n9988), .B2(n9145), .ZN(
        n8012) );
  INV_X1 U4359 ( .A(n8013), .ZN(n9985) );
  AOI22_X1 U4360 ( .A1(ram[3405]), .A2(n8000), .B1(n9988), .B2(n9169), .ZN(
        n8013) );
  INV_X1 U4361 ( .A(n8014), .ZN(n9986) );
  AOI22_X1 U4362 ( .A1(ram[3406]), .A2(n8000), .B1(n9988), .B2(n9193), .ZN(
        n8014) );
  INV_X1 U4363 ( .A(n8015), .ZN(n9987) );
  AOI22_X1 U4364 ( .A1(ram[3407]), .A2(n8000), .B1(n9988), .B2(n9217), .ZN(
        n8015) );
  INV_X1 U4365 ( .A(n8033), .ZN(n9938) );
  AOI22_X1 U4366 ( .A1(ram[3424]), .A2(n8034), .B1(n9954), .B2(n8857), .ZN(
        n8033) );
  INV_X1 U4367 ( .A(n8035), .ZN(n9939) );
  AOI22_X1 U4368 ( .A1(ram[3425]), .A2(n8034), .B1(n9954), .B2(n8881), .ZN(
        n8035) );
  INV_X1 U4369 ( .A(n8036), .ZN(n9940) );
  AOI22_X1 U4370 ( .A1(ram[3426]), .A2(n8034), .B1(n9954), .B2(n8905), .ZN(
        n8036) );
  INV_X1 U4371 ( .A(n8037), .ZN(n9941) );
  AOI22_X1 U4372 ( .A1(ram[3427]), .A2(n8034), .B1(n9954), .B2(n8929), .ZN(
        n8037) );
  INV_X1 U4373 ( .A(n8038), .ZN(n9942) );
  AOI22_X1 U4374 ( .A1(ram[3428]), .A2(n8034), .B1(n9954), .B2(n8953), .ZN(
        n8038) );
  INV_X1 U4375 ( .A(n8039), .ZN(n9943) );
  AOI22_X1 U4376 ( .A1(ram[3429]), .A2(n8034), .B1(n9954), .B2(n8977), .ZN(
        n8039) );
  INV_X1 U4377 ( .A(n8040), .ZN(n9944) );
  AOI22_X1 U4378 ( .A1(ram[3430]), .A2(n8034), .B1(n9954), .B2(n9001), .ZN(
        n8040) );
  INV_X1 U4379 ( .A(n8041), .ZN(n9945) );
  AOI22_X1 U4380 ( .A1(ram[3431]), .A2(n8034), .B1(n9954), .B2(n9025), .ZN(
        n8041) );
  INV_X1 U4381 ( .A(n8042), .ZN(n9946) );
  AOI22_X1 U4382 ( .A1(ram[3432]), .A2(n8034), .B1(n9954), .B2(n9049), .ZN(
        n8042) );
  INV_X1 U4383 ( .A(n8043), .ZN(n9947) );
  AOI22_X1 U4384 ( .A1(ram[3433]), .A2(n8034), .B1(n9954), .B2(n9073), .ZN(
        n8043) );
  INV_X1 U4385 ( .A(n8044), .ZN(n9948) );
  AOI22_X1 U4386 ( .A1(ram[3434]), .A2(n8034), .B1(n9954), .B2(n9097), .ZN(
        n8044) );
  INV_X1 U4387 ( .A(n8045), .ZN(n9949) );
  AOI22_X1 U4388 ( .A1(ram[3435]), .A2(n8034), .B1(n9954), .B2(n9121), .ZN(
        n8045) );
  INV_X1 U4389 ( .A(n8046), .ZN(n9950) );
  AOI22_X1 U4390 ( .A1(ram[3436]), .A2(n8034), .B1(n9954), .B2(n9145), .ZN(
        n8046) );
  INV_X1 U4391 ( .A(n8047), .ZN(n9951) );
  AOI22_X1 U4392 ( .A1(ram[3437]), .A2(n8034), .B1(n9954), .B2(n9169), .ZN(
        n8047) );
  INV_X1 U4393 ( .A(n8048), .ZN(n9952) );
  AOI22_X1 U4394 ( .A1(ram[3438]), .A2(n8034), .B1(n9954), .B2(n9193), .ZN(
        n8048) );
  INV_X1 U4395 ( .A(n8049), .ZN(n9953) );
  AOI22_X1 U4396 ( .A1(ram[3439]), .A2(n8034), .B1(n9954), .B2(n9217), .ZN(
        n8049) );
  INV_X1 U4397 ( .A(n8067), .ZN(n9904) );
  AOI22_X1 U4398 ( .A1(ram[3456]), .A2(n8068), .B1(n9920), .B2(n8857), .ZN(
        n8067) );
  INV_X1 U4399 ( .A(n8069), .ZN(n9905) );
  AOI22_X1 U4400 ( .A1(ram[3457]), .A2(n8068), .B1(n9920), .B2(n8881), .ZN(
        n8069) );
  INV_X1 U4401 ( .A(n8070), .ZN(n9906) );
  AOI22_X1 U4402 ( .A1(ram[3458]), .A2(n8068), .B1(n9920), .B2(n8905), .ZN(
        n8070) );
  INV_X1 U4403 ( .A(n8071), .ZN(n9907) );
  AOI22_X1 U4404 ( .A1(ram[3459]), .A2(n8068), .B1(n9920), .B2(n8929), .ZN(
        n8071) );
  INV_X1 U4405 ( .A(n8072), .ZN(n9908) );
  AOI22_X1 U4406 ( .A1(ram[3460]), .A2(n8068), .B1(n9920), .B2(n8953), .ZN(
        n8072) );
  INV_X1 U4407 ( .A(n8073), .ZN(n9909) );
  AOI22_X1 U4408 ( .A1(ram[3461]), .A2(n8068), .B1(n9920), .B2(n8977), .ZN(
        n8073) );
  INV_X1 U4409 ( .A(n8074), .ZN(n9910) );
  AOI22_X1 U4410 ( .A1(ram[3462]), .A2(n8068), .B1(n9920), .B2(n9001), .ZN(
        n8074) );
  INV_X1 U4411 ( .A(n8075), .ZN(n9911) );
  AOI22_X1 U4412 ( .A1(ram[3463]), .A2(n8068), .B1(n9920), .B2(n9025), .ZN(
        n8075) );
  INV_X1 U4413 ( .A(n8076), .ZN(n9912) );
  AOI22_X1 U4414 ( .A1(ram[3464]), .A2(n8068), .B1(n9920), .B2(n9049), .ZN(
        n8076) );
  INV_X1 U4415 ( .A(n8077), .ZN(n9913) );
  AOI22_X1 U4416 ( .A1(ram[3465]), .A2(n8068), .B1(n9920), .B2(n9073), .ZN(
        n8077) );
  INV_X1 U4417 ( .A(n8078), .ZN(n9914) );
  AOI22_X1 U4418 ( .A1(ram[3466]), .A2(n8068), .B1(n9920), .B2(n9097), .ZN(
        n8078) );
  INV_X1 U4419 ( .A(n8079), .ZN(n9915) );
  AOI22_X1 U4420 ( .A1(ram[3467]), .A2(n8068), .B1(n9920), .B2(n9121), .ZN(
        n8079) );
  INV_X1 U4421 ( .A(n8080), .ZN(n9916) );
  AOI22_X1 U4422 ( .A1(ram[3468]), .A2(n8068), .B1(n9920), .B2(n9145), .ZN(
        n8080) );
  INV_X1 U4423 ( .A(n8081), .ZN(n9917) );
  AOI22_X1 U4424 ( .A1(ram[3469]), .A2(n8068), .B1(n9920), .B2(n9169), .ZN(
        n8081) );
  INV_X1 U4425 ( .A(n8082), .ZN(n9918) );
  AOI22_X1 U4426 ( .A1(ram[3470]), .A2(n8068), .B1(n9920), .B2(n9193), .ZN(
        n8082) );
  INV_X1 U4427 ( .A(n8083), .ZN(n9919) );
  AOI22_X1 U4428 ( .A1(ram[3471]), .A2(n8068), .B1(n9920), .B2(n9217), .ZN(
        n8083) );
  INV_X1 U4429 ( .A(n8101), .ZN(n9870) );
  AOI22_X1 U4430 ( .A1(ram[3488]), .A2(n8102), .B1(n9886), .B2(n8857), .ZN(
        n8101) );
  INV_X1 U4431 ( .A(n8103), .ZN(n9871) );
  AOI22_X1 U4432 ( .A1(ram[3489]), .A2(n8102), .B1(n9886), .B2(n8881), .ZN(
        n8103) );
  INV_X1 U4433 ( .A(n8104), .ZN(n9872) );
  AOI22_X1 U4434 ( .A1(ram[3490]), .A2(n8102), .B1(n9886), .B2(n8905), .ZN(
        n8104) );
  INV_X1 U4435 ( .A(n8105), .ZN(n9873) );
  AOI22_X1 U4436 ( .A1(ram[3491]), .A2(n8102), .B1(n9886), .B2(n8929), .ZN(
        n8105) );
  INV_X1 U4437 ( .A(n8106), .ZN(n9874) );
  AOI22_X1 U4438 ( .A1(ram[3492]), .A2(n8102), .B1(n9886), .B2(n8953), .ZN(
        n8106) );
  INV_X1 U4439 ( .A(n8107), .ZN(n9875) );
  AOI22_X1 U4440 ( .A1(ram[3493]), .A2(n8102), .B1(n9886), .B2(n8977), .ZN(
        n8107) );
  INV_X1 U4441 ( .A(n8108), .ZN(n9876) );
  AOI22_X1 U4442 ( .A1(ram[3494]), .A2(n8102), .B1(n9886), .B2(n9001), .ZN(
        n8108) );
  INV_X1 U4443 ( .A(n8109), .ZN(n9877) );
  AOI22_X1 U4444 ( .A1(ram[3495]), .A2(n8102), .B1(n9886), .B2(n9025), .ZN(
        n8109) );
  INV_X1 U4445 ( .A(n8110), .ZN(n9878) );
  AOI22_X1 U4446 ( .A1(ram[3496]), .A2(n8102), .B1(n9886), .B2(n9049), .ZN(
        n8110) );
  INV_X1 U4447 ( .A(n8111), .ZN(n9879) );
  AOI22_X1 U4448 ( .A1(ram[3497]), .A2(n8102), .B1(n9886), .B2(n9073), .ZN(
        n8111) );
  INV_X1 U4449 ( .A(n8112), .ZN(n9880) );
  AOI22_X1 U4450 ( .A1(ram[3498]), .A2(n8102), .B1(n9886), .B2(n9097), .ZN(
        n8112) );
  INV_X1 U4451 ( .A(n8113), .ZN(n9881) );
  AOI22_X1 U4452 ( .A1(ram[3499]), .A2(n8102), .B1(n9886), .B2(n9121), .ZN(
        n8113) );
  INV_X1 U4453 ( .A(n8114), .ZN(n9882) );
  AOI22_X1 U4454 ( .A1(ram[3500]), .A2(n8102), .B1(n9886), .B2(n9145), .ZN(
        n8114) );
  INV_X1 U4455 ( .A(n8115), .ZN(n9883) );
  AOI22_X1 U4456 ( .A1(ram[3501]), .A2(n8102), .B1(n9886), .B2(n9169), .ZN(
        n8115) );
  INV_X1 U4457 ( .A(n8116), .ZN(n9884) );
  AOI22_X1 U4458 ( .A1(ram[3502]), .A2(n8102), .B1(n9886), .B2(n9193), .ZN(
        n8116) );
  INV_X1 U4459 ( .A(n8117), .ZN(n9885) );
  AOI22_X1 U4460 ( .A1(ram[3503]), .A2(n8102), .B1(n9886), .B2(n9217), .ZN(
        n8117) );
  INV_X1 U4461 ( .A(n8135), .ZN(n9836) );
  AOI22_X1 U4462 ( .A1(ram[3520]), .A2(n8136), .B1(n9852), .B2(n8856), .ZN(
        n8135) );
  INV_X1 U4463 ( .A(n8137), .ZN(n9837) );
  AOI22_X1 U4464 ( .A1(ram[3521]), .A2(n8136), .B1(n9852), .B2(n8880), .ZN(
        n8137) );
  INV_X1 U4465 ( .A(n8138), .ZN(n9838) );
  AOI22_X1 U4466 ( .A1(ram[3522]), .A2(n8136), .B1(n9852), .B2(n8904), .ZN(
        n8138) );
  INV_X1 U4467 ( .A(n8139), .ZN(n9839) );
  AOI22_X1 U4468 ( .A1(ram[3523]), .A2(n8136), .B1(n9852), .B2(n8928), .ZN(
        n8139) );
  INV_X1 U4469 ( .A(n8140), .ZN(n9840) );
  AOI22_X1 U4470 ( .A1(ram[3524]), .A2(n8136), .B1(n9852), .B2(n8952), .ZN(
        n8140) );
  INV_X1 U4471 ( .A(n8141), .ZN(n9841) );
  AOI22_X1 U4472 ( .A1(ram[3525]), .A2(n8136), .B1(n9852), .B2(n8976), .ZN(
        n8141) );
  INV_X1 U4473 ( .A(n8142), .ZN(n9842) );
  AOI22_X1 U4474 ( .A1(ram[3526]), .A2(n8136), .B1(n9852), .B2(n9000), .ZN(
        n8142) );
  INV_X1 U4475 ( .A(n8143), .ZN(n9843) );
  AOI22_X1 U4476 ( .A1(ram[3527]), .A2(n8136), .B1(n9852), .B2(n9024), .ZN(
        n8143) );
  INV_X1 U4477 ( .A(n8144), .ZN(n9844) );
  AOI22_X1 U4478 ( .A1(ram[3528]), .A2(n8136), .B1(n9852), .B2(n9048), .ZN(
        n8144) );
  INV_X1 U4479 ( .A(n8145), .ZN(n9845) );
  AOI22_X1 U4480 ( .A1(ram[3529]), .A2(n8136), .B1(n9852), .B2(n9072), .ZN(
        n8145) );
  INV_X1 U4481 ( .A(n8146), .ZN(n9846) );
  AOI22_X1 U4482 ( .A1(ram[3530]), .A2(n8136), .B1(n9852), .B2(n9096), .ZN(
        n8146) );
  INV_X1 U4483 ( .A(n8147), .ZN(n9847) );
  AOI22_X1 U4484 ( .A1(ram[3531]), .A2(n8136), .B1(n9852), .B2(n9120), .ZN(
        n8147) );
  INV_X1 U4485 ( .A(n8148), .ZN(n9848) );
  AOI22_X1 U4486 ( .A1(ram[3532]), .A2(n8136), .B1(n9852), .B2(n9144), .ZN(
        n8148) );
  INV_X1 U4487 ( .A(n8149), .ZN(n9849) );
  AOI22_X1 U4488 ( .A1(ram[3533]), .A2(n8136), .B1(n9852), .B2(n9168), .ZN(
        n8149) );
  INV_X1 U4489 ( .A(n8150), .ZN(n9850) );
  AOI22_X1 U4490 ( .A1(ram[3534]), .A2(n8136), .B1(n9852), .B2(n9192), .ZN(
        n8150) );
  INV_X1 U4491 ( .A(n8151), .ZN(n9851) );
  AOI22_X1 U4492 ( .A1(ram[3535]), .A2(n8136), .B1(n9852), .B2(n9216), .ZN(
        n8151) );
  INV_X1 U4493 ( .A(n8169), .ZN(n9802) );
  AOI22_X1 U4494 ( .A1(ram[3552]), .A2(n8170), .B1(n9818), .B2(n8856), .ZN(
        n8169) );
  INV_X1 U4495 ( .A(n8171), .ZN(n9803) );
  AOI22_X1 U4496 ( .A1(ram[3553]), .A2(n8170), .B1(n9818), .B2(n8880), .ZN(
        n8171) );
  INV_X1 U4497 ( .A(n8172), .ZN(n9804) );
  AOI22_X1 U4498 ( .A1(ram[3554]), .A2(n8170), .B1(n9818), .B2(n8904), .ZN(
        n8172) );
  INV_X1 U4499 ( .A(n8173), .ZN(n9805) );
  AOI22_X1 U4500 ( .A1(ram[3555]), .A2(n8170), .B1(n9818), .B2(n8928), .ZN(
        n8173) );
  INV_X1 U4501 ( .A(n8174), .ZN(n9806) );
  AOI22_X1 U4502 ( .A1(ram[3556]), .A2(n8170), .B1(n9818), .B2(n8952), .ZN(
        n8174) );
  INV_X1 U4503 ( .A(n8175), .ZN(n9807) );
  AOI22_X1 U4504 ( .A1(ram[3557]), .A2(n8170), .B1(n9818), .B2(n8976), .ZN(
        n8175) );
  INV_X1 U4505 ( .A(n8176), .ZN(n9808) );
  AOI22_X1 U4506 ( .A1(ram[3558]), .A2(n8170), .B1(n9818), .B2(n9000), .ZN(
        n8176) );
  INV_X1 U4507 ( .A(n8177), .ZN(n9809) );
  AOI22_X1 U4508 ( .A1(ram[3559]), .A2(n8170), .B1(n9818), .B2(n9024), .ZN(
        n8177) );
  INV_X1 U4509 ( .A(n8178), .ZN(n9810) );
  AOI22_X1 U4510 ( .A1(ram[3560]), .A2(n8170), .B1(n9818), .B2(n9048), .ZN(
        n8178) );
  INV_X1 U4511 ( .A(n8179), .ZN(n9811) );
  AOI22_X1 U4512 ( .A1(ram[3561]), .A2(n8170), .B1(n9818), .B2(n9072), .ZN(
        n8179) );
  INV_X1 U4513 ( .A(n8180), .ZN(n9812) );
  AOI22_X1 U4514 ( .A1(ram[3562]), .A2(n8170), .B1(n9818), .B2(n9096), .ZN(
        n8180) );
  INV_X1 U4515 ( .A(n8181), .ZN(n9813) );
  AOI22_X1 U4516 ( .A1(ram[3563]), .A2(n8170), .B1(n9818), .B2(n9120), .ZN(
        n8181) );
  INV_X1 U4517 ( .A(n8182), .ZN(n9814) );
  AOI22_X1 U4518 ( .A1(ram[3564]), .A2(n8170), .B1(n9818), .B2(n9144), .ZN(
        n8182) );
  INV_X1 U4519 ( .A(n8183), .ZN(n9815) );
  AOI22_X1 U4520 ( .A1(ram[3565]), .A2(n8170), .B1(n9818), .B2(n9168), .ZN(
        n8183) );
  INV_X1 U4521 ( .A(n8184), .ZN(n9816) );
  AOI22_X1 U4522 ( .A1(ram[3566]), .A2(n8170), .B1(n9818), .B2(n9192), .ZN(
        n8184) );
  INV_X1 U4523 ( .A(n8185), .ZN(n9817) );
  AOI22_X1 U4524 ( .A1(ram[3567]), .A2(n8170), .B1(n9818), .B2(n9216), .ZN(
        n8185) );
  INV_X1 U4525 ( .A(n8203), .ZN(n9768) );
  AOI22_X1 U4526 ( .A1(ram[3584]), .A2(n8204), .B1(n9784), .B2(n8856), .ZN(
        n8203) );
  INV_X1 U4527 ( .A(n8205), .ZN(n9769) );
  AOI22_X1 U4528 ( .A1(ram[3585]), .A2(n8204), .B1(n9784), .B2(n8880), .ZN(
        n8205) );
  INV_X1 U4529 ( .A(n8206), .ZN(n9770) );
  AOI22_X1 U4530 ( .A1(ram[3586]), .A2(n8204), .B1(n9784), .B2(n8904), .ZN(
        n8206) );
  INV_X1 U4531 ( .A(n8207), .ZN(n9771) );
  AOI22_X1 U4532 ( .A1(ram[3587]), .A2(n8204), .B1(n9784), .B2(n8928), .ZN(
        n8207) );
  INV_X1 U4533 ( .A(n8208), .ZN(n9772) );
  AOI22_X1 U4534 ( .A1(ram[3588]), .A2(n8204), .B1(n9784), .B2(n8952), .ZN(
        n8208) );
  INV_X1 U4535 ( .A(n8209), .ZN(n9773) );
  AOI22_X1 U4536 ( .A1(ram[3589]), .A2(n8204), .B1(n9784), .B2(n8976), .ZN(
        n8209) );
  INV_X1 U4537 ( .A(n8210), .ZN(n9774) );
  AOI22_X1 U4538 ( .A1(ram[3590]), .A2(n8204), .B1(n9784), .B2(n9000), .ZN(
        n8210) );
  INV_X1 U4539 ( .A(n8211), .ZN(n9775) );
  AOI22_X1 U4540 ( .A1(ram[3591]), .A2(n8204), .B1(n9784), .B2(n9024), .ZN(
        n8211) );
  INV_X1 U4541 ( .A(n8212), .ZN(n9776) );
  AOI22_X1 U4542 ( .A1(ram[3592]), .A2(n8204), .B1(n9784), .B2(n9048), .ZN(
        n8212) );
  INV_X1 U4543 ( .A(n8213), .ZN(n9777) );
  AOI22_X1 U4544 ( .A1(ram[3593]), .A2(n8204), .B1(n9784), .B2(n9072), .ZN(
        n8213) );
  INV_X1 U4545 ( .A(n8214), .ZN(n9778) );
  AOI22_X1 U4546 ( .A1(ram[3594]), .A2(n8204), .B1(n9784), .B2(n9096), .ZN(
        n8214) );
  INV_X1 U4547 ( .A(n8215), .ZN(n9779) );
  AOI22_X1 U4548 ( .A1(ram[3595]), .A2(n8204), .B1(n9784), .B2(n9120), .ZN(
        n8215) );
  INV_X1 U4549 ( .A(n8216), .ZN(n9780) );
  AOI22_X1 U4550 ( .A1(ram[3596]), .A2(n8204), .B1(n9784), .B2(n9144), .ZN(
        n8216) );
  INV_X1 U4551 ( .A(n8217), .ZN(n9781) );
  AOI22_X1 U4552 ( .A1(ram[3597]), .A2(n8204), .B1(n9784), .B2(n9168), .ZN(
        n8217) );
  INV_X1 U4553 ( .A(n8218), .ZN(n9782) );
  AOI22_X1 U4554 ( .A1(ram[3598]), .A2(n8204), .B1(n9784), .B2(n9192), .ZN(
        n8218) );
  INV_X1 U4555 ( .A(n8219), .ZN(n9783) );
  AOI22_X1 U4556 ( .A1(ram[3599]), .A2(n8204), .B1(n9784), .B2(n9216), .ZN(
        n8219) );
  INV_X1 U4557 ( .A(n8238), .ZN(n9734) );
  AOI22_X1 U4558 ( .A1(ram[3616]), .A2(n8239), .B1(n9750), .B2(n8856), .ZN(
        n8238) );
  INV_X1 U4559 ( .A(n8240), .ZN(n9735) );
  AOI22_X1 U4560 ( .A1(ram[3617]), .A2(n8239), .B1(n9750), .B2(n8880), .ZN(
        n8240) );
  INV_X1 U4561 ( .A(n8241), .ZN(n9736) );
  AOI22_X1 U4562 ( .A1(ram[3618]), .A2(n8239), .B1(n9750), .B2(n8904), .ZN(
        n8241) );
  INV_X1 U4563 ( .A(n8242), .ZN(n9737) );
  AOI22_X1 U4564 ( .A1(ram[3619]), .A2(n8239), .B1(n9750), .B2(n8928), .ZN(
        n8242) );
  INV_X1 U4565 ( .A(n8243), .ZN(n9738) );
  AOI22_X1 U4566 ( .A1(ram[3620]), .A2(n8239), .B1(n9750), .B2(n8952), .ZN(
        n8243) );
  INV_X1 U4567 ( .A(n8244), .ZN(n9739) );
  AOI22_X1 U4568 ( .A1(ram[3621]), .A2(n8239), .B1(n9750), .B2(n8976), .ZN(
        n8244) );
  INV_X1 U4569 ( .A(n8245), .ZN(n9740) );
  AOI22_X1 U4570 ( .A1(ram[3622]), .A2(n8239), .B1(n9750), .B2(n9000), .ZN(
        n8245) );
  INV_X1 U4571 ( .A(n8246), .ZN(n9741) );
  AOI22_X1 U4572 ( .A1(ram[3623]), .A2(n8239), .B1(n9750), .B2(n9024), .ZN(
        n8246) );
  INV_X1 U4573 ( .A(n8247), .ZN(n9742) );
  AOI22_X1 U4574 ( .A1(ram[3624]), .A2(n8239), .B1(n9750), .B2(n9048), .ZN(
        n8247) );
  INV_X1 U4575 ( .A(n8248), .ZN(n9743) );
  AOI22_X1 U4576 ( .A1(ram[3625]), .A2(n8239), .B1(n9750), .B2(n9072), .ZN(
        n8248) );
  INV_X1 U4577 ( .A(n8249), .ZN(n9744) );
  AOI22_X1 U4578 ( .A1(ram[3626]), .A2(n8239), .B1(n9750), .B2(n9096), .ZN(
        n8249) );
  INV_X1 U4579 ( .A(n8250), .ZN(n9745) );
  AOI22_X1 U4580 ( .A1(ram[3627]), .A2(n8239), .B1(n9750), .B2(n9120), .ZN(
        n8250) );
  INV_X1 U4581 ( .A(n8251), .ZN(n9746) );
  AOI22_X1 U4582 ( .A1(ram[3628]), .A2(n8239), .B1(n9750), .B2(n9144), .ZN(
        n8251) );
  INV_X1 U4583 ( .A(n8252), .ZN(n9747) );
  AOI22_X1 U4584 ( .A1(ram[3629]), .A2(n8239), .B1(n9750), .B2(n9168), .ZN(
        n8252) );
  INV_X1 U4585 ( .A(n8253), .ZN(n9748) );
  AOI22_X1 U4586 ( .A1(ram[3630]), .A2(n8239), .B1(n9750), .B2(n9192), .ZN(
        n8253) );
  INV_X1 U4587 ( .A(n8254), .ZN(n9749) );
  AOI22_X1 U4588 ( .A1(ram[3631]), .A2(n8239), .B1(n9750), .B2(n9216), .ZN(
        n8254) );
  INV_X1 U4589 ( .A(n8272), .ZN(n9700) );
  AOI22_X1 U4590 ( .A1(ram[3648]), .A2(n8273), .B1(n9716), .B2(n8856), .ZN(
        n8272) );
  INV_X1 U4591 ( .A(n8274), .ZN(n9701) );
  AOI22_X1 U4592 ( .A1(ram[3649]), .A2(n8273), .B1(n9716), .B2(n8880), .ZN(
        n8274) );
  INV_X1 U4593 ( .A(n8275), .ZN(n9702) );
  AOI22_X1 U4594 ( .A1(ram[3650]), .A2(n8273), .B1(n9716), .B2(n8904), .ZN(
        n8275) );
  INV_X1 U4595 ( .A(n8276), .ZN(n9703) );
  AOI22_X1 U4596 ( .A1(ram[3651]), .A2(n8273), .B1(n9716), .B2(n8928), .ZN(
        n8276) );
  INV_X1 U4597 ( .A(n8277), .ZN(n9704) );
  AOI22_X1 U4598 ( .A1(ram[3652]), .A2(n8273), .B1(n9716), .B2(n8952), .ZN(
        n8277) );
  INV_X1 U4599 ( .A(n8278), .ZN(n9705) );
  AOI22_X1 U4600 ( .A1(ram[3653]), .A2(n8273), .B1(n9716), .B2(n8976), .ZN(
        n8278) );
  INV_X1 U4601 ( .A(n8279), .ZN(n9706) );
  AOI22_X1 U4602 ( .A1(ram[3654]), .A2(n8273), .B1(n9716), .B2(n9000), .ZN(
        n8279) );
  INV_X1 U4603 ( .A(n8280), .ZN(n9707) );
  AOI22_X1 U4604 ( .A1(ram[3655]), .A2(n8273), .B1(n9716), .B2(n9024), .ZN(
        n8280) );
  INV_X1 U4605 ( .A(n8281), .ZN(n9708) );
  AOI22_X1 U4606 ( .A1(ram[3656]), .A2(n8273), .B1(n9716), .B2(n9048), .ZN(
        n8281) );
  INV_X1 U4607 ( .A(n8282), .ZN(n9709) );
  AOI22_X1 U4608 ( .A1(ram[3657]), .A2(n8273), .B1(n9716), .B2(n9072), .ZN(
        n8282) );
  INV_X1 U4609 ( .A(n8283), .ZN(n9710) );
  AOI22_X1 U4610 ( .A1(ram[3658]), .A2(n8273), .B1(n9716), .B2(n9096), .ZN(
        n8283) );
  INV_X1 U4611 ( .A(n8284), .ZN(n9711) );
  AOI22_X1 U4612 ( .A1(ram[3659]), .A2(n8273), .B1(n9716), .B2(n9120), .ZN(
        n8284) );
  INV_X1 U4613 ( .A(n8285), .ZN(n9712) );
  AOI22_X1 U4614 ( .A1(ram[3660]), .A2(n8273), .B1(n9716), .B2(n9144), .ZN(
        n8285) );
  INV_X1 U4615 ( .A(n8286), .ZN(n9713) );
  AOI22_X1 U4616 ( .A1(ram[3661]), .A2(n8273), .B1(n9716), .B2(n9168), .ZN(
        n8286) );
  INV_X1 U4617 ( .A(n8287), .ZN(n9714) );
  AOI22_X1 U4618 ( .A1(ram[3662]), .A2(n8273), .B1(n9716), .B2(n9192), .ZN(
        n8287) );
  INV_X1 U4619 ( .A(n8288), .ZN(n9715) );
  AOI22_X1 U4620 ( .A1(ram[3663]), .A2(n8273), .B1(n9716), .B2(n9216), .ZN(
        n8288) );
  INV_X1 U4621 ( .A(n8306), .ZN(n9666) );
  AOI22_X1 U4622 ( .A1(ram[3680]), .A2(n8307), .B1(n9682), .B2(n8856), .ZN(
        n8306) );
  INV_X1 U4623 ( .A(n8308), .ZN(n9667) );
  AOI22_X1 U4624 ( .A1(ram[3681]), .A2(n8307), .B1(n9682), .B2(n8880), .ZN(
        n8308) );
  INV_X1 U4625 ( .A(n8309), .ZN(n9668) );
  AOI22_X1 U4626 ( .A1(ram[3682]), .A2(n8307), .B1(n9682), .B2(n8904), .ZN(
        n8309) );
  INV_X1 U4627 ( .A(n8310), .ZN(n9669) );
  AOI22_X1 U4628 ( .A1(ram[3683]), .A2(n8307), .B1(n9682), .B2(n8928), .ZN(
        n8310) );
  INV_X1 U4629 ( .A(n8311), .ZN(n9670) );
  AOI22_X1 U4630 ( .A1(ram[3684]), .A2(n8307), .B1(n9682), .B2(n8952), .ZN(
        n8311) );
  INV_X1 U4631 ( .A(n8312), .ZN(n9671) );
  AOI22_X1 U4632 ( .A1(ram[3685]), .A2(n8307), .B1(n9682), .B2(n8976), .ZN(
        n8312) );
  INV_X1 U4633 ( .A(n8313), .ZN(n9672) );
  AOI22_X1 U4634 ( .A1(ram[3686]), .A2(n8307), .B1(n9682), .B2(n9000), .ZN(
        n8313) );
  INV_X1 U4635 ( .A(n8314), .ZN(n9673) );
  AOI22_X1 U4636 ( .A1(ram[3687]), .A2(n8307), .B1(n9682), .B2(n9024), .ZN(
        n8314) );
  INV_X1 U4637 ( .A(n8315), .ZN(n9674) );
  AOI22_X1 U4638 ( .A1(ram[3688]), .A2(n8307), .B1(n9682), .B2(n9048), .ZN(
        n8315) );
  INV_X1 U4639 ( .A(n8316), .ZN(n9675) );
  AOI22_X1 U4640 ( .A1(ram[3689]), .A2(n8307), .B1(n9682), .B2(n9072), .ZN(
        n8316) );
  INV_X1 U4641 ( .A(n8317), .ZN(n9676) );
  AOI22_X1 U4642 ( .A1(ram[3690]), .A2(n8307), .B1(n9682), .B2(n9096), .ZN(
        n8317) );
  INV_X1 U4643 ( .A(n8318), .ZN(n9677) );
  AOI22_X1 U4644 ( .A1(ram[3691]), .A2(n8307), .B1(n9682), .B2(n9120), .ZN(
        n8318) );
  INV_X1 U4645 ( .A(n8319), .ZN(n9678) );
  AOI22_X1 U4646 ( .A1(ram[3692]), .A2(n8307), .B1(n9682), .B2(n9144), .ZN(
        n8319) );
  INV_X1 U4647 ( .A(n8320), .ZN(n9679) );
  AOI22_X1 U4648 ( .A1(ram[3693]), .A2(n8307), .B1(n9682), .B2(n9168), .ZN(
        n8320) );
  INV_X1 U4649 ( .A(n8321), .ZN(n9680) );
  AOI22_X1 U4650 ( .A1(ram[3694]), .A2(n8307), .B1(n9682), .B2(n9192), .ZN(
        n8321) );
  INV_X1 U4651 ( .A(n8322), .ZN(n9681) );
  AOI22_X1 U4652 ( .A1(ram[3695]), .A2(n8307), .B1(n9682), .B2(n9216), .ZN(
        n8322) );
  INV_X1 U4653 ( .A(n8340), .ZN(n9632) );
  AOI22_X1 U4654 ( .A1(ram[3712]), .A2(n8341), .B1(n9648), .B2(n8855), .ZN(
        n8340) );
  INV_X1 U4655 ( .A(n8342), .ZN(n9633) );
  AOI22_X1 U4656 ( .A1(ram[3713]), .A2(n8341), .B1(n9648), .B2(n8879), .ZN(
        n8342) );
  INV_X1 U4657 ( .A(n8343), .ZN(n9634) );
  AOI22_X1 U4658 ( .A1(ram[3714]), .A2(n8341), .B1(n9648), .B2(n8903), .ZN(
        n8343) );
  INV_X1 U4659 ( .A(n8344), .ZN(n9635) );
  AOI22_X1 U4660 ( .A1(ram[3715]), .A2(n8341), .B1(n9648), .B2(n8927), .ZN(
        n8344) );
  INV_X1 U4661 ( .A(n8345), .ZN(n9636) );
  AOI22_X1 U4662 ( .A1(ram[3716]), .A2(n8341), .B1(n9648), .B2(n8951), .ZN(
        n8345) );
  INV_X1 U4663 ( .A(n8346), .ZN(n9637) );
  AOI22_X1 U4664 ( .A1(ram[3717]), .A2(n8341), .B1(n9648), .B2(n8975), .ZN(
        n8346) );
  INV_X1 U4665 ( .A(n8347), .ZN(n9638) );
  AOI22_X1 U4666 ( .A1(ram[3718]), .A2(n8341), .B1(n9648), .B2(n8999), .ZN(
        n8347) );
  INV_X1 U4667 ( .A(n8348), .ZN(n9639) );
  AOI22_X1 U4668 ( .A1(ram[3719]), .A2(n8341), .B1(n9648), .B2(n9023), .ZN(
        n8348) );
  INV_X1 U4669 ( .A(n8349), .ZN(n9640) );
  AOI22_X1 U4670 ( .A1(ram[3720]), .A2(n8341), .B1(n9648), .B2(n9047), .ZN(
        n8349) );
  INV_X1 U4671 ( .A(n8350), .ZN(n9641) );
  AOI22_X1 U4672 ( .A1(ram[3721]), .A2(n8341), .B1(n9648), .B2(n9071), .ZN(
        n8350) );
  INV_X1 U4673 ( .A(n8351), .ZN(n9642) );
  AOI22_X1 U4674 ( .A1(ram[3722]), .A2(n8341), .B1(n9648), .B2(n9095), .ZN(
        n8351) );
  INV_X1 U4675 ( .A(n8352), .ZN(n9643) );
  AOI22_X1 U4676 ( .A1(ram[3723]), .A2(n8341), .B1(n9648), .B2(n9119), .ZN(
        n8352) );
  INV_X1 U4677 ( .A(n8353), .ZN(n9644) );
  AOI22_X1 U4678 ( .A1(ram[3724]), .A2(n8341), .B1(n9648), .B2(n9143), .ZN(
        n8353) );
  INV_X1 U4679 ( .A(n8354), .ZN(n9645) );
  AOI22_X1 U4680 ( .A1(ram[3725]), .A2(n8341), .B1(n9648), .B2(n9167), .ZN(
        n8354) );
  INV_X1 U4681 ( .A(n8355), .ZN(n9646) );
  AOI22_X1 U4682 ( .A1(ram[3726]), .A2(n8341), .B1(n9648), .B2(n9191), .ZN(
        n8355) );
  INV_X1 U4683 ( .A(n8356), .ZN(n9647) );
  AOI22_X1 U4684 ( .A1(ram[3727]), .A2(n8341), .B1(n9648), .B2(n9215), .ZN(
        n8356) );
  INV_X1 U4685 ( .A(n8374), .ZN(n9598) );
  AOI22_X1 U4686 ( .A1(ram[3744]), .A2(n8375), .B1(n9614), .B2(n8855), .ZN(
        n8374) );
  INV_X1 U4687 ( .A(n8376), .ZN(n9599) );
  AOI22_X1 U4688 ( .A1(ram[3745]), .A2(n8375), .B1(n9614), .B2(n8879), .ZN(
        n8376) );
  INV_X1 U4689 ( .A(n8377), .ZN(n9600) );
  AOI22_X1 U4690 ( .A1(ram[3746]), .A2(n8375), .B1(n9614), .B2(n8903), .ZN(
        n8377) );
  INV_X1 U4691 ( .A(n8378), .ZN(n9601) );
  AOI22_X1 U4692 ( .A1(ram[3747]), .A2(n8375), .B1(n9614), .B2(n8927), .ZN(
        n8378) );
  INV_X1 U4693 ( .A(n8379), .ZN(n9602) );
  AOI22_X1 U4694 ( .A1(ram[3748]), .A2(n8375), .B1(n9614), .B2(n8951), .ZN(
        n8379) );
  INV_X1 U4695 ( .A(n8380), .ZN(n9603) );
  AOI22_X1 U4696 ( .A1(ram[3749]), .A2(n8375), .B1(n9614), .B2(n8975), .ZN(
        n8380) );
  INV_X1 U4697 ( .A(n8381), .ZN(n9604) );
  AOI22_X1 U4698 ( .A1(ram[3750]), .A2(n8375), .B1(n9614), .B2(n8999), .ZN(
        n8381) );
  INV_X1 U4699 ( .A(n8382), .ZN(n9605) );
  AOI22_X1 U4700 ( .A1(ram[3751]), .A2(n8375), .B1(n9614), .B2(n9023), .ZN(
        n8382) );
  INV_X1 U4701 ( .A(n8383), .ZN(n9606) );
  AOI22_X1 U4702 ( .A1(ram[3752]), .A2(n8375), .B1(n9614), .B2(n9047), .ZN(
        n8383) );
  INV_X1 U4703 ( .A(n8384), .ZN(n9607) );
  AOI22_X1 U4704 ( .A1(ram[3753]), .A2(n8375), .B1(n9614), .B2(n9071), .ZN(
        n8384) );
  INV_X1 U4705 ( .A(n8385), .ZN(n9608) );
  AOI22_X1 U4706 ( .A1(ram[3754]), .A2(n8375), .B1(n9614), .B2(n9095), .ZN(
        n8385) );
  INV_X1 U4707 ( .A(n8386), .ZN(n9609) );
  AOI22_X1 U4708 ( .A1(ram[3755]), .A2(n8375), .B1(n9614), .B2(n9119), .ZN(
        n8386) );
  INV_X1 U4709 ( .A(n8387), .ZN(n9610) );
  AOI22_X1 U4710 ( .A1(ram[3756]), .A2(n8375), .B1(n9614), .B2(n9143), .ZN(
        n8387) );
  INV_X1 U4711 ( .A(n8388), .ZN(n9611) );
  AOI22_X1 U4712 ( .A1(ram[3757]), .A2(n8375), .B1(n9614), .B2(n9167), .ZN(
        n8388) );
  INV_X1 U4713 ( .A(n8389), .ZN(n9612) );
  AOI22_X1 U4714 ( .A1(ram[3758]), .A2(n8375), .B1(n9614), .B2(n9191), .ZN(
        n8389) );
  INV_X1 U4715 ( .A(n8390), .ZN(n9613) );
  AOI22_X1 U4716 ( .A1(ram[3759]), .A2(n8375), .B1(n9614), .B2(n9215), .ZN(
        n8390) );
  INV_X1 U4717 ( .A(n8408), .ZN(n9564) );
  AOI22_X1 U4718 ( .A1(ram[3776]), .A2(n8409), .B1(n9580), .B2(n8855), .ZN(
        n8408) );
  INV_X1 U4719 ( .A(n8410), .ZN(n9565) );
  AOI22_X1 U4720 ( .A1(ram[3777]), .A2(n8409), .B1(n9580), .B2(n8879), .ZN(
        n8410) );
  INV_X1 U4721 ( .A(n8411), .ZN(n9566) );
  AOI22_X1 U4722 ( .A1(ram[3778]), .A2(n8409), .B1(n9580), .B2(n8903), .ZN(
        n8411) );
  INV_X1 U4723 ( .A(n8412), .ZN(n9567) );
  AOI22_X1 U4724 ( .A1(ram[3779]), .A2(n8409), .B1(n9580), .B2(n8927), .ZN(
        n8412) );
  INV_X1 U4725 ( .A(n8413), .ZN(n9568) );
  AOI22_X1 U4726 ( .A1(ram[3780]), .A2(n8409), .B1(n9580), .B2(n8951), .ZN(
        n8413) );
  INV_X1 U4727 ( .A(n8414), .ZN(n9569) );
  AOI22_X1 U4728 ( .A1(ram[3781]), .A2(n8409), .B1(n9580), .B2(n8975), .ZN(
        n8414) );
  INV_X1 U4729 ( .A(n8415), .ZN(n9570) );
  AOI22_X1 U4730 ( .A1(ram[3782]), .A2(n8409), .B1(n9580), .B2(n8999), .ZN(
        n8415) );
  INV_X1 U4731 ( .A(n8416), .ZN(n9571) );
  AOI22_X1 U4732 ( .A1(ram[3783]), .A2(n8409), .B1(n9580), .B2(n9023), .ZN(
        n8416) );
  INV_X1 U4733 ( .A(n8417), .ZN(n9572) );
  AOI22_X1 U4734 ( .A1(ram[3784]), .A2(n8409), .B1(n9580), .B2(n9047), .ZN(
        n8417) );
  INV_X1 U4735 ( .A(n8418), .ZN(n9573) );
  AOI22_X1 U4736 ( .A1(ram[3785]), .A2(n8409), .B1(n9580), .B2(n9071), .ZN(
        n8418) );
  INV_X1 U4737 ( .A(n8419), .ZN(n9574) );
  AOI22_X1 U4738 ( .A1(ram[3786]), .A2(n8409), .B1(n9580), .B2(n9095), .ZN(
        n8419) );
  INV_X1 U4739 ( .A(n8420), .ZN(n9575) );
  AOI22_X1 U4740 ( .A1(ram[3787]), .A2(n8409), .B1(n9580), .B2(n9119), .ZN(
        n8420) );
  INV_X1 U4741 ( .A(n8421), .ZN(n9576) );
  AOI22_X1 U4742 ( .A1(ram[3788]), .A2(n8409), .B1(n9580), .B2(n9143), .ZN(
        n8421) );
  INV_X1 U4743 ( .A(n8422), .ZN(n9577) );
  AOI22_X1 U4744 ( .A1(ram[3789]), .A2(n8409), .B1(n9580), .B2(n9167), .ZN(
        n8422) );
  INV_X1 U4745 ( .A(n8423), .ZN(n9578) );
  AOI22_X1 U4746 ( .A1(ram[3790]), .A2(n8409), .B1(n9580), .B2(n9191), .ZN(
        n8423) );
  INV_X1 U4747 ( .A(n8424), .ZN(n9579) );
  AOI22_X1 U4748 ( .A1(ram[3791]), .A2(n8409), .B1(n9580), .B2(n9215), .ZN(
        n8424) );
  INV_X1 U4749 ( .A(n8442), .ZN(n9530) );
  AOI22_X1 U4750 ( .A1(ram[3808]), .A2(n8443), .B1(n9546), .B2(n8855), .ZN(
        n8442) );
  INV_X1 U4751 ( .A(n8444), .ZN(n9531) );
  AOI22_X1 U4752 ( .A1(ram[3809]), .A2(n8443), .B1(n9546), .B2(n8879), .ZN(
        n8444) );
  INV_X1 U4753 ( .A(n8445), .ZN(n9532) );
  AOI22_X1 U4754 ( .A1(ram[3810]), .A2(n8443), .B1(n9546), .B2(n8903), .ZN(
        n8445) );
  INV_X1 U4755 ( .A(n8446), .ZN(n9533) );
  AOI22_X1 U4756 ( .A1(ram[3811]), .A2(n8443), .B1(n9546), .B2(n8927), .ZN(
        n8446) );
  INV_X1 U4757 ( .A(n8447), .ZN(n9534) );
  AOI22_X1 U4758 ( .A1(ram[3812]), .A2(n8443), .B1(n9546), .B2(n8951), .ZN(
        n8447) );
  INV_X1 U4759 ( .A(n8448), .ZN(n9535) );
  AOI22_X1 U4760 ( .A1(ram[3813]), .A2(n8443), .B1(n9546), .B2(n8975), .ZN(
        n8448) );
  INV_X1 U4761 ( .A(n8449), .ZN(n9536) );
  AOI22_X1 U4762 ( .A1(ram[3814]), .A2(n8443), .B1(n9546), .B2(n8999), .ZN(
        n8449) );
  INV_X1 U4763 ( .A(n8450), .ZN(n9537) );
  AOI22_X1 U4764 ( .A1(ram[3815]), .A2(n8443), .B1(n9546), .B2(n9023), .ZN(
        n8450) );
  INV_X1 U4765 ( .A(n8451), .ZN(n9538) );
  AOI22_X1 U4766 ( .A1(ram[3816]), .A2(n8443), .B1(n9546), .B2(n9047), .ZN(
        n8451) );
  INV_X1 U4767 ( .A(n8452), .ZN(n9539) );
  AOI22_X1 U4768 ( .A1(ram[3817]), .A2(n8443), .B1(n9546), .B2(n9071), .ZN(
        n8452) );
  INV_X1 U4769 ( .A(n8453), .ZN(n9540) );
  AOI22_X1 U4770 ( .A1(ram[3818]), .A2(n8443), .B1(n9546), .B2(n9095), .ZN(
        n8453) );
  INV_X1 U4771 ( .A(n8454), .ZN(n9541) );
  AOI22_X1 U4772 ( .A1(ram[3819]), .A2(n8443), .B1(n9546), .B2(n9119), .ZN(
        n8454) );
  INV_X1 U4773 ( .A(n8455), .ZN(n9542) );
  AOI22_X1 U4774 ( .A1(ram[3820]), .A2(n8443), .B1(n9546), .B2(n9143), .ZN(
        n8455) );
  INV_X1 U4775 ( .A(n8456), .ZN(n9543) );
  AOI22_X1 U4776 ( .A1(ram[3821]), .A2(n8443), .B1(n9546), .B2(n9167), .ZN(
        n8456) );
  INV_X1 U4777 ( .A(n8457), .ZN(n9544) );
  AOI22_X1 U4778 ( .A1(ram[3822]), .A2(n8443), .B1(n9546), .B2(n9191), .ZN(
        n8457) );
  INV_X1 U4779 ( .A(n8458), .ZN(n9545) );
  AOI22_X1 U4780 ( .A1(ram[3823]), .A2(n8443), .B1(n9546), .B2(n9215), .ZN(
        n8458) );
  INV_X1 U4781 ( .A(n8476), .ZN(n9496) );
  AOI22_X1 U4782 ( .A1(ram[3840]), .A2(n8477), .B1(n9512), .B2(n8855), .ZN(
        n8476) );
  INV_X1 U4783 ( .A(n8478), .ZN(n9497) );
  AOI22_X1 U4784 ( .A1(ram[3841]), .A2(n8477), .B1(n9512), .B2(n8879), .ZN(
        n8478) );
  INV_X1 U4785 ( .A(n8479), .ZN(n9498) );
  AOI22_X1 U4786 ( .A1(ram[3842]), .A2(n8477), .B1(n9512), .B2(n8903), .ZN(
        n8479) );
  INV_X1 U4787 ( .A(n8480), .ZN(n9499) );
  AOI22_X1 U4788 ( .A1(ram[3843]), .A2(n8477), .B1(n9512), .B2(n8927), .ZN(
        n8480) );
  INV_X1 U4789 ( .A(n8481), .ZN(n9500) );
  AOI22_X1 U4790 ( .A1(ram[3844]), .A2(n8477), .B1(n9512), .B2(n8951), .ZN(
        n8481) );
  INV_X1 U4791 ( .A(n8482), .ZN(n9501) );
  AOI22_X1 U4792 ( .A1(ram[3845]), .A2(n8477), .B1(n9512), .B2(n8975), .ZN(
        n8482) );
  INV_X1 U4793 ( .A(n8483), .ZN(n9502) );
  AOI22_X1 U4794 ( .A1(ram[3846]), .A2(n8477), .B1(n9512), .B2(n8999), .ZN(
        n8483) );
  INV_X1 U4795 ( .A(n8484), .ZN(n9503) );
  AOI22_X1 U4796 ( .A1(ram[3847]), .A2(n8477), .B1(n9512), .B2(n9023), .ZN(
        n8484) );
  INV_X1 U4797 ( .A(n8485), .ZN(n9504) );
  AOI22_X1 U4798 ( .A1(ram[3848]), .A2(n8477), .B1(n9512), .B2(n9047), .ZN(
        n8485) );
  INV_X1 U4799 ( .A(n8486), .ZN(n9505) );
  AOI22_X1 U4800 ( .A1(ram[3849]), .A2(n8477), .B1(n9512), .B2(n9071), .ZN(
        n8486) );
  INV_X1 U4801 ( .A(n8487), .ZN(n9506) );
  AOI22_X1 U4802 ( .A1(ram[3850]), .A2(n8477), .B1(n9512), .B2(n9095), .ZN(
        n8487) );
  INV_X1 U4803 ( .A(n8488), .ZN(n9507) );
  AOI22_X1 U4804 ( .A1(ram[3851]), .A2(n8477), .B1(n9512), .B2(n9119), .ZN(
        n8488) );
  INV_X1 U4805 ( .A(n8489), .ZN(n9508) );
  AOI22_X1 U4806 ( .A1(ram[3852]), .A2(n8477), .B1(n9512), .B2(n9143), .ZN(
        n8489) );
  INV_X1 U4807 ( .A(n8490), .ZN(n9509) );
  AOI22_X1 U4808 ( .A1(ram[3853]), .A2(n8477), .B1(n9512), .B2(n9167), .ZN(
        n8490) );
  INV_X1 U4809 ( .A(n8491), .ZN(n9510) );
  AOI22_X1 U4810 ( .A1(ram[3854]), .A2(n8477), .B1(n9512), .B2(n9191), .ZN(
        n8491) );
  INV_X1 U4811 ( .A(n8492), .ZN(n9511) );
  AOI22_X1 U4812 ( .A1(ram[3855]), .A2(n8477), .B1(n9512), .B2(n9215), .ZN(
        n8492) );
  INV_X1 U4813 ( .A(n8514), .ZN(n9462) );
  AOI22_X1 U4814 ( .A1(ram[3872]), .A2(n8515), .B1(n9478), .B2(n8855), .ZN(
        n8514) );
  INV_X1 U4815 ( .A(n8516), .ZN(n9463) );
  AOI22_X1 U4816 ( .A1(ram[3873]), .A2(n8515), .B1(n9478), .B2(n8879), .ZN(
        n8516) );
  INV_X1 U4817 ( .A(n8517), .ZN(n9464) );
  AOI22_X1 U4818 ( .A1(ram[3874]), .A2(n8515), .B1(n9478), .B2(n8903), .ZN(
        n8517) );
  INV_X1 U4819 ( .A(n8518), .ZN(n9465) );
  AOI22_X1 U4820 ( .A1(ram[3875]), .A2(n8515), .B1(n9478), .B2(n8927), .ZN(
        n8518) );
  INV_X1 U4821 ( .A(n8519), .ZN(n9466) );
  AOI22_X1 U4822 ( .A1(ram[3876]), .A2(n8515), .B1(n9478), .B2(n8951), .ZN(
        n8519) );
  INV_X1 U4823 ( .A(n8520), .ZN(n9467) );
  AOI22_X1 U4824 ( .A1(ram[3877]), .A2(n8515), .B1(n9478), .B2(n8975), .ZN(
        n8520) );
  INV_X1 U4825 ( .A(n8521), .ZN(n9468) );
  AOI22_X1 U4826 ( .A1(ram[3878]), .A2(n8515), .B1(n9478), .B2(n8999), .ZN(
        n8521) );
  INV_X1 U4827 ( .A(n8522), .ZN(n9469) );
  AOI22_X1 U4828 ( .A1(ram[3879]), .A2(n8515), .B1(n9478), .B2(n9023), .ZN(
        n8522) );
  INV_X1 U4829 ( .A(n8523), .ZN(n9470) );
  AOI22_X1 U4830 ( .A1(ram[3880]), .A2(n8515), .B1(n9478), .B2(n9047), .ZN(
        n8523) );
  INV_X1 U4831 ( .A(n8524), .ZN(n9471) );
  AOI22_X1 U4832 ( .A1(ram[3881]), .A2(n8515), .B1(n9478), .B2(n9071), .ZN(
        n8524) );
  INV_X1 U4833 ( .A(n8525), .ZN(n9472) );
  AOI22_X1 U4834 ( .A1(ram[3882]), .A2(n8515), .B1(n9478), .B2(n9095), .ZN(
        n8525) );
  INV_X1 U4835 ( .A(n8526), .ZN(n9473) );
  AOI22_X1 U4836 ( .A1(ram[3883]), .A2(n8515), .B1(n9478), .B2(n9119), .ZN(
        n8526) );
  INV_X1 U4837 ( .A(n8527), .ZN(n9474) );
  AOI22_X1 U4838 ( .A1(ram[3884]), .A2(n8515), .B1(n9478), .B2(n9143), .ZN(
        n8527) );
  INV_X1 U4839 ( .A(n8528), .ZN(n9475) );
  AOI22_X1 U4840 ( .A1(ram[3885]), .A2(n8515), .B1(n9478), .B2(n9167), .ZN(
        n8528) );
  INV_X1 U4841 ( .A(n8529), .ZN(n9476) );
  AOI22_X1 U4842 ( .A1(ram[3886]), .A2(n8515), .B1(n9478), .B2(n9191), .ZN(
        n8529) );
  INV_X1 U4843 ( .A(n8530), .ZN(n9477) );
  AOI22_X1 U4844 ( .A1(ram[3887]), .A2(n8515), .B1(n9478), .B2(n9215), .ZN(
        n8530) );
  INV_X1 U4845 ( .A(n8550), .ZN(n9428) );
  AOI22_X1 U4846 ( .A1(ram[3904]), .A2(n8551), .B1(n9444), .B2(n8854), .ZN(
        n8550) );
  INV_X1 U4847 ( .A(n8552), .ZN(n9429) );
  AOI22_X1 U4848 ( .A1(ram[3905]), .A2(n8551), .B1(n9444), .B2(n8878), .ZN(
        n8552) );
  INV_X1 U4849 ( .A(n8553), .ZN(n9430) );
  AOI22_X1 U4850 ( .A1(ram[3906]), .A2(n8551), .B1(n9444), .B2(n8902), .ZN(
        n8553) );
  INV_X1 U4851 ( .A(n8554), .ZN(n9431) );
  AOI22_X1 U4852 ( .A1(ram[3907]), .A2(n8551), .B1(n9444), .B2(n8926), .ZN(
        n8554) );
  INV_X1 U4853 ( .A(n8555), .ZN(n9432) );
  AOI22_X1 U4854 ( .A1(ram[3908]), .A2(n8551), .B1(n9444), .B2(n8950), .ZN(
        n8555) );
  INV_X1 U4855 ( .A(n8556), .ZN(n9433) );
  AOI22_X1 U4856 ( .A1(ram[3909]), .A2(n8551), .B1(n9444), .B2(n8974), .ZN(
        n8556) );
  INV_X1 U4857 ( .A(n8557), .ZN(n9434) );
  AOI22_X1 U4858 ( .A1(ram[3910]), .A2(n8551), .B1(n9444), .B2(n8998), .ZN(
        n8557) );
  INV_X1 U4859 ( .A(n8558), .ZN(n9435) );
  AOI22_X1 U4860 ( .A1(ram[3911]), .A2(n8551), .B1(n9444), .B2(n9022), .ZN(
        n8558) );
  INV_X1 U4861 ( .A(n8559), .ZN(n9436) );
  AOI22_X1 U4862 ( .A1(ram[3912]), .A2(n8551), .B1(n9444), .B2(n9046), .ZN(
        n8559) );
  INV_X1 U4863 ( .A(n8560), .ZN(n9437) );
  AOI22_X1 U4864 ( .A1(ram[3913]), .A2(n8551), .B1(n9444), .B2(n9070), .ZN(
        n8560) );
  INV_X1 U4865 ( .A(n8561), .ZN(n9438) );
  AOI22_X1 U4866 ( .A1(ram[3914]), .A2(n8551), .B1(n9444), .B2(n9094), .ZN(
        n8561) );
  INV_X1 U4867 ( .A(n8562), .ZN(n9439) );
  AOI22_X1 U4868 ( .A1(ram[3915]), .A2(n8551), .B1(n9444), .B2(n9118), .ZN(
        n8562) );
  INV_X1 U4869 ( .A(n8563), .ZN(n9440) );
  AOI22_X1 U4870 ( .A1(ram[3916]), .A2(n8551), .B1(n9444), .B2(n9142), .ZN(
        n8563) );
  INV_X1 U4871 ( .A(n8564), .ZN(n9441) );
  AOI22_X1 U4872 ( .A1(ram[3917]), .A2(n8551), .B1(n9444), .B2(n9166), .ZN(
        n8564) );
  INV_X1 U4873 ( .A(n8565), .ZN(n9442) );
  AOI22_X1 U4874 ( .A1(ram[3918]), .A2(n8551), .B1(n9444), .B2(n9190), .ZN(
        n8565) );
  INV_X1 U4875 ( .A(n8566), .ZN(n9443) );
  AOI22_X1 U4876 ( .A1(ram[3919]), .A2(n8551), .B1(n9444), .B2(n9214), .ZN(
        n8566) );
  INV_X1 U4877 ( .A(n8585), .ZN(n9394) );
  AOI22_X1 U4878 ( .A1(ram[3936]), .A2(n8586), .B1(n9410), .B2(n8854), .ZN(
        n8585) );
  INV_X1 U4879 ( .A(n8587), .ZN(n9395) );
  AOI22_X1 U4880 ( .A1(ram[3937]), .A2(n8586), .B1(n9410), .B2(n8878), .ZN(
        n8587) );
  INV_X1 U4881 ( .A(n8588), .ZN(n9396) );
  AOI22_X1 U4882 ( .A1(ram[3938]), .A2(n8586), .B1(n9410), .B2(n8902), .ZN(
        n8588) );
  INV_X1 U4883 ( .A(n8589), .ZN(n9397) );
  AOI22_X1 U4884 ( .A1(ram[3939]), .A2(n8586), .B1(n9410), .B2(n8926), .ZN(
        n8589) );
  INV_X1 U4885 ( .A(n8590), .ZN(n9398) );
  AOI22_X1 U4886 ( .A1(ram[3940]), .A2(n8586), .B1(n9410), .B2(n8950), .ZN(
        n8590) );
  INV_X1 U4887 ( .A(n8591), .ZN(n9399) );
  AOI22_X1 U4888 ( .A1(ram[3941]), .A2(n8586), .B1(n9410), .B2(n8974), .ZN(
        n8591) );
  INV_X1 U4889 ( .A(n8592), .ZN(n9400) );
  AOI22_X1 U4890 ( .A1(ram[3942]), .A2(n8586), .B1(n9410), .B2(n8998), .ZN(
        n8592) );
  INV_X1 U4891 ( .A(n8593), .ZN(n9401) );
  AOI22_X1 U4892 ( .A1(ram[3943]), .A2(n8586), .B1(n9410), .B2(n9022), .ZN(
        n8593) );
  INV_X1 U4893 ( .A(n8594), .ZN(n9402) );
  AOI22_X1 U4894 ( .A1(ram[3944]), .A2(n8586), .B1(n9410), .B2(n9046), .ZN(
        n8594) );
  INV_X1 U4895 ( .A(n8595), .ZN(n9403) );
  AOI22_X1 U4896 ( .A1(ram[3945]), .A2(n8586), .B1(n9410), .B2(n9070), .ZN(
        n8595) );
  INV_X1 U4897 ( .A(n8596), .ZN(n9404) );
  AOI22_X1 U4898 ( .A1(ram[3946]), .A2(n8586), .B1(n9410), .B2(n9094), .ZN(
        n8596) );
  INV_X1 U4899 ( .A(n8597), .ZN(n9405) );
  AOI22_X1 U4900 ( .A1(ram[3947]), .A2(n8586), .B1(n9410), .B2(n9118), .ZN(
        n8597) );
  INV_X1 U4901 ( .A(n8598), .ZN(n9406) );
  AOI22_X1 U4902 ( .A1(ram[3948]), .A2(n8586), .B1(n9410), .B2(n9142), .ZN(
        n8598) );
  INV_X1 U4903 ( .A(n8599), .ZN(n9407) );
  AOI22_X1 U4904 ( .A1(ram[3949]), .A2(n8586), .B1(n9410), .B2(n9166), .ZN(
        n8599) );
  INV_X1 U4905 ( .A(n8600), .ZN(n9408) );
  AOI22_X1 U4906 ( .A1(ram[3950]), .A2(n8586), .B1(n9410), .B2(n9190), .ZN(
        n8600) );
  INV_X1 U4907 ( .A(n8601), .ZN(n9409) );
  AOI22_X1 U4908 ( .A1(ram[3951]), .A2(n8586), .B1(n9410), .B2(n9214), .ZN(
        n8601) );
  INV_X1 U4909 ( .A(n8619), .ZN(n9360) );
  AOI22_X1 U4910 ( .A1(ram[3968]), .A2(n8620), .B1(n9376), .B2(n8854), .ZN(
        n8619) );
  INV_X1 U4911 ( .A(n8621), .ZN(n9361) );
  AOI22_X1 U4912 ( .A1(ram[3969]), .A2(n8620), .B1(n9376), .B2(n8878), .ZN(
        n8621) );
  INV_X1 U4913 ( .A(n8622), .ZN(n9362) );
  AOI22_X1 U4914 ( .A1(ram[3970]), .A2(n8620), .B1(n9376), .B2(n8902), .ZN(
        n8622) );
  INV_X1 U4915 ( .A(n8623), .ZN(n9363) );
  AOI22_X1 U4916 ( .A1(ram[3971]), .A2(n8620), .B1(n9376), .B2(n8926), .ZN(
        n8623) );
  INV_X1 U4917 ( .A(n8624), .ZN(n9364) );
  AOI22_X1 U4918 ( .A1(ram[3972]), .A2(n8620), .B1(n9376), .B2(n8950), .ZN(
        n8624) );
  INV_X1 U4919 ( .A(n8625), .ZN(n9365) );
  AOI22_X1 U4920 ( .A1(ram[3973]), .A2(n8620), .B1(n9376), .B2(n8974), .ZN(
        n8625) );
  INV_X1 U4921 ( .A(n8626), .ZN(n9366) );
  AOI22_X1 U4922 ( .A1(ram[3974]), .A2(n8620), .B1(n9376), .B2(n8998), .ZN(
        n8626) );
  INV_X1 U4923 ( .A(n8627), .ZN(n9367) );
  AOI22_X1 U4924 ( .A1(ram[3975]), .A2(n8620), .B1(n9376), .B2(n9022), .ZN(
        n8627) );
  INV_X1 U4925 ( .A(n8628), .ZN(n9368) );
  AOI22_X1 U4926 ( .A1(ram[3976]), .A2(n8620), .B1(n9376), .B2(n9046), .ZN(
        n8628) );
  INV_X1 U4927 ( .A(n8629), .ZN(n9369) );
  AOI22_X1 U4928 ( .A1(ram[3977]), .A2(n8620), .B1(n9376), .B2(n9070), .ZN(
        n8629) );
  INV_X1 U4929 ( .A(n8630), .ZN(n9370) );
  AOI22_X1 U4930 ( .A1(ram[3978]), .A2(n8620), .B1(n9376), .B2(n9094), .ZN(
        n8630) );
  INV_X1 U4931 ( .A(n8631), .ZN(n9371) );
  AOI22_X1 U4932 ( .A1(ram[3979]), .A2(n8620), .B1(n9376), .B2(n9118), .ZN(
        n8631) );
  INV_X1 U4933 ( .A(n8632), .ZN(n9372) );
  AOI22_X1 U4934 ( .A1(ram[3980]), .A2(n8620), .B1(n9376), .B2(n9142), .ZN(
        n8632) );
  INV_X1 U4935 ( .A(n8633), .ZN(n9373) );
  AOI22_X1 U4936 ( .A1(ram[3981]), .A2(n8620), .B1(n9376), .B2(n9166), .ZN(
        n8633) );
  INV_X1 U4937 ( .A(n8634), .ZN(n9374) );
  AOI22_X1 U4938 ( .A1(ram[3982]), .A2(n8620), .B1(n9376), .B2(n9190), .ZN(
        n8634) );
  INV_X1 U4939 ( .A(n8635), .ZN(n9375) );
  AOI22_X1 U4940 ( .A1(ram[3983]), .A2(n8620), .B1(n9376), .B2(n9214), .ZN(
        n8635) );
  INV_X1 U4941 ( .A(n8654), .ZN(n9326) );
  AOI22_X1 U4942 ( .A1(ram[4000]), .A2(n8655), .B1(n9342), .B2(n8854), .ZN(
        n8654) );
  INV_X1 U4943 ( .A(n8656), .ZN(n9327) );
  AOI22_X1 U4944 ( .A1(ram[4001]), .A2(n8655), .B1(n9342), .B2(n8878), .ZN(
        n8656) );
  INV_X1 U4945 ( .A(n8657), .ZN(n9328) );
  AOI22_X1 U4946 ( .A1(ram[4002]), .A2(n8655), .B1(n9342), .B2(n8902), .ZN(
        n8657) );
  INV_X1 U4947 ( .A(n8658), .ZN(n9329) );
  AOI22_X1 U4948 ( .A1(ram[4003]), .A2(n8655), .B1(n9342), .B2(n8926), .ZN(
        n8658) );
  INV_X1 U4949 ( .A(n8659), .ZN(n9330) );
  AOI22_X1 U4950 ( .A1(ram[4004]), .A2(n8655), .B1(n9342), .B2(n8950), .ZN(
        n8659) );
  INV_X1 U4951 ( .A(n8660), .ZN(n9331) );
  AOI22_X1 U4952 ( .A1(ram[4005]), .A2(n8655), .B1(n9342), .B2(n8974), .ZN(
        n8660) );
  INV_X1 U4953 ( .A(n8661), .ZN(n9332) );
  AOI22_X1 U4954 ( .A1(ram[4006]), .A2(n8655), .B1(n9342), .B2(n8998), .ZN(
        n8661) );
  INV_X1 U4955 ( .A(n8662), .ZN(n9333) );
  AOI22_X1 U4956 ( .A1(ram[4007]), .A2(n8655), .B1(n9342), .B2(n9022), .ZN(
        n8662) );
  INV_X1 U4957 ( .A(n8663), .ZN(n9334) );
  AOI22_X1 U4958 ( .A1(ram[4008]), .A2(n8655), .B1(n9342), .B2(n9046), .ZN(
        n8663) );
  INV_X1 U4959 ( .A(n8664), .ZN(n9335) );
  AOI22_X1 U4960 ( .A1(ram[4009]), .A2(n8655), .B1(n9342), .B2(n9070), .ZN(
        n8664) );
  INV_X1 U4961 ( .A(n8665), .ZN(n9336) );
  AOI22_X1 U4962 ( .A1(ram[4010]), .A2(n8655), .B1(n9342), .B2(n9094), .ZN(
        n8665) );
  INV_X1 U4963 ( .A(n8666), .ZN(n9337) );
  AOI22_X1 U4964 ( .A1(ram[4011]), .A2(n8655), .B1(n9342), .B2(n9118), .ZN(
        n8666) );
  INV_X1 U4965 ( .A(n8667), .ZN(n9338) );
  AOI22_X1 U4966 ( .A1(ram[4012]), .A2(n8655), .B1(n9342), .B2(n9142), .ZN(
        n8667) );
  INV_X1 U4967 ( .A(n8668), .ZN(n9339) );
  AOI22_X1 U4968 ( .A1(ram[4013]), .A2(n8655), .B1(n9342), .B2(n9166), .ZN(
        n8668) );
  INV_X1 U4969 ( .A(n8669), .ZN(n9340) );
  AOI22_X1 U4970 ( .A1(ram[4014]), .A2(n8655), .B1(n9342), .B2(n9190), .ZN(
        n8669) );
  INV_X1 U4971 ( .A(n8670), .ZN(n9341) );
  AOI22_X1 U4972 ( .A1(ram[4015]), .A2(n8655), .B1(n9342), .B2(n9214), .ZN(
        n8670) );
  INV_X1 U4973 ( .A(n8688), .ZN(n9292) );
  AOI22_X1 U4974 ( .A1(ram[4032]), .A2(n8689), .B1(n9308), .B2(n8854), .ZN(
        n8688) );
  INV_X1 U4975 ( .A(n8690), .ZN(n9293) );
  AOI22_X1 U4976 ( .A1(ram[4033]), .A2(n8689), .B1(n9308), .B2(n8878), .ZN(
        n8690) );
  INV_X1 U4977 ( .A(n8691), .ZN(n9294) );
  AOI22_X1 U4978 ( .A1(ram[4034]), .A2(n8689), .B1(n9308), .B2(n8902), .ZN(
        n8691) );
  INV_X1 U4979 ( .A(n8692), .ZN(n9295) );
  AOI22_X1 U4980 ( .A1(ram[4035]), .A2(n8689), .B1(n9308), .B2(n8926), .ZN(
        n8692) );
  INV_X1 U4981 ( .A(n8693), .ZN(n9296) );
  AOI22_X1 U4982 ( .A1(ram[4036]), .A2(n8689), .B1(n9308), .B2(n8950), .ZN(
        n8693) );
  INV_X1 U4983 ( .A(n8694), .ZN(n9297) );
  AOI22_X1 U4984 ( .A1(ram[4037]), .A2(n8689), .B1(n9308), .B2(n8974), .ZN(
        n8694) );
  INV_X1 U4985 ( .A(n8695), .ZN(n9298) );
  AOI22_X1 U4986 ( .A1(ram[4038]), .A2(n8689), .B1(n9308), .B2(n8998), .ZN(
        n8695) );
  INV_X1 U4987 ( .A(n8696), .ZN(n9299) );
  AOI22_X1 U4988 ( .A1(ram[4039]), .A2(n8689), .B1(n9308), .B2(n9022), .ZN(
        n8696) );
  INV_X1 U4989 ( .A(n8697), .ZN(n9300) );
  AOI22_X1 U4990 ( .A1(ram[4040]), .A2(n8689), .B1(n9308), .B2(n9046), .ZN(
        n8697) );
  INV_X1 U4991 ( .A(n8698), .ZN(n9301) );
  AOI22_X1 U4992 ( .A1(ram[4041]), .A2(n8689), .B1(n9308), .B2(n9070), .ZN(
        n8698) );
  INV_X1 U4993 ( .A(n8699), .ZN(n9302) );
  AOI22_X1 U4994 ( .A1(ram[4042]), .A2(n8689), .B1(n9308), .B2(n9094), .ZN(
        n8699) );
  INV_X1 U4995 ( .A(n8700), .ZN(n9303) );
  AOI22_X1 U4996 ( .A1(ram[4043]), .A2(n8689), .B1(n9308), .B2(n9118), .ZN(
        n8700) );
  INV_X1 U4997 ( .A(n8701), .ZN(n9304) );
  AOI22_X1 U4998 ( .A1(ram[4044]), .A2(n8689), .B1(n9308), .B2(n9142), .ZN(
        n8701) );
  INV_X1 U4999 ( .A(n8702), .ZN(n9305) );
  AOI22_X1 U5000 ( .A1(ram[4045]), .A2(n8689), .B1(n9308), .B2(n9166), .ZN(
        n8702) );
  INV_X1 U5001 ( .A(n8703), .ZN(n9306) );
  AOI22_X1 U5002 ( .A1(ram[4046]), .A2(n8689), .B1(n9308), .B2(n9190), .ZN(
        n8703) );
  INV_X1 U5003 ( .A(n8704), .ZN(n9307) );
  AOI22_X1 U5004 ( .A1(ram[4047]), .A2(n8689), .B1(n9308), .B2(n9214), .ZN(
        n8704) );
  INV_X1 U5005 ( .A(n8723), .ZN(n9258) );
  AOI22_X1 U5006 ( .A1(ram[4064]), .A2(n8724), .B1(n9274), .B2(n8854), .ZN(
        n8723) );
  INV_X1 U5007 ( .A(n8725), .ZN(n9259) );
  AOI22_X1 U5008 ( .A1(ram[4065]), .A2(n8724), .B1(n9274), .B2(n8878), .ZN(
        n8725) );
  INV_X1 U5009 ( .A(n8726), .ZN(n9260) );
  AOI22_X1 U5010 ( .A1(ram[4066]), .A2(n8724), .B1(n9274), .B2(n8902), .ZN(
        n8726) );
  INV_X1 U5011 ( .A(n8727), .ZN(n9261) );
  AOI22_X1 U5012 ( .A1(ram[4067]), .A2(n8724), .B1(n9274), .B2(n8926), .ZN(
        n8727) );
  INV_X1 U5013 ( .A(n8728), .ZN(n9262) );
  AOI22_X1 U5014 ( .A1(ram[4068]), .A2(n8724), .B1(n9274), .B2(n8950), .ZN(
        n8728) );
  INV_X1 U5015 ( .A(n8729), .ZN(n9263) );
  AOI22_X1 U5016 ( .A1(ram[4069]), .A2(n8724), .B1(n9274), .B2(n8974), .ZN(
        n8729) );
  INV_X1 U5017 ( .A(n8730), .ZN(n9264) );
  AOI22_X1 U5018 ( .A1(ram[4070]), .A2(n8724), .B1(n9274), .B2(n8998), .ZN(
        n8730) );
  INV_X1 U5019 ( .A(n8731), .ZN(n9265) );
  AOI22_X1 U5020 ( .A1(ram[4071]), .A2(n8724), .B1(n9274), .B2(n9022), .ZN(
        n8731) );
  INV_X1 U5021 ( .A(n8732), .ZN(n9266) );
  AOI22_X1 U5022 ( .A1(ram[4072]), .A2(n8724), .B1(n9274), .B2(n9046), .ZN(
        n8732) );
  INV_X1 U5023 ( .A(n8733), .ZN(n9267) );
  AOI22_X1 U5024 ( .A1(ram[4073]), .A2(n8724), .B1(n9274), .B2(n9070), .ZN(
        n8733) );
  INV_X1 U5025 ( .A(n8734), .ZN(n9268) );
  AOI22_X1 U5026 ( .A1(ram[4074]), .A2(n8724), .B1(n9274), .B2(n9094), .ZN(
        n8734) );
  INV_X1 U5027 ( .A(n8735), .ZN(n9269) );
  AOI22_X1 U5028 ( .A1(ram[4075]), .A2(n8724), .B1(n9274), .B2(n9118), .ZN(
        n8735) );
  INV_X1 U5029 ( .A(n8736), .ZN(n9270) );
  AOI22_X1 U5030 ( .A1(ram[4076]), .A2(n8724), .B1(n9274), .B2(n9142), .ZN(
        n8736) );
  INV_X1 U5031 ( .A(n8737), .ZN(n9271) );
  AOI22_X1 U5032 ( .A1(ram[4077]), .A2(n8724), .B1(n9274), .B2(n9166), .ZN(
        n8737) );
  INV_X1 U5033 ( .A(n8738), .ZN(n9272) );
  AOI22_X1 U5034 ( .A1(ram[4078]), .A2(n8724), .B1(n9274), .B2(n9190), .ZN(
        n8738) );
  INV_X1 U5035 ( .A(n8739), .ZN(n9273) );
  AOI22_X1 U5036 ( .A1(ram[4079]), .A2(n8724), .B1(n9274), .B2(n9214), .ZN(
        n8739) );
  INV_X1 U5037 ( .A(n4376), .ZN(n13559) );
  AOI22_X1 U5038 ( .A1(ram[16]), .A2(n4377), .B1(n13575), .B2(n8875), .ZN(
        n4376) );
  INV_X1 U5039 ( .A(n4378), .ZN(n13560) );
  AOI22_X1 U5040 ( .A1(ram[17]), .A2(n4377), .B1(n13575), .B2(n8899), .ZN(
        n4378) );
  INV_X1 U5041 ( .A(n4379), .ZN(n13561) );
  AOI22_X1 U5042 ( .A1(ram[18]), .A2(n4377), .B1(n13575), .B2(n8923), .ZN(
        n4379) );
  INV_X1 U5043 ( .A(n4380), .ZN(n13562) );
  AOI22_X1 U5044 ( .A1(ram[19]), .A2(n4377), .B1(n13575), .B2(n8947), .ZN(
        n4380) );
  INV_X1 U5045 ( .A(n4381), .ZN(n13563) );
  AOI22_X1 U5046 ( .A1(ram[20]), .A2(n4377), .B1(n13575), .B2(n8971), .ZN(
        n4381) );
  INV_X1 U5047 ( .A(n4382), .ZN(n13564) );
  AOI22_X1 U5048 ( .A1(ram[21]), .A2(n4377), .B1(n13575), .B2(n8995), .ZN(
        n4382) );
  INV_X1 U5049 ( .A(n4383), .ZN(n13565) );
  AOI22_X1 U5050 ( .A1(ram[22]), .A2(n4377), .B1(n13575), .B2(n9019), .ZN(
        n4383) );
  INV_X1 U5051 ( .A(n4384), .ZN(n13566) );
  AOI22_X1 U5052 ( .A1(ram[23]), .A2(n4377), .B1(n13575), .B2(n9043), .ZN(
        n4384) );
  INV_X1 U5053 ( .A(n4385), .ZN(n13567) );
  AOI22_X1 U5054 ( .A1(ram[24]), .A2(n4377), .B1(n13575), .B2(n9067), .ZN(
        n4385) );
  INV_X1 U5055 ( .A(n4386), .ZN(n13568) );
  AOI22_X1 U5056 ( .A1(ram[25]), .A2(n4377), .B1(n13575), .B2(n9091), .ZN(
        n4386) );
  INV_X1 U5057 ( .A(n4387), .ZN(n13569) );
  AOI22_X1 U5058 ( .A1(ram[26]), .A2(n4377), .B1(n13575), .B2(n9115), .ZN(
        n4387) );
  INV_X1 U5059 ( .A(n4388), .ZN(n13570) );
  AOI22_X1 U5060 ( .A1(ram[27]), .A2(n4377), .B1(n13575), .B2(n9139), .ZN(
        n4388) );
  INV_X1 U5061 ( .A(n4389), .ZN(n13571) );
  AOI22_X1 U5062 ( .A1(ram[28]), .A2(n4377), .B1(n13575), .B2(n9163), .ZN(
        n4389) );
  INV_X1 U5063 ( .A(n4390), .ZN(n13572) );
  AOI22_X1 U5064 ( .A1(ram[29]), .A2(n4377), .B1(n13575), .B2(n9187), .ZN(
        n4390) );
  INV_X1 U5065 ( .A(n4391), .ZN(n13573) );
  AOI22_X1 U5066 ( .A1(ram[30]), .A2(n4377), .B1(n13575), .B2(n9211), .ZN(
        n4391) );
  INV_X1 U5067 ( .A(n4392), .ZN(n13574) );
  AOI22_X1 U5068 ( .A1(ram[31]), .A2(n4377), .B1(n13575), .B2(n9235), .ZN(
        n4392) );
  INV_X1 U5069 ( .A(n4412), .ZN(n13525) );
  AOI22_X1 U5070 ( .A1(ram[48]), .A2(n4413), .B1(n13541), .B2(n8875), .ZN(
        n4412) );
  INV_X1 U5071 ( .A(n4414), .ZN(n13526) );
  AOI22_X1 U5072 ( .A1(ram[49]), .A2(n4413), .B1(n13541), .B2(n8899), .ZN(
        n4414) );
  INV_X1 U5073 ( .A(n4415), .ZN(n13527) );
  AOI22_X1 U5074 ( .A1(ram[50]), .A2(n4413), .B1(n13541), .B2(n8923), .ZN(
        n4415) );
  INV_X1 U5075 ( .A(n4416), .ZN(n13528) );
  AOI22_X1 U5076 ( .A1(ram[51]), .A2(n4413), .B1(n13541), .B2(n8947), .ZN(
        n4416) );
  INV_X1 U5077 ( .A(n4417), .ZN(n13529) );
  AOI22_X1 U5078 ( .A1(ram[52]), .A2(n4413), .B1(n13541), .B2(n8971), .ZN(
        n4417) );
  INV_X1 U5079 ( .A(n4418), .ZN(n13530) );
  AOI22_X1 U5080 ( .A1(ram[53]), .A2(n4413), .B1(n13541), .B2(n8995), .ZN(
        n4418) );
  INV_X1 U5081 ( .A(n4419), .ZN(n13531) );
  AOI22_X1 U5082 ( .A1(ram[54]), .A2(n4413), .B1(n13541), .B2(n9019), .ZN(
        n4419) );
  INV_X1 U5083 ( .A(n4420), .ZN(n13532) );
  AOI22_X1 U5084 ( .A1(ram[55]), .A2(n4413), .B1(n13541), .B2(n9043), .ZN(
        n4420) );
  INV_X1 U5085 ( .A(n4421), .ZN(n13533) );
  AOI22_X1 U5086 ( .A1(ram[56]), .A2(n4413), .B1(n13541), .B2(n9067), .ZN(
        n4421) );
  INV_X1 U5087 ( .A(n4422), .ZN(n13534) );
  AOI22_X1 U5088 ( .A1(ram[57]), .A2(n4413), .B1(n13541), .B2(n9091), .ZN(
        n4422) );
  INV_X1 U5089 ( .A(n4423), .ZN(n13535) );
  AOI22_X1 U5090 ( .A1(ram[58]), .A2(n4413), .B1(n13541), .B2(n9115), .ZN(
        n4423) );
  INV_X1 U5091 ( .A(n4424), .ZN(n13536) );
  AOI22_X1 U5092 ( .A1(ram[59]), .A2(n4413), .B1(n13541), .B2(n9139), .ZN(
        n4424) );
  INV_X1 U5093 ( .A(n4425), .ZN(n13537) );
  AOI22_X1 U5094 ( .A1(ram[60]), .A2(n4413), .B1(n13541), .B2(n9163), .ZN(
        n4425) );
  INV_X1 U5095 ( .A(n4426), .ZN(n13538) );
  AOI22_X1 U5096 ( .A1(ram[61]), .A2(n4413), .B1(n13541), .B2(n9187), .ZN(
        n4426) );
  INV_X1 U5097 ( .A(n4427), .ZN(n13539) );
  AOI22_X1 U5098 ( .A1(ram[62]), .A2(n4413), .B1(n13541), .B2(n9211), .ZN(
        n4427) );
  INV_X1 U5099 ( .A(n4428), .ZN(n13540) );
  AOI22_X1 U5100 ( .A1(ram[63]), .A2(n4413), .B1(n13541), .B2(n9235), .ZN(
        n4428) );
  INV_X1 U5101 ( .A(n4448), .ZN(n13491) );
  AOI22_X1 U5102 ( .A1(ram[80]), .A2(n4449), .B1(n13507), .B2(n8874), .ZN(
        n4448) );
  INV_X1 U5103 ( .A(n4450), .ZN(n13492) );
  AOI22_X1 U5104 ( .A1(ram[81]), .A2(n4449), .B1(n13507), .B2(n8898), .ZN(
        n4450) );
  INV_X1 U5105 ( .A(n4451), .ZN(n13493) );
  AOI22_X1 U5106 ( .A1(ram[82]), .A2(n4449), .B1(n13507), .B2(n8922), .ZN(
        n4451) );
  INV_X1 U5107 ( .A(n4452), .ZN(n13494) );
  AOI22_X1 U5108 ( .A1(ram[83]), .A2(n4449), .B1(n13507), .B2(n8946), .ZN(
        n4452) );
  INV_X1 U5109 ( .A(n4453), .ZN(n13495) );
  AOI22_X1 U5110 ( .A1(ram[84]), .A2(n4449), .B1(n13507), .B2(n8970), .ZN(
        n4453) );
  INV_X1 U5111 ( .A(n4454), .ZN(n13496) );
  AOI22_X1 U5112 ( .A1(ram[85]), .A2(n4449), .B1(n13507), .B2(n8994), .ZN(
        n4454) );
  INV_X1 U5113 ( .A(n4455), .ZN(n13497) );
  AOI22_X1 U5114 ( .A1(ram[86]), .A2(n4449), .B1(n13507), .B2(n9018), .ZN(
        n4455) );
  INV_X1 U5115 ( .A(n4456), .ZN(n13498) );
  AOI22_X1 U5116 ( .A1(ram[87]), .A2(n4449), .B1(n13507), .B2(n9042), .ZN(
        n4456) );
  INV_X1 U5117 ( .A(n4457), .ZN(n13499) );
  AOI22_X1 U5118 ( .A1(ram[88]), .A2(n4449), .B1(n13507), .B2(n9066), .ZN(
        n4457) );
  INV_X1 U5119 ( .A(n4458), .ZN(n13500) );
  AOI22_X1 U5120 ( .A1(ram[89]), .A2(n4449), .B1(n13507), .B2(n9090), .ZN(
        n4458) );
  INV_X1 U5121 ( .A(n4459), .ZN(n13501) );
  AOI22_X1 U5122 ( .A1(ram[90]), .A2(n4449), .B1(n13507), .B2(n9114), .ZN(
        n4459) );
  INV_X1 U5123 ( .A(n4460), .ZN(n13502) );
  AOI22_X1 U5124 ( .A1(ram[91]), .A2(n4449), .B1(n13507), .B2(n9138), .ZN(
        n4460) );
  INV_X1 U5125 ( .A(n4461), .ZN(n13503) );
  AOI22_X1 U5126 ( .A1(ram[92]), .A2(n4449), .B1(n13507), .B2(n9162), .ZN(
        n4461) );
  INV_X1 U5127 ( .A(n4462), .ZN(n13504) );
  AOI22_X1 U5128 ( .A1(ram[93]), .A2(n4449), .B1(n13507), .B2(n9186), .ZN(
        n4462) );
  INV_X1 U5129 ( .A(n4463), .ZN(n13505) );
  AOI22_X1 U5130 ( .A1(ram[94]), .A2(n4449), .B1(n13507), .B2(n9210), .ZN(
        n4463) );
  INV_X1 U5131 ( .A(n4464), .ZN(n13506) );
  AOI22_X1 U5132 ( .A1(ram[95]), .A2(n4449), .B1(n13507), .B2(n9234), .ZN(
        n4464) );
  INV_X1 U5133 ( .A(n4484), .ZN(n13457) );
  AOI22_X1 U5134 ( .A1(ram[112]), .A2(n4485), .B1(n13473), .B2(n8874), .ZN(
        n4484) );
  INV_X1 U5135 ( .A(n4486), .ZN(n13458) );
  AOI22_X1 U5136 ( .A1(ram[113]), .A2(n4485), .B1(n13473), .B2(n8898), .ZN(
        n4486) );
  INV_X1 U5137 ( .A(n4487), .ZN(n13459) );
  AOI22_X1 U5138 ( .A1(ram[114]), .A2(n4485), .B1(n13473), .B2(n8922), .ZN(
        n4487) );
  INV_X1 U5139 ( .A(n4488), .ZN(n13460) );
  AOI22_X1 U5140 ( .A1(ram[115]), .A2(n4485), .B1(n13473), .B2(n8946), .ZN(
        n4488) );
  INV_X1 U5141 ( .A(n4489), .ZN(n13461) );
  AOI22_X1 U5142 ( .A1(ram[116]), .A2(n4485), .B1(n13473), .B2(n8970), .ZN(
        n4489) );
  INV_X1 U5143 ( .A(n4490), .ZN(n13462) );
  AOI22_X1 U5144 ( .A1(ram[117]), .A2(n4485), .B1(n13473), .B2(n8994), .ZN(
        n4490) );
  INV_X1 U5145 ( .A(n4491), .ZN(n13463) );
  AOI22_X1 U5146 ( .A1(ram[118]), .A2(n4485), .B1(n13473), .B2(n9018), .ZN(
        n4491) );
  INV_X1 U5147 ( .A(n4492), .ZN(n13464) );
  AOI22_X1 U5148 ( .A1(ram[119]), .A2(n4485), .B1(n13473), .B2(n9042), .ZN(
        n4492) );
  INV_X1 U5149 ( .A(n4493), .ZN(n13465) );
  AOI22_X1 U5150 ( .A1(ram[120]), .A2(n4485), .B1(n13473), .B2(n9066), .ZN(
        n4493) );
  INV_X1 U5151 ( .A(n4494), .ZN(n13466) );
  AOI22_X1 U5152 ( .A1(ram[121]), .A2(n4485), .B1(n13473), .B2(n9090), .ZN(
        n4494) );
  INV_X1 U5153 ( .A(n4495), .ZN(n13467) );
  AOI22_X1 U5154 ( .A1(ram[122]), .A2(n4485), .B1(n13473), .B2(n9114), .ZN(
        n4495) );
  INV_X1 U5155 ( .A(n4496), .ZN(n13468) );
  AOI22_X1 U5156 ( .A1(ram[123]), .A2(n4485), .B1(n13473), .B2(n9138), .ZN(
        n4496) );
  INV_X1 U5157 ( .A(n4497), .ZN(n13469) );
  AOI22_X1 U5158 ( .A1(ram[124]), .A2(n4485), .B1(n13473), .B2(n9162), .ZN(
        n4497) );
  INV_X1 U5159 ( .A(n4498), .ZN(n13470) );
  AOI22_X1 U5160 ( .A1(ram[125]), .A2(n4485), .B1(n13473), .B2(n9186), .ZN(
        n4498) );
  INV_X1 U5161 ( .A(n4499), .ZN(n13471) );
  AOI22_X1 U5162 ( .A1(ram[126]), .A2(n4485), .B1(n13473), .B2(n9210), .ZN(
        n4499) );
  INV_X1 U5163 ( .A(n4500), .ZN(n13472) );
  AOI22_X1 U5164 ( .A1(ram[127]), .A2(n4485), .B1(n13473), .B2(n9234), .ZN(
        n4500) );
  INV_X1 U5165 ( .A(n4520), .ZN(n13423) );
  AOI22_X1 U5166 ( .A1(ram[144]), .A2(n4521), .B1(n13439), .B2(n8874), .ZN(
        n4520) );
  INV_X1 U5167 ( .A(n4522), .ZN(n13424) );
  AOI22_X1 U5168 ( .A1(ram[145]), .A2(n4521), .B1(n13439), .B2(n8898), .ZN(
        n4522) );
  INV_X1 U5169 ( .A(n4523), .ZN(n13425) );
  AOI22_X1 U5170 ( .A1(ram[146]), .A2(n4521), .B1(n13439), .B2(n8922), .ZN(
        n4523) );
  INV_X1 U5171 ( .A(n4524), .ZN(n13426) );
  AOI22_X1 U5172 ( .A1(ram[147]), .A2(n4521), .B1(n13439), .B2(n8946), .ZN(
        n4524) );
  INV_X1 U5173 ( .A(n4525), .ZN(n13427) );
  AOI22_X1 U5174 ( .A1(ram[148]), .A2(n4521), .B1(n13439), .B2(n8970), .ZN(
        n4525) );
  INV_X1 U5175 ( .A(n4526), .ZN(n13428) );
  AOI22_X1 U5176 ( .A1(ram[149]), .A2(n4521), .B1(n13439), .B2(n8994), .ZN(
        n4526) );
  INV_X1 U5177 ( .A(n4527), .ZN(n13429) );
  AOI22_X1 U5178 ( .A1(ram[150]), .A2(n4521), .B1(n13439), .B2(n9018), .ZN(
        n4527) );
  INV_X1 U5179 ( .A(n4528), .ZN(n13430) );
  AOI22_X1 U5180 ( .A1(ram[151]), .A2(n4521), .B1(n13439), .B2(n9042), .ZN(
        n4528) );
  INV_X1 U5181 ( .A(n4529), .ZN(n13431) );
  AOI22_X1 U5182 ( .A1(ram[152]), .A2(n4521), .B1(n13439), .B2(n9066), .ZN(
        n4529) );
  INV_X1 U5183 ( .A(n4530), .ZN(n13432) );
  AOI22_X1 U5184 ( .A1(ram[153]), .A2(n4521), .B1(n13439), .B2(n9090), .ZN(
        n4530) );
  INV_X1 U5185 ( .A(n4531), .ZN(n13433) );
  AOI22_X1 U5186 ( .A1(ram[154]), .A2(n4521), .B1(n13439), .B2(n9114), .ZN(
        n4531) );
  INV_X1 U5187 ( .A(n4532), .ZN(n13434) );
  AOI22_X1 U5188 ( .A1(ram[155]), .A2(n4521), .B1(n13439), .B2(n9138), .ZN(
        n4532) );
  INV_X1 U5189 ( .A(n4533), .ZN(n13435) );
  AOI22_X1 U5190 ( .A1(ram[156]), .A2(n4521), .B1(n13439), .B2(n9162), .ZN(
        n4533) );
  INV_X1 U5191 ( .A(n4534), .ZN(n13436) );
  AOI22_X1 U5192 ( .A1(ram[157]), .A2(n4521), .B1(n13439), .B2(n9186), .ZN(
        n4534) );
  INV_X1 U5193 ( .A(n4535), .ZN(n13437) );
  AOI22_X1 U5194 ( .A1(ram[158]), .A2(n4521), .B1(n13439), .B2(n9210), .ZN(
        n4535) );
  INV_X1 U5195 ( .A(n4536), .ZN(n13438) );
  AOI22_X1 U5196 ( .A1(ram[159]), .A2(n4521), .B1(n13439), .B2(n9234), .ZN(
        n4536) );
  INV_X1 U5197 ( .A(n4556), .ZN(n13389) );
  AOI22_X1 U5198 ( .A1(ram[176]), .A2(n4557), .B1(n13405), .B2(n8874), .ZN(
        n4556) );
  INV_X1 U5199 ( .A(n4558), .ZN(n13390) );
  AOI22_X1 U5200 ( .A1(ram[177]), .A2(n4557), .B1(n13405), .B2(n8898), .ZN(
        n4558) );
  INV_X1 U5201 ( .A(n4559), .ZN(n13391) );
  AOI22_X1 U5202 ( .A1(ram[178]), .A2(n4557), .B1(n13405), .B2(n8922), .ZN(
        n4559) );
  INV_X1 U5203 ( .A(n4560), .ZN(n13392) );
  AOI22_X1 U5204 ( .A1(ram[179]), .A2(n4557), .B1(n13405), .B2(n8946), .ZN(
        n4560) );
  INV_X1 U5205 ( .A(n4561), .ZN(n13393) );
  AOI22_X1 U5206 ( .A1(ram[180]), .A2(n4557), .B1(n13405), .B2(n8970), .ZN(
        n4561) );
  INV_X1 U5207 ( .A(n4562), .ZN(n13394) );
  AOI22_X1 U5208 ( .A1(ram[181]), .A2(n4557), .B1(n13405), .B2(n8994), .ZN(
        n4562) );
  INV_X1 U5209 ( .A(n4563), .ZN(n13395) );
  AOI22_X1 U5210 ( .A1(ram[182]), .A2(n4557), .B1(n13405), .B2(n9018), .ZN(
        n4563) );
  INV_X1 U5211 ( .A(n4564), .ZN(n13396) );
  AOI22_X1 U5212 ( .A1(ram[183]), .A2(n4557), .B1(n13405), .B2(n9042), .ZN(
        n4564) );
  INV_X1 U5213 ( .A(n4565), .ZN(n13397) );
  AOI22_X1 U5214 ( .A1(ram[184]), .A2(n4557), .B1(n13405), .B2(n9066), .ZN(
        n4565) );
  INV_X1 U5215 ( .A(n4566), .ZN(n13398) );
  AOI22_X1 U5216 ( .A1(ram[185]), .A2(n4557), .B1(n13405), .B2(n9090), .ZN(
        n4566) );
  INV_X1 U5217 ( .A(n4567), .ZN(n13399) );
  AOI22_X1 U5218 ( .A1(ram[186]), .A2(n4557), .B1(n13405), .B2(n9114), .ZN(
        n4567) );
  INV_X1 U5219 ( .A(n4568), .ZN(n13400) );
  AOI22_X1 U5220 ( .A1(ram[187]), .A2(n4557), .B1(n13405), .B2(n9138), .ZN(
        n4568) );
  INV_X1 U5221 ( .A(n4569), .ZN(n13401) );
  AOI22_X1 U5222 ( .A1(ram[188]), .A2(n4557), .B1(n13405), .B2(n9162), .ZN(
        n4569) );
  INV_X1 U5223 ( .A(n4570), .ZN(n13402) );
  AOI22_X1 U5224 ( .A1(ram[189]), .A2(n4557), .B1(n13405), .B2(n9186), .ZN(
        n4570) );
  INV_X1 U5225 ( .A(n4571), .ZN(n13403) );
  AOI22_X1 U5226 ( .A1(ram[190]), .A2(n4557), .B1(n13405), .B2(n9210), .ZN(
        n4571) );
  INV_X1 U5227 ( .A(n4572), .ZN(n13404) );
  AOI22_X1 U5228 ( .A1(ram[191]), .A2(n4557), .B1(n13405), .B2(n9234), .ZN(
        n4572) );
  INV_X1 U5229 ( .A(n4592), .ZN(n13355) );
  AOI22_X1 U5230 ( .A1(ram[208]), .A2(n4593), .B1(n13371), .B2(n8874), .ZN(
        n4592) );
  INV_X1 U5231 ( .A(n4594), .ZN(n13356) );
  AOI22_X1 U5232 ( .A1(ram[209]), .A2(n4593), .B1(n13371), .B2(n8898), .ZN(
        n4594) );
  INV_X1 U5233 ( .A(n4595), .ZN(n13357) );
  AOI22_X1 U5234 ( .A1(ram[210]), .A2(n4593), .B1(n13371), .B2(n8922), .ZN(
        n4595) );
  INV_X1 U5235 ( .A(n4596), .ZN(n13358) );
  AOI22_X1 U5236 ( .A1(ram[211]), .A2(n4593), .B1(n13371), .B2(n8946), .ZN(
        n4596) );
  INV_X1 U5237 ( .A(n4597), .ZN(n13359) );
  AOI22_X1 U5238 ( .A1(ram[212]), .A2(n4593), .B1(n13371), .B2(n8970), .ZN(
        n4597) );
  INV_X1 U5239 ( .A(n4598), .ZN(n13360) );
  AOI22_X1 U5240 ( .A1(ram[213]), .A2(n4593), .B1(n13371), .B2(n8994), .ZN(
        n4598) );
  INV_X1 U5241 ( .A(n4599), .ZN(n13361) );
  AOI22_X1 U5242 ( .A1(ram[214]), .A2(n4593), .B1(n13371), .B2(n9018), .ZN(
        n4599) );
  INV_X1 U5243 ( .A(n4600), .ZN(n13362) );
  AOI22_X1 U5244 ( .A1(ram[215]), .A2(n4593), .B1(n13371), .B2(n9042), .ZN(
        n4600) );
  INV_X1 U5245 ( .A(n4601), .ZN(n13363) );
  AOI22_X1 U5246 ( .A1(ram[216]), .A2(n4593), .B1(n13371), .B2(n9066), .ZN(
        n4601) );
  INV_X1 U5247 ( .A(n4602), .ZN(n13364) );
  AOI22_X1 U5248 ( .A1(ram[217]), .A2(n4593), .B1(n13371), .B2(n9090), .ZN(
        n4602) );
  INV_X1 U5249 ( .A(n4603), .ZN(n13365) );
  AOI22_X1 U5250 ( .A1(ram[218]), .A2(n4593), .B1(n13371), .B2(n9114), .ZN(
        n4603) );
  INV_X1 U5251 ( .A(n4604), .ZN(n13366) );
  AOI22_X1 U5252 ( .A1(ram[219]), .A2(n4593), .B1(n13371), .B2(n9138), .ZN(
        n4604) );
  INV_X1 U5253 ( .A(n4605), .ZN(n13367) );
  AOI22_X1 U5254 ( .A1(ram[220]), .A2(n4593), .B1(n13371), .B2(n9162), .ZN(
        n4605) );
  INV_X1 U5255 ( .A(n4606), .ZN(n13368) );
  AOI22_X1 U5256 ( .A1(ram[221]), .A2(n4593), .B1(n13371), .B2(n9186), .ZN(
        n4606) );
  INV_X1 U5257 ( .A(n4607), .ZN(n13369) );
  AOI22_X1 U5258 ( .A1(ram[222]), .A2(n4593), .B1(n13371), .B2(n9210), .ZN(
        n4607) );
  INV_X1 U5259 ( .A(n4608), .ZN(n13370) );
  AOI22_X1 U5260 ( .A1(ram[223]), .A2(n4593), .B1(n13371), .B2(n9234), .ZN(
        n4608) );
  INV_X1 U5261 ( .A(n4628), .ZN(n13321) );
  AOI22_X1 U5262 ( .A1(ram[240]), .A2(n4629), .B1(n13337), .B2(n8874), .ZN(
        n4628) );
  INV_X1 U5263 ( .A(n4630), .ZN(n13322) );
  AOI22_X1 U5264 ( .A1(ram[241]), .A2(n4629), .B1(n13337), .B2(n8898), .ZN(
        n4630) );
  INV_X1 U5265 ( .A(n4631), .ZN(n13323) );
  AOI22_X1 U5266 ( .A1(ram[242]), .A2(n4629), .B1(n13337), .B2(n8922), .ZN(
        n4631) );
  INV_X1 U5267 ( .A(n4632), .ZN(n13324) );
  AOI22_X1 U5268 ( .A1(ram[243]), .A2(n4629), .B1(n13337), .B2(n8946), .ZN(
        n4632) );
  INV_X1 U5269 ( .A(n4633), .ZN(n13325) );
  AOI22_X1 U5270 ( .A1(ram[244]), .A2(n4629), .B1(n13337), .B2(n8970), .ZN(
        n4633) );
  INV_X1 U5271 ( .A(n4634), .ZN(n13326) );
  AOI22_X1 U5272 ( .A1(ram[245]), .A2(n4629), .B1(n13337), .B2(n8994), .ZN(
        n4634) );
  INV_X1 U5273 ( .A(n4635), .ZN(n13327) );
  AOI22_X1 U5274 ( .A1(ram[246]), .A2(n4629), .B1(n13337), .B2(n9018), .ZN(
        n4635) );
  INV_X1 U5275 ( .A(n4636), .ZN(n13328) );
  AOI22_X1 U5276 ( .A1(ram[247]), .A2(n4629), .B1(n13337), .B2(n9042), .ZN(
        n4636) );
  INV_X1 U5277 ( .A(n4637), .ZN(n13329) );
  AOI22_X1 U5278 ( .A1(ram[248]), .A2(n4629), .B1(n13337), .B2(n9066), .ZN(
        n4637) );
  INV_X1 U5279 ( .A(n4638), .ZN(n13330) );
  AOI22_X1 U5280 ( .A1(ram[249]), .A2(n4629), .B1(n13337), .B2(n9090), .ZN(
        n4638) );
  INV_X1 U5281 ( .A(n4639), .ZN(n13331) );
  AOI22_X1 U5282 ( .A1(ram[250]), .A2(n4629), .B1(n13337), .B2(n9114), .ZN(
        n4639) );
  INV_X1 U5283 ( .A(n4640), .ZN(n13332) );
  AOI22_X1 U5284 ( .A1(ram[251]), .A2(n4629), .B1(n13337), .B2(n9138), .ZN(
        n4640) );
  INV_X1 U5285 ( .A(n4641), .ZN(n13333) );
  AOI22_X1 U5286 ( .A1(ram[252]), .A2(n4629), .B1(n13337), .B2(n9162), .ZN(
        n4641) );
  INV_X1 U5287 ( .A(n4642), .ZN(n13334) );
  AOI22_X1 U5288 ( .A1(ram[253]), .A2(n4629), .B1(n13337), .B2(n9186), .ZN(
        n4642) );
  INV_X1 U5289 ( .A(n4643), .ZN(n13335) );
  AOI22_X1 U5290 ( .A1(ram[254]), .A2(n4629), .B1(n13337), .B2(n9210), .ZN(
        n4643) );
  INV_X1 U5291 ( .A(n4644), .ZN(n13336) );
  AOI22_X1 U5292 ( .A1(ram[255]), .A2(n4629), .B1(n13337), .B2(n9234), .ZN(
        n4644) );
  INV_X1 U5293 ( .A(n4666), .ZN(n13287) );
  AOI22_X1 U5294 ( .A1(ram[272]), .A2(n4667), .B1(n13303), .B2(n8873), .ZN(
        n4666) );
  INV_X1 U5295 ( .A(n4668), .ZN(n13288) );
  AOI22_X1 U5296 ( .A1(ram[273]), .A2(n4667), .B1(n13303), .B2(n8897), .ZN(
        n4668) );
  INV_X1 U5297 ( .A(n4669), .ZN(n13289) );
  AOI22_X1 U5298 ( .A1(ram[274]), .A2(n4667), .B1(n13303), .B2(n8921), .ZN(
        n4669) );
  INV_X1 U5299 ( .A(n4670), .ZN(n13290) );
  AOI22_X1 U5300 ( .A1(ram[275]), .A2(n4667), .B1(n13303), .B2(n8945), .ZN(
        n4670) );
  INV_X1 U5301 ( .A(n4671), .ZN(n13291) );
  AOI22_X1 U5302 ( .A1(ram[276]), .A2(n4667), .B1(n13303), .B2(n8969), .ZN(
        n4671) );
  INV_X1 U5303 ( .A(n4672), .ZN(n13292) );
  AOI22_X1 U5304 ( .A1(ram[277]), .A2(n4667), .B1(n13303), .B2(n8993), .ZN(
        n4672) );
  INV_X1 U5305 ( .A(n4673), .ZN(n13293) );
  AOI22_X1 U5306 ( .A1(ram[278]), .A2(n4667), .B1(n13303), .B2(n9017), .ZN(
        n4673) );
  INV_X1 U5307 ( .A(n4674), .ZN(n13294) );
  AOI22_X1 U5308 ( .A1(ram[279]), .A2(n4667), .B1(n13303), .B2(n9041), .ZN(
        n4674) );
  INV_X1 U5309 ( .A(n4675), .ZN(n13295) );
  AOI22_X1 U5310 ( .A1(ram[280]), .A2(n4667), .B1(n13303), .B2(n9065), .ZN(
        n4675) );
  INV_X1 U5311 ( .A(n4676), .ZN(n13296) );
  AOI22_X1 U5312 ( .A1(ram[281]), .A2(n4667), .B1(n13303), .B2(n9089), .ZN(
        n4676) );
  INV_X1 U5313 ( .A(n4677), .ZN(n13297) );
  AOI22_X1 U5314 ( .A1(ram[282]), .A2(n4667), .B1(n13303), .B2(n9113), .ZN(
        n4677) );
  INV_X1 U5315 ( .A(n4678), .ZN(n13298) );
  AOI22_X1 U5316 ( .A1(ram[283]), .A2(n4667), .B1(n13303), .B2(n9137), .ZN(
        n4678) );
  INV_X1 U5317 ( .A(n4679), .ZN(n13299) );
  AOI22_X1 U5318 ( .A1(ram[284]), .A2(n4667), .B1(n13303), .B2(n9161), .ZN(
        n4679) );
  INV_X1 U5319 ( .A(n4680), .ZN(n13300) );
  AOI22_X1 U5320 ( .A1(ram[285]), .A2(n4667), .B1(n13303), .B2(n9185), .ZN(
        n4680) );
  INV_X1 U5321 ( .A(n4681), .ZN(n13301) );
  AOI22_X1 U5322 ( .A1(ram[286]), .A2(n4667), .B1(n13303), .B2(n9209), .ZN(
        n4681) );
  INV_X1 U5323 ( .A(n4682), .ZN(n13302) );
  AOI22_X1 U5324 ( .A1(ram[287]), .A2(n4667), .B1(n13303), .B2(n9233), .ZN(
        n4682) );
  INV_X1 U5325 ( .A(n4700), .ZN(n13253) );
  AOI22_X1 U5326 ( .A1(ram[304]), .A2(n4701), .B1(n13269), .B2(n8873), .ZN(
        n4700) );
  INV_X1 U5327 ( .A(n4702), .ZN(n13254) );
  AOI22_X1 U5328 ( .A1(ram[305]), .A2(n4701), .B1(n13269), .B2(n8897), .ZN(
        n4702) );
  INV_X1 U5329 ( .A(n4703), .ZN(n13255) );
  AOI22_X1 U5330 ( .A1(ram[306]), .A2(n4701), .B1(n13269), .B2(n8921), .ZN(
        n4703) );
  INV_X1 U5331 ( .A(n4704), .ZN(n13256) );
  AOI22_X1 U5332 ( .A1(ram[307]), .A2(n4701), .B1(n13269), .B2(n8945), .ZN(
        n4704) );
  INV_X1 U5333 ( .A(n4705), .ZN(n13257) );
  AOI22_X1 U5334 ( .A1(ram[308]), .A2(n4701), .B1(n13269), .B2(n8969), .ZN(
        n4705) );
  INV_X1 U5335 ( .A(n4706), .ZN(n13258) );
  AOI22_X1 U5336 ( .A1(ram[309]), .A2(n4701), .B1(n13269), .B2(n8993), .ZN(
        n4706) );
  INV_X1 U5337 ( .A(n4707), .ZN(n13259) );
  AOI22_X1 U5338 ( .A1(ram[310]), .A2(n4701), .B1(n13269), .B2(n9017), .ZN(
        n4707) );
  INV_X1 U5339 ( .A(n4708), .ZN(n13260) );
  AOI22_X1 U5340 ( .A1(ram[311]), .A2(n4701), .B1(n13269), .B2(n9041), .ZN(
        n4708) );
  INV_X1 U5341 ( .A(n4709), .ZN(n13261) );
  AOI22_X1 U5342 ( .A1(ram[312]), .A2(n4701), .B1(n13269), .B2(n9065), .ZN(
        n4709) );
  INV_X1 U5343 ( .A(n4710), .ZN(n13262) );
  AOI22_X1 U5344 ( .A1(ram[313]), .A2(n4701), .B1(n13269), .B2(n9089), .ZN(
        n4710) );
  INV_X1 U5345 ( .A(n4711), .ZN(n13263) );
  AOI22_X1 U5346 ( .A1(ram[314]), .A2(n4701), .B1(n13269), .B2(n9113), .ZN(
        n4711) );
  INV_X1 U5347 ( .A(n4712), .ZN(n13264) );
  AOI22_X1 U5348 ( .A1(ram[315]), .A2(n4701), .B1(n13269), .B2(n9137), .ZN(
        n4712) );
  INV_X1 U5349 ( .A(n4713), .ZN(n13265) );
  AOI22_X1 U5350 ( .A1(ram[316]), .A2(n4701), .B1(n13269), .B2(n9161), .ZN(
        n4713) );
  INV_X1 U5351 ( .A(n4714), .ZN(n13266) );
  AOI22_X1 U5352 ( .A1(ram[317]), .A2(n4701), .B1(n13269), .B2(n9185), .ZN(
        n4714) );
  INV_X1 U5353 ( .A(n4715), .ZN(n13267) );
  AOI22_X1 U5354 ( .A1(ram[318]), .A2(n4701), .B1(n13269), .B2(n9209), .ZN(
        n4715) );
  INV_X1 U5355 ( .A(n4716), .ZN(n13268) );
  AOI22_X1 U5356 ( .A1(ram[319]), .A2(n4701), .B1(n13269), .B2(n9233), .ZN(
        n4716) );
  INV_X1 U5357 ( .A(n4734), .ZN(n13219) );
  AOI22_X1 U5358 ( .A1(ram[336]), .A2(n4735), .B1(n13235), .B2(n8873), .ZN(
        n4734) );
  INV_X1 U5359 ( .A(n4736), .ZN(n13220) );
  AOI22_X1 U5360 ( .A1(ram[337]), .A2(n4735), .B1(n13235), .B2(n8897), .ZN(
        n4736) );
  INV_X1 U5361 ( .A(n4737), .ZN(n13221) );
  AOI22_X1 U5362 ( .A1(ram[338]), .A2(n4735), .B1(n13235), .B2(n8921), .ZN(
        n4737) );
  INV_X1 U5363 ( .A(n4738), .ZN(n13222) );
  AOI22_X1 U5364 ( .A1(ram[339]), .A2(n4735), .B1(n13235), .B2(n8945), .ZN(
        n4738) );
  INV_X1 U5365 ( .A(n4739), .ZN(n13223) );
  AOI22_X1 U5366 ( .A1(ram[340]), .A2(n4735), .B1(n13235), .B2(n8969), .ZN(
        n4739) );
  INV_X1 U5367 ( .A(n4740), .ZN(n13224) );
  AOI22_X1 U5368 ( .A1(ram[341]), .A2(n4735), .B1(n13235), .B2(n8993), .ZN(
        n4740) );
  INV_X1 U5369 ( .A(n4741), .ZN(n13225) );
  AOI22_X1 U5370 ( .A1(ram[342]), .A2(n4735), .B1(n13235), .B2(n9017), .ZN(
        n4741) );
  INV_X1 U5371 ( .A(n4742), .ZN(n13226) );
  AOI22_X1 U5372 ( .A1(ram[343]), .A2(n4735), .B1(n13235), .B2(n9041), .ZN(
        n4742) );
  INV_X1 U5373 ( .A(n4743), .ZN(n13227) );
  AOI22_X1 U5374 ( .A1(ram[344]), .A2(n4735), .B1(n13235), .B2(n9065), .ZN(
        n4743) );
  INV_X1 U5375 ( .A(n4744), .ZN(n13228) );
  AOI22_X1 U5376 ( .A1(ram[345]), .A2(n4735), .B1(n13235), .B2(n9089), .ZN(
        n4744) );
  INV_X1 U5377 ( .A(n4745), .ZN(n13229) );
  AOI22_X1 U5378 ( .A1(ram[346]), .A2(n4735), .B1(n13235), .B2(n9113), .ZN(
        n4745) );
  INV_X1 U5379 ( .A(n4746), .ZN(n13230) );
  AOI22_X1 U5380 ( .A1(ram[347]), .A2(n4735), .B1(n13235), .B2(n9137), .ZN(
        n4746) );
  INV_X1 U5381 ( .A(n4747), .ZN(n13231) );
  AOI22_X1 U5382 ( .A1(ram[348]), .A2(n4735), .B1(n13235), .B2(n9161), .ZN(
        n4747) );
  INV_X1 U5383 ( .A(n4748), .ZN(n13232) );
  AOI22_X1 U5384 ( .A1(ram[349]), .A2(n4735), .B1(n13235), .B2(n9185), .ZN(
        n4748) );
  INV_X1 U5385 ( .A(n4749), .ZN(n13233) );
  AOI22_X1 U5386 ( .A1(ram[350]), .A2(n4735), .B1(n13235), .B2(n9209), .ZN(
        n4749) );
  INV_X1 U5387 ( .A(n4750), .ZN(n13234) );
  AOI22_X1 U5388 ( .A1(ram[351]), .A2(n4735), .B1(n13235), .B2(n9233), .ZN(
        n4750) );
  INV_X1 U5389 ( .A(n4768), .ZN(n13185) );
  AOI22_X1 U5390 ( .A1(ram[368]), .A2(n4769), .B1(n13201), .B2(n8873), .ZN(
        n4768) );
  INV_X1 U5391 ( .A(n4770), .ZN(n13186) );
  AOI22_X1 U5392 ( .A1(ram[369]), .A2(n4769), .B1(n13201), .B2(n8897), .ZN(
        n4770) );
  INV_X1 U5393 ( .A(n4771), .ZN(n13187) );
  AOI22_X1 U5394 ( .A1(ram[370]), .A2(n4769), .B1(n13201), .B2(n8921), .ZN(
        n4771) );
  INV_X1 U5395 ( .A(n4772), .ZN(n13188) );
  AOI22_X1 U5396 ( .A1(ram[371]), .A2(n4769), .B1(n13201), .B2(n8945), .ZN(
        n4772) );
  INV_X1 U5397 ( .A(n4773), .ZN(n13189) );
  AOI22_X1 U5398 ( .A1(ram[372]), .A2(n4769), .B1(n13201), .B2(n8969), .ZN(
        n4773) );
  INV_X1 U5399 ( .A(n4774), .ZN(n13190) );
  AOI22_X1 U5400 ( .A1(ram[373]), .A2(n4769), .B1(n13201), .B2(n8993), .ZN(
        n4774) );
  INV_X1 U5401 ( .A(n4775), .ZN(n13191) );
  AOI22_X1 U5402 ( .A1(ram[374]), .A2(n4769), .B1(n13201), .B2(n9017), .ZN(
        n4775) );
  INV_X1 U5403 ( .A(n4776), .ZN(n13192) );
  AOI22_X1 U5404 ( .A1(ram[375]), .A2(n4769), .B1(n13201), .B2(n9041), .ZN(
        n4776) );
  INV_X1 U5405 ( .A(n4777), .ZN(n13193) );
  AOI22_X1 U5406 ( .A1(ram[376]), .A2(n4769), .B1(n13201), .B2(n9065), .ZN(
        n4777) );
  INV_X1 U5407 ( .A(n4778), .ZN(n13194) );
  AOI22_X1 U5408 ( .A1(ram[377]), .A2(n4769), .B1(n13201), .B2(n9089), .ZN(
        n4778) );
  INV_X1 U5409 ( .A(n4779), .ZN(n13195) );
  AOI22_X1 U5410 ( .A1(ram[378]), .A2(n4769), .B1(n13201), .B2(n9113), .ZN(
        n4779) );
  INV_X1 U5411 ( .A(n4780), .ZN(n13196) );
  AOI22_X1 U5412 ( .A1(ram[379]), .A2(n4769), .B1(n13201), .B2(n9137), .ZN(
        n4780) );
  INV_X1 U5413 ( .A(n4781), .ZN(n13197) );
  AOI22_X1 U5414 ( .A1(ram[380]), .A2(n4769), .B1(n13201), .B2(n9161), .ZN(
        n4781) );
  INV_X1 U5415 ( .A(n4782), .ZN(n13198) );
  AOI22_X1 U5416 ( .A1(ram[381]), .A2(n4769), .B1(n13201), .B2(n9185), .ZN(
        n4782) );
  INV_X1 U5417 ( .A(n4783), .ZN(n13199) );
  AOI22_X1 U5418 ( .A1(ram[382]), .A2(n4769), .B1(n13201), .B2(n9209), .ZN(
        n4783) );
  INV_X1 U5419 ( .A(n4784), .ZN(n13200) );
  AOI22_X1 U5420 ( .A1(ram[383]), .A2(n4769), .B1(n13201), .B2(n9233), .ZN(
        n4784) );
  INV_X1 U5421 ( .A(n4802), .ZN(n13151) );
  AOI22_X1 U5422 ( .A1(ram[400]), .A2(n4803), .B1(n13167), .B2(n8873), .ZN(
        n4802) );
  INV_X1 U5423 ( .A(n4804), .ZN(n13152) );
  AOI22_X1 U5424 ( .A1(ram[401]), .A2(n4803), .B1(n13167), .B2(n8897), .ZN(
        n4804) );
  INV_X1 U5425 ( .A(n4805), .ZN(n13153) );
  AOI22_X1 U5426 ( .A1(ram[402]), .A2(n4803), .B1(n13167), .B2(n8921), .ZN(
        n4805) );
  INV_X1 U5427 ( .A(n4806), .ZN(n13154) );
  AOI22_X1 U5428 ( .A1(ram[403]), .A2(n4803), .B1(n13167), .B2(n8945), .ZN(
        n4806) );
  INV_X1 U5429 ( .A(n4807), .ZN(n13155) );
  AOI22_X1 U5430 ( .A1(ram[404]), .A2(n4803), .B1(n13167), .B2(n8969), .ZN(
        n4807) );
  INV_X1 U5431 ( .A(n4808), .ZN(n13156) );
  AOI22_X1 U5432 ( .A1(ram[405]), .A2(n4803), .B1(n13167), .B2(n8993), .ZN(
        n4808) );
  INV_X1 U5433 ( .A(n4809), .ZN(n13157) );
  AOI22_X1 U5434 ( .A1(ram[406]), .A2(n4803), .B1(n13167), .B2(n9017), .ZN(
        n4809) );
  INV_X1 U5435 ( .A(n4810), .ZN(n13158) );
  AOI22_X1 U5436 ( .A1(ram[407]), .A2(n4803), .B1(n13167), .B2(n9041), .ZN(
        n4810) );
  INV_X1 U5437 ( .A(n4811), .ZN(n13159) );
  AOI22_X1 U5438 ( .A1(ram[408]), .A2(n4803), .B1(n13167), .B2(n9065), .ZN(
        n4811) );
  INV_X1 U5439 ( .A(n4812), .ZN(n13160) );
  AOI22_X1 U5440 ( .A1(ram[409]), .A2(n4803), .B1(n13167), .B2(n9089), .ZN(
        n4812) );
  INV_X1 U5441 ( .A(n4813), .ZN(n13161) );
  AOI22_X1 U5442 ( .A1(ram[410]), .A2(n4803), .B1(n13167), .B2(n9113), .ZN(
        n4813) );
  INV_X1 U5443 ( .A(n4814), .ZN(n13162) );
  AOI22_X1 U5444 ( .A1(ram[411]), .A2(n4803), .B1(n13167), .B2(n9137), .ZN(
        n4814) );
  INV_X1 U5445 ( .A(n4815), .ZN(n13163) );
  AOI22_X1 U5446 ( .A1(ram[412]), .A2(n4803), .B1(n13167), .B2(n9161), .ZN(
        n4815) );
  INV_X1 U5447 ( .A(n4816), .ZN(n13164) );
  AOI22_X1 U5448 ( .A1(ram[413]), .A2(n4803), .B1(n13167), .B2(n9185), .ZN(
        n4816) );
  INV_X1 U5449 ( .A(n4817), .ZN(n13165) );
  AOI22_X1 U5450 ( .A1(ram[414]), .A2(n4803), .B1(n13167), .B2(n9209), .ZN(
        n4817) );
  INV_X1 U5451 ( .A(n4818), .ZN(n13166) );
  AOI22_X1 U5452 ( .A1(ram[415]), .A2(n4803), .B1(n13167), .B2(n9233), .ZN(
        n4818) );
  INV_X1 U5453 ( .A(n4836), .ZN(n13117) );
  AOI22_X1 U5454 ( .A1(ram[432]), .A2(n4837), .B1(n13133), .B2(n8873), .ZN(
        n4836) );
  INV_X1 U5455 ( .A(n4838), .ZN(n13118) );
  AOI22_X1 U5456 ( .A1(ram[433]), .A2(n4837), .B1(n13133), .B2(n8897), .ZN(
        n4838) );
  INV_X1 U5457 ( .A(n4839), .ZN(n13119) );
  AOI22_X1 U5458 ( .A1(ram[434]), .A2(n4837), .B1(n13133), .B2(n8921), .ZN(
        n4839) );
  INV_X1 U5459 ( .A(n4840), .ZN(n13120) );
  AOI22_X1 U5460 ( .A1(ram[435]), .A2(n4837), .B1(n13133), .B2(n8945), .ZN(
        n4840) );
  INV_X1 U5461 ( .A(n4841), .ZN(n13121) );
  AOI22_X1 U5462 ( .A1(ram[436]), .A2(n4837), .B1(n13133), .B2(n8969), .ZN(
        n4841) );
  INV_X1 U5463 ( .A(n4842), .ZN(n13122) );
  AOI22_X1 U5464 ( .A1(ram[437]), .A2(n4837), .B1(n13133), .B2(n8993), .ZN(
        n4842) );
  INV_X1 U5465 ( .A(n4843), .ZN(n13123) );
  AOI22_X1 U5466 ( .A1(ram[438]), .A2(n4837), .B1(n13133), .B2(n9017), .ZN(
        n4843) );
  INV_X1 U5467 ( .A(n4844), .ZN(n13124) );
  AOI22_X1 U5468 ( .A1(ram[439]), .A2(n4837), .B1(n13133), .B2(n9041), .ZN(
        n4844) );
  INV_X1 U5469 ( .A(n4845), .ZN(n13125) );
  AOI22_X1 U5470 ( .A1(ram[440]), .A2(n4837), .B1(n13133), .B2(n9065), .ZN(
        n4845) );
  INV_X1 U5471 ( .A(n4846), .ZN(n13126) );
  AOI22_X1 U5472 ( .A1(ram[441]), .A2(n4837), .B1(n13133), .B2(n9089), .ZN(
        n4846) );
  INV_X1 U5473 ( .A(n4847), .ZN(n13127) );
  AOI22_X1 U5474 ( .A1(ram[442]), .A2(n4837), .B1(n13133), .B2(n9113), .ZN(
        n4847) );
  INV_X1 U5475 ( .A(n4848), .ZN(n13128) );
  AOI22_X1 U5476 ( .A1(ram[443]), .A2(n4837), .B1(n13133), .B2(n9137), .ZN(
        n4848) );
  INV_X1 U5477 ( .A(n4849), .ZN(n13129) );
  AOI22_X1 U5478 ( .A1(ram[444]), .A2(n4837), .B1(n13133), .B2(n9161), .ZN(
        n4849) );
  INV_X1 U5479 ( .A(n4850), .ZN(n13130) );
  AOI22_X1 U5480 ( .A1(ram[445]), .A2(n4837), .B1(n13133), .B2(n9185), .ZN(
        n4850) );
  INV_X1 U5481 ( .A(n4851), .ZN(n13131) );
  AOI22_X1 U5482 ( .A1(ram[446]), .A2(n4837), .B1(n13133), .B2(n9209), .ZN(
        n4851) );
  INV_X1 U5483 ( .A(n4852), .ZN(n13132) );
  AOI22_X1 U5484 ( .A1(ram[447]), .A2(n4837), .B1(n13133), .B2(n9233), .ZN(
        n4852) );
  INV_X1 U5485 ( .A(n4870), .ZN(n13083) );
  AOI22_X1 U5486 ( .A1(ram[464]), .A2(n4871), .B1(n13099), .B2(n8872), .ZN(
        n4870) );
  INV_X1 U5487 ( .A(n4872), .ZN(n13084) );
  AOI22_X1 U5488 ( .A1(ram[465]), .A2(n4871), .B1(n13099), .B2(n8896), .ZN(
        n4872) );
  INV_X1 U5489 ( .A(n4873), .ZN(n13085) );
  AOI22_X1 U5490 ( .A1(ram[466]), .A2(n4871), .B1(n13099), .B2(n8920), .ZN(
        n4873) );
  INV_X1 U5491 ( .A(n4874), .ZN(n13086) );
  AOI22_X1 U5492 ( .A1(ram[467]), .A2(n4871), .B1(n13099), .B2(n8944), .ZN(
        n4874) );
  INV_X1 U5493 ( .A(n4875), .ZN(n13087) );
  AOI22_X1 U5494 ( .A1(ram[468]), .A2(n4871), .B1(n13099), .B2(n8968), .ZN(
        n4875) );
  INV_X1 U5495 ( .A(n4876), .ZN(n13088) );
  AOI22_X1 U5496 ( .A1(ram[469]), .A2(n4871), .B1(n13099), .B2(n8992), .ZN(
        n4876) );
  INV_X1 U5497 ( .A(n4877), .ZN(n13089) );
  AOI22_X1 U5498 ( .A1(ram[470]), .A2(n4871), .B1(n13099), .B2(n9016), .ZN(
        n4877) );
  INV_X1 U5499 ( .A(n4878), .ZN(n13090) );
  AOI22_X1 U5500 ( .A1(ram[471]), .A2(n4871), .B1(n13099), .B2(n9040), .ZN(
        n4878) );
  INV_X1 U5501 ( .A(n4879), .ZN(n13091) );
  AOI22_X1 U5502 ( .A1(ram[472]), .A2(n4871), .B1(n13099), .B2(n9064), .ZN(
        n4879) );
  INV_X1 U5503 ( .A(n4880), .ZN(n13092) );
  AOI22_X1 U5504 ( .A1(ram[473]), .A2(n4871), .B1(n13099), .B2(n9088), .ZN(
        n4880) );
  INV_X1 U5505 ( .A(n4881), .ZN(n13093) );
  AOI22_X1 U5506 ( .A1(ram[474]), .A2(n4871), .B1(n13099), .B2(n9112), .ZN(
        n4881) );
  INV_X1 U5507 ( .A(n4882), .ZN(n13094) );
  AOI22_X1 U5508 ( .A1(ram[475]), .A2(n4871), .B1(n13099), .B2(n9136), .ZN(
        n4882) );
  INV_X1 U5509 ( .A(n4883), .ZN(n13095) );
  AOI22_X1 U5510 ( .A1(ram[476]), .A2(n4871), .B1(n13099), .B2(n9160), .ZN(
        n4883) );
  INV_X1 U5511 ( .A(n4884), .ZN(n13096) );
  AOI22_X1 U5512 ( .A1(ram[477]), .A2(n4871), .B1(n13099), .B2(n9184), .ZN(
        n4884) );
  INV_X1 U5513 ( .A(n4885), .ZN(n13097) );
  AOI22_X1 U5514 ( .A1(ram[478]), .A2(n4871), .B1(n13099), .B2(n9208), .ZN(
        n4885) );
  INV_X1 U5515 ( .A(n4886), .ZN(n13098) );
  AOI22_X1 U5516 ( .A1(ram[479]), .A2(n4871), .B1(n13099), .B2(n9232), .ZN(
        n4886) );
  INV_X1 U5517 ( .A(n4904), .ZN(n13049) );
  AOI22_X1 U5518 ( .A1(ram[496]), .A2(n4905), .B1(n13065), .B2(n8872), .ZN(
        n4904) );
  INV_X1 U5519 ( .A(n4906), .ZN(n13050) );
  AOI22_X1 U5520 ( .A1(ram[497]), .A2(n4905), .B1(n13065), .B2(n8896), .ZN(
        n4906) );
  INV_X1 U5521 ( .A(n4907), .ZN(n13051) );
  AOI22_X1 U5522 ( .A1(ram[498]), .A2(n4905), .B1(n13065), .B2(n8920), .ZN(
        n4907) );
  INV_X1 U5523 ( .A(n4908), .ZN(n13052) );
  AOI22_X1 U5524 ( .A1(ram[499]), .A2(n4905), .B1(n13065), .B2(n8944), .ZN(
        n4908) );
  INV_X1 U5525 ( .A(n4909), .ZN(n13053) );
  AOI22_X1 U5526 ( .A1(ram[500]), .A2(n4905), .B1(n13065), .B2(n8968), .ZN(
        n4909) );
  INV_X1 U5527 ( .A(n4910), .ZN(n13054) );
  AOI22_X1 U5528 ( .A1(ram[501]), .A2(n4905), .B1(n13065), .B2(n8992), .ZN(
        n4910) );
  INV_X1 U5529 ( .A(n4911), .ZN(n13055) );
  AOI22_X1 U5530 ( .A1(ram[502]), .A2(n4905), .B1(n13065), .B2(n9016), .ZN(
        n4911) );
  INV_X1 U5531 ( .A(n4912), .ZN(n13056) );
  AOI22_X1 U5532 ( .A1(ram[503]), .A2(n4905), .B1(n13065), .B2(n9040), .ZN(
        n4912) );
  INV_X1 U5533 ( .A(n4913), .ZN(n13057) );
  AOI22_X1 U5534 ( .A1(ram[504]), .A2(n4905), .B1(n13065), .B2(n9064), .ZN(
        n4913) );
  INV_X1 U5535 ( .A(n4914), .ZN(n13058) );
  AOI22_X1 U5536 ( .A1(ram[505]), .A2(n4905), .B1(n13065), .B2(n9088), .ZN(
        n4914) );
  INV_X1 U5537 ( .A(n4915), .ZN(n13059) );
  AOI22_X1 U5538 ( .A1(ram[506]), .A2(n4905), .B1(n13065), .B2(n9112), .ZN(
        n4915) );
  INV_X1 U5539 ( .A(n4916), .ZN(n13060) );
  AOI22_X1 U5540 ( .A1(ram[507]), .A2(n4905), .B1(n13065), .B2(n9136), .ZN(
        n4916) );
  INV_X1 U5541 ( .A(n4917), .ZN(n13061) );
  AOI22_X1 U5542 ( .A1(ram[508]), .A2(n4905), .B1(n13065), .B2(n9160), .ZN(
        n4917) );
  INV_X1 U5543 ( .A(n4918), .ZN(n13062) );
  AOI22_X1 U5544 ( .A1(ram[509]), .A2(n4905), .B1(n13065), .B2(n9184), .ZN(
        n4918) );
  INV_X1 U5545 ( .A(n4919), .ZN(n13063) );
  AOI22_X1 U5546 ( .A1(ram[510]), .A2(n4905), .B1(n13065), .B2(n9208), .ZN(
        n4919) );
  INV_X1 U5547 ( .A(n4920), .ZN(n13064) );
  AOI22_X1 U5548 ( .A1(ram[511]), .A2(n4905), .B1(n13065), .B2(n9232), .ZN(
        n4920) );
  INV_X1 U5549 ( .A(n4940), .ZN(n13015) );
  AOI22_X1 U5550 ( .A1(ram[528]), .A2(n4941), .B1(n13031), .B2(n8872), .ZN(
        n4940) );
  INV_X1 U5551 ( .A(n4942), .ZN(n13016) );
  AOI22_X1 U5552 ( .A1(ram[529]), .A2(n4941), .B1(n13031), .B2(n8896), .ZN(
        n4942) );
  INV_X1 U5553 ( .A(n4943), .ZN(n13017) );
  AOI22_X1 U5554 ( .A1(ram[530]), .A2(n4941), .B1(n13031), .B2(n8920), .ZN(
        n4943) );
  INV_X1 U5555 ( .A(n4944), .ZN(n13018) );
  AOI22_X1 U5556 ( .A1(ram[531]), .A2(n4941), .B1(n13031), .B2(n8944), .ZN(
        n4944) );
  INV_X1 U5557 ( .A(n4945), .ZN(n13019) );
  AOI22_X1 U5558 ( .A1(ram[532]), .A2(n4941), .B1(n13031), .B2(n8968), .ZN(
        n4945) );
  INV_X1 U5559 ( .A(n4946), .ZN(n13020) );
  AOI22_X1 U5560 ( .A1(ram[533]), .A2(n4941), .B1(n13031), .B2(n8992), .ZN(
        n4946) );
  INV_X1 U5561 ( .A(n4947), .ZN(n13021) );
  AOI22_X1 U5562 ( .A1(ram[534]), .A2(n4941), .B1(n13031), .B2(n9016), .ZN(
        n4947) );
  INV_X1 U5563 ( .A(n4948), .ZN(n13022) );
  AOI22_X1 U5564 ( .A1(ram[535]), .A2(n4941), .B1(n13031), .B2(n9040), .ZN(
        n4948) );
  INV_X1 U5565 ( .A(n4949), .ZN(n13023) );
  AOI22_X1 U5566 ( .A1(ram[536]), .A2(n4941), .B1(n13031), .B2(n9064), .ZN(
        n4949) );
  INV_X1 U5567 ( .A(n4950), .ZN(n13024) );
  AOI22_X1 U5568 ( .A1(ram[537]), .A2(n4941), .B1(n13031), .B2(n9088), .ZN(
        n4950) );
  INV_X1 U5569 ( .A(n4951), .ZN(n13025) );
  AOI22_X1 U5570 ( .A1(ram[538]), .A2(n4941), .B1(n13031), .B2(n9112), .ZN(
        n4951) );
  INV_X1 U5571 ( .A(n4952), .ZN(n13026) );
  AOI22_X1 U5572 ( .A1(ram[539]), .A2(n4941), .B1(n13031), .B2(n9136), .ZN(
        n4952) );
  INV_X1 U5573 ( .A(n4953), .ZN(n13027) );
  AOI22_X1 U5574 ( .A1(ram[540]), .A2(n4941), .B1(n13031), .B2(n9160), .ZN(
        n4953) );
  INV_X1 U5575 ( .A(n4954), .ZN(n13028) );
  AOI22_X1 U5576 ( .A1(ram[541]), .A2(n4941), .B1(n13031), .B2(n9184), .ZN(
        n4954) );
  INV_X1 U5577 ( .A(n4955), .ZN(n13029) );
  AOI22_X1 U5578 ( .A1(ram[542]), .A2(n4941), .B1(n13031), .B2(n9208), .ZN(
        n4955) );
  INV_X1 U5579 ( .A(n4956), .ZN(n13030) );
  AOI22_X1 U5580 ( .A1(ram[543]), .A2(n4941), .B1(n13031), .B2(n9232), .ZN(
        n4956) );
  INV_X1 U5581 ( .A(n4974), .ZN(n12981) );
  AOI22_X1 U5582 ( .A1(ram[560]), .A2(n4975), .B1(n12997), .B2(n8872), .ZN(
        n4974) );
  INV_X1 U5583 ( .A(n4976), .ZN(n12982) );
  AOI22_X1 U5584 ( .A1(ram[561]), .A2(n4975), .B1(n12997), .B2(n8896), .ZN(
        n4976) );
  INV_X1 U5585 ( .A(n4977), .ZN(n12983) );
  AOI22_X1 U5586 ( .A1(ram[562]), .A2(n4975), .B1(n12997), .B2(n8920), .ZN(
        n4977) );
  INV_X1 U5587 ( .A(n4978), .ZN(n12984) );
  AOI22_X1 U5588 ( .A1(ram[563]), .A2(n4975), .B1(n12997), .B2(n8944), .ZN(
        n4978) );
  INV_X1 U5589 ( .A(n4979), .ZN(n12985) );
  AOI22_X1 U5590 ( .A1(ram[564]), .A2(n4975), .B1(n12997), .B2(n8968), .ZN(
        n4979) );
  INV_X1 U5591 ( .A(n4980), .ZN(n12986) );
  AOI22_X1 U5592 ( .A1(ram[565]), .A2(n4975), .B1(n12997), .B2(n8992), .ZN(
        n4980) );
  INV_X1 U5593 ( .A(n4981), .ZN(n12987) );
  AOI22_X1 U5594 ( .A1(ram[566]), .A2(n4975), .B1(n12997), .B2(n9016), .ZN(
        n4981) );
  INV_X1 U5595 ( .A(n4982), .ZN(n12988) );
  AOI22_X1 U5596 ( .A1(ram[567]), .A2(n4975), .B1(n12997), .B2(n9040), .ZN(
        n4982) );
  INV_X1 U5597 ( .A(n4983), .ZN(n12989) );
  AOI22_X1 U5598 ( .A1(ram[568]), .A2(n4975), .B1(n12997), .B2(n9064), .ZN(
        n4983) );
  INV_X1 U5599 ( .A(n4984), .ZN(n12990) );
  AOI22_X1 U5600 ( .A1(ram[569]), .A2(n4975), .B1(n12997), .B2(n9088), .ZN(
        n4984) );
  INV_X1 U5601 ( .A(n4985), .ZN(n12991) );
  AOI22_X1 U5602 ( .A1(ram[570]), .A2(n4975), .B1(n12997), .B2(n9112), .ZN(
        n4985) );
  INV_X1 U5603 ( .A(n4986), .ZN(n12992) );
  AOI22_X1 U5604 ( .A1(ram[571]), .A2(n4975), .B1(n12997), .B2(n9136), .ZN(
        n4986) );
  INV_X1 U5605 ( .A(n4987), .ZN(n12993) );
  AOI22_X1 U5606 ( .A1(ram[572]), .A2(n4975), .B1(n12997), .B2(n9160), .ZN(
        n4987) );
  INV_X1 U5607 ( .A(n4988), .ZN(n12994) );
  AOI22_X1 U5608 ( .A1(ram[573]), .A2(n4975), .B1(n12997), .B2(n9184), .ZN(
        n4988) );
  INV_X1 U5609 ( .A(n4989), .ZN(n12995) );
  AOI22_X1 U5610 ( .A1(ram[574]), .A2(n4975), .B1(n12997), .B2(n9208), .ZN(
        n4989) );
  INV_X1 U5611 ( .A(n4990), .ZN(n12996) );
  AOI22_X1 U5612 ( .A1(ram[575]), .A2(n4975), .B1(n12997), .B2(n9232), .ZN(
        n4990) );
  INV_X1 U5613 ( .A(n5008), .ZN(n12947) );
  AOI22_X1 U5614 ( .A1(ram[592]), .A2(n5009), .B1(n12963), .B2(n8872), .ZN(
        n5008) );
  INV_X1 U5615 ( .A(n5010), .ZN(n12948) );
  AOI22_X1 U5616 ( .A1(ram[593]), .A2(n5009), .B1(n12963), .B2(n8896), .ZN(
        n5010) );
  INV_X1 U5617 ( .A(n5011), .ZN(n12949) );
  AOI22_X1 U5618 ( .A1(ram[594]), .A2(n5009), .B1(n12963), .B2(n8920), .ZN(
        n5011) );
  INV_X1 U5619 ( .A(n5012), .ZN(n12950) );
  AOI22_X1 U5620 ( .A1(ram[595]), .A2(n5009), .B1(n12963), .B2(n8944), .ZN(
        n5012) );
  INV_X1 U5621 ( .A(n5013), .ZN(n12951) );
  AOI22_X1 U5622 ( .A1(ram[596]), .A2(n5009), .B1(n12963), .B2(n8968), .ZN(
        n5013) );
  INV_X1 U5623 ( .A(n5014), .ZN(n12952) );
  AOI22_X1 U5624 ( .A1(ram[597]), .A2(n5009), .B1(n12963), .B2(n8992), .ZN(
        n5014) );
  INV_X1 U5625 ( .A(n5015), .ZN(n12953) );
  AOI22_X1 U5626 ( .A1(ram[598]), .A2(n5009), .B1(n12963), .B2(n9016), .ZN(
        n5015) );
  INV_X1 U5627 ( .A(n5016), .ZN(n12954) );
  AOI22_X1 U5628 ( .A1(ram[599]), .A2(n5009), .B1(n12963), .B2(n9040), .ZN(
        n5016) );
  INV_X1 U5629 ( .A(n5017), .ZN(n12955) );
  AOI22_X1 U5630 ( .A1(ram[600]), .A2(n5009), .B1(n12963), .B2(n9064), .ZN(
        n5017) );
  INV_X1 U5631 ( .A(n5018), .ZN(n12956) );
  AOI22_X1 U5632 ( .A1(ram[601]), .A2(n5009), .B1(n12963), .B2(n9088), .ZN(
        n5018) );
  INV_X1 U5633 ( .A(n5019), .ZN(n12957) );
  AOI22_X1 U5634 ( .A1(ram[602]), .A2(n5009), .B1(n12963), .B2(n9112), .ZN(
        n5019) );
  INV_X1 U5635 ( .A(n5020), .ZN(n12958) );
  AOI22_X1 U5636 ( .A1(ram[603]), .A2(n5009), .B1(n12963), .B2(n9136), .ZN(
        n5020) );
  INV_X1 U5637 ( .A(n5021), .ZN(n12959) );
  AOI22_X1 U5638 ( .A1(ram[604]), .A2(n5009), .B1(n12963), .B2(n9160), .ZN(
        n5021) );
  INV_X1 U5639 ( .A(n5022), .ZN(n12960) );
  AOI22_X1 U5640 ( .A1(ram[605]), .A2(n5009), .B1(n12963), .B2(n9184), .ZN(
        n5022) );
  INV_X1 U5641 ( .A(n5023), .ZN(n12961) );
  AOI22_X1 U5642 ( .A1(ram[606]), .A2(n5009), .B1(n12963), .B2(n9208), .ZN(
        n5023) );
  INV_X1 U5643 ( .A(n5024), .ZN(n12962) );
  AOI22_X1 U5644 ( .A1(ram[607]), .A2(n5009), .B1(n12963), .B2(n9232), .ZN(
        n5024) );
  INV_X1 U5645 ( .A(n5042), .ZN(n12913) );
  AOI22_X1 U5646 ( .A1(ram[624]), .A2(n5043), .B1(n12929), .B2(n8872), .ZN(
        n5042) );
  INV_X1 U5647 ( .A(n5044), .ZN(n12914) );
  AOI22_X1 U5648 ( .A1(ram[625]), .A2(n5043), .B1(n12929), .B2(n8896), .ZN(
        n5044) );
  INV_X1 U5649 ( .A(n5045), .ZN(n12915) );
  AOI22_X1 U5650 ( .A1(ram[626]), .A2(n5043), .B1(n12929), .B2(n8920), .ZN(
        n5045) );
  INV_X1 U5651 ( .A(n5046), .ZN(n12916) );
  AOI22_X1 U5652 ( .A1(ram[627]), .A2(n5043), .B1(n12929), .B2(n8944), .ZN(
        n5046) );
  INV_X1 U5653 ( .A(n5047), .ZN(n12917) );
  AOI22_X1 U5654 ( .A1(ram[628]), .A2(n5043), .B1(n12929), .B2(n8968), .ZN(
        n5047) );
  INV_X1 U5655 ( .A(n5048), .ZN(n12918) );
  AOI22_X1 U5656 ( .A1(ram[629]), .A2(n5043), .B1(n12929), .B2(n8992), .ZN(
        n5048) );
  INV_X1 U5657 ( .A(n5049), .ZN(n12919) );
  AOI22_X1 U5658 ( .A1(ram[630]), .A2(n5043), .B1(n12929), .B2(n9016), .ZN(
        n5049) );
  INV_X1 U5659 ( .A(n5050), .ZN(n12920) );
  AOI22_X1 U5660 ( .A1(ram[631]), .A2(n5043), .B1(n12929), .B2(n9040), .ZN(
        n5050) );
  INV_X1 U5661 ( .A(n5051), .ZN(n12921) );
  AOI22_X1 U5662 ( .A1(ram[632]), .A2(n5043), .B1(n12929), .B2(n9064), .ZN(
        n5051) );
  INV_X1 U5663 ( .A(n5052), .ZN(n12922) );
  AOI22_X1 U5664 ( .A1(ram[633]), .A2(n5043), .B1(n12929), .B2(n9088), .ZN(
        n5052) );
  INV_X1 U5665 ( .A(n5053), .ZN(n12923) );
  AOI22_X1 U5666 ( .A1(ram[634]), .A2(n5043), .B1(n12929), .B2(n9112), .ZN(
        n5053) );
  INV_X1 U5667 ( .A(n5054), .ZN(n12924) );
  AOI22_X1 U5668 ( .A1(ram[635]), .A2(n5043), .B1(n12929), .B2(n9136), .ZN(
        n5054) );
  INV_X1 U5669 ( .A(n5055), .ZN(n12925) );
  AOI22_X1 U5670 ( .A1(ram[636]), .A2(n5043), .B1(n12929), .B2(n9160), .ZN(
        n5055) );
  INV_X1 U5671 ( .A(n5056), .ZN(n12926) );
  AOI22_X1 U5672 ( .A1(ram[637]), .A2(n5043), .B1(n12929), .B2(n9184), .ZN(
        n5056) );
  INV_X1 U5673 ( .A(n5057), .ZN(n12927) );
  AOI22_X1 U5674 ( .A1(ram[638]), .A2(n5043), .B1(n12929), .B2(n9208), .ZN(
        n5057) );
  INV_X1 U5675 ( .A(n5058), .ZN(n12928) );
  AOI22_X1 U5676 ( .A1(ram[639]), .A2(n5043), .B1(n12929), .B2(n9232), .ZN(
        n5058) );
  INV_X1 U5677 ( .A(n5076), .ZN(n12879) );
  AOI22_X1 U5678 ( .A1(ram[656]), .A2(n5077), .B1(n12895), .B2(n8871), .ZN(
        n5076) );
  INV_X1 U5679 ( .A(n5078), .ZN(n12880) );
  AOI22_X1 U5680 ( .A1(ram[657]), .A2(n5077), .B1(n12895), .B2(n8895), .ZN(
        n5078) );
  INV_X1 U5681 ( .A(n5079), .ZN(n12881) );
  AOI22_X1 U5682 ( .A1(ram[658]), .A2(n5077), .B1(n12895), .B2(n8919), .ZN(
        n5079) );
  INV_X1 U5683 ( .A(n5080), .ZN(n12882) );
  AOI22_X1 U5684 ( .A1(ram[659]), .A2(n5077), .B1(n12895), .B2(n8943), .ZN(
        n5080) );
  INV_X1 U5685 ( .A(n5081), .ZN(n12883) );
  AOI22_X1 U5686 ( .A1(ram[660]), .A2(n5077), .B1(n12895), .B2(n8967), .ZN(
        n5081) );
  INV_X1 U5687 ( .A(n5082), .ZN(n12884) );
  AOI22_X1 U5688 ( .A1(ram[661]), .A2(n5077), .B1(n12895), .B2(n8991), .ZN(
        n5082) );
  INV_X1 U5689 ( .A(n5083), .ZN(n12885) );
  AOI22_X1 U5690 ( .A1(ram[662]), .A2(n5077), .B1(n12895), .B2(n9015), .ZN(
        n5083) );
  INV_X1 U5691 ( .A(n5084), .ZN(n12886) );
  AOI22_X1 U5692 ( .A1(ram[663]), .A2(n5077), .B1(n12895), .B2(n9039), .ZN(
        n5084) );
  INV_X1 U5693 ( .A(n5085), .ZN(n12887) );
  AOI22_X1 U5694 ( .A1(ram[664]), .A2(n5077), .B1(n12895), .B2(n9063), .ZN(
        n5085) );
  INV_X1 U5695 ( .A(n5086), .ZN(n12888) );
  AOI22_X1 U5696 ( .A1(ram[665]), .A2(n5077), .B1(n12895), .B2(n9087), .ZN(
        n5086) );
  INV_X1 U5697 ( .A(n5087), .ZN(n12889) );
  AOI22_X1 U5698 ( .A1(ram[666]), .A2(n5077), .B1(n12895), .B2(n9111), .ZN(
        n5087) );
  INV_X1 U5699 ( .A(n5088), .ZN(n12890) );
  AOI22_X1 U5700 ( .A1(ram[667]), .A2(n5077), .B1(n12895), .B2(n9135), .ZN(
        n5088) );
  INV_X1 U5701 ( .A(n5089), .ZN(n12891) );
  AOI22_X1 U5702 ( .A1(ram[668]), .A2(n5077), .B1(n12895), .B2(n9159), .ZN(
        n5089) );
  INV_X1 U5703 ( .A(n5090), .ZN(n12892) );
  AOI22_X1 U5704 ( .A1(ram[669]), .A2(n5077), .B1(n12895), .B2(n9183), .ZN(
        n5090) );
  INV_X1 U5705 ( .A(n5091), .ZN(n12893) );
  AOI22_X1 U5706 ( .A1(ram[670]), .A2(n5077), .B1(n12895), .B2(n9207), .ZN(
        n5091) );
  INV_X1 U5707 ( .A(n5092), .ZN(n12894) );
  AOI22_X1 U5708 ( .A1(ram[671]), .A2(n5077), .B1(n12895), .B2(n9231), .ZN(
        n5092) );
  INV_X1 U5709 ( .A(n5110), .ZN(n12845) );
  AOI22_X1 U5710 ( .A1(ram[688]), .A2(n5111), .B1(n12861), .B2(n8871), .ZN(
        n5110) );
  INV_X1 U5711 ( .A(n5112), .ZN(n12846) );
  AOI22_X1 U5712 ( .A1(ram[689]), .A2(n5111), .B1(n12861), .B2(n8895), .ZN(
        n5112) );
  INV_X1 U5713 ( .A(n5113), .ZN(n12847) );
  AOI22_X1 U5714 ( .A1(ram[690]), .A2(n5111), .B1(n12861), .B2(n8919), .ZN(
        n5113) );
  INV_X1 U5715 ( .A(n5114), .ZN(n12848) );
  AOI22_X1 U5716 ( .A1(ram[691]), .A2(n5111), .B1(n12861), .B2(n8943), .ZN(
        n5114) );
  INV_X1 U5717 ( .A(n5115), .ZN(n12849) );
  AOI22_X1 U5718 ( .A1(ram[692]), .A2(n5111), .B1(n12861), .B2(n8967), .ZN(
        n5115) );
  INV_X1 U5719 ( .A(n5116), .ZN(n12850) );
  AOI22_X1 U5720 ( .A1(ram[693]), .A2(n5111), .B1(n12861), .B2(n8991), .ZN(
        n5116) );
  INV_X1 U5721 ( .A(n5117), .ZN(n12851) );
  AOI22_X1 U5722 ( .A1(ram[694]), .A2(n5111), .B1(n12861), .B2(n9015), .ZN(
        n5117) );
  INV_X1 U5723 ( .A(n5118), .ZN(n12852) );
  AOI22_X1 U5724 ( .A1(ram[695]), .A2(n5111), .B1(n12861), .B2(n9039), .ZN(
        n5118) );
  INV_X1 U5725 ( .A(n5119), .ZN(n12853) );
  AOI22_X1 U5726 ( .A1(ram[696]), .A2(n5111), .B1(n12861), .B2(n9063), .ZN(
        n5119) );
  INV_X1 U5727 ( .A(n5120), .ZN(n12854) );
  AOI22_X1 U5728 ( .A1(ram[697]), .A2(n5111), .B1(n12861), .B2(n9087), .ZN(
        n5120) );
  INV_X1 U5729 ( .A(n5121), .ZN(n12855) );
  AOI22_X1 U5730 ( .A1(ram[698]), .A2(n5111), .B1(n12861), .B2(n9111), .ZN(
        n5121) );
  INV_X1 U5731 ( .A(n5122), .ZN(n12856) );
  AOI22_X1 U5732 ( .A1(ram[699]), .A2(n5111), .B1(n12861), .B2(n9135), .ZN(
        n5122) );
  INV_X1 U5733 ( .A(n5123), .ZN(n12857) );
  AOI22_X1 U5734 ( .A1(ram[700]), .A2(n5111), .B1(n12861), .B2(n9159), .ZN(
        n5123) );
  INV_X1 U5735 ( .A(n5124), .ZN(n12858) );
  AOI22_X1 U5736 ( .A1(ram[701]), .A2(n5111), .B1(n12861), .B2(n9183), .ZN(
        n5124) );
  INV_X1 U5737 ( .A(n5125), .ZN(n12859) );
  AOI22_X1 U5738 ( .A1(ram[702]), .A2(n5111), .B1(n12861), .B2(n9207), .ZN(
        n5125) );
  INV_X1 U5739 ( .A(n5126), .ZN(n12860) );
  AOI22_X1 U5740 ( .A1(ram[703]), .A2(n5111), .B1(n12861), .B2(n9231), .ZN(
        n5126) );
  INV_X1 U5741 ( .A(n5144), .ZN(n12811) );
  AOI22_X1 U5742 ( .A1(ram[720]), .A2(n5145), .B1(n12827), .B2(n8871), .ZN(
        n5144) );
  INV_X1 U5743 ( .A(n5146), .ZN(n12812) );
  AOI22_X1 U5744 ( .A1(ram[721]), .A2(n5145), .B1(n12827), .B2(n8895), .ZN(
        n5146) );
  INV_X1 U5745 ( .A(n5147), .ZN(n12813) );
  AOI22_X1 U5746 ( .A1(ram[722]), .A2(n5145), .B1(n12827), .B2(n8919), .ZN(
        n5147) );
  INV_X1 U5747 ( .A(n5148), .ZN(n12814) );
  AOI22_X1 U5748 ( .A1(ram[723]), .A2(n5145), .B1(n12827), .B2(n8943), .ZN(
        n5148) );
  INV_X1 U5749 ( .A(n5149), .ZN(n12815) );
  AOI22_X1 U5750 ( .A1(ram[724]), .A2(n5145), .B1(n12827), .B2(n8967), .ZN(
        n5149) );
  INV_X1 U5751 ( .A(n5150), .ZN(n12816) );
  AOI22_X1 U5752 ( .A1(ram[725]), .A2(n5145), .B1(n12827), .B2(n8991), .ZN(
        n5150) );
  INV_X1 U5753 ( .A(n5151), .ZN(n12817) );
  AOI22_X1 U5754 ( .A1(ram[726]), .A2(n5145), .B1(n12827), .B2(n9015), .ZN(
        n5151) );
  INV_X1 U5755 ( .A(n5152), .ZN(n12818) );
  AOI22_X1 U5756 ( .A1(ram[727]), .A2(n5145), .B1(n12827), .B2(n9039), .ZN(
        n5152) );
  INV_X1 U5757 ( .A(n5153), .ZN(n12819) );
  AOI22_X1 U5758 ( .A1(ram[728]), .A2(n5145), .B1(n12827), .B2(n9063), .ZN(
        n5153) );
  INV_X1 U5759 ( .A(n5154), .ZN(n12820) );
  AOI22_X1 U5760 ( .A1(ram[729]), .A2(n5145), .B1(n12827), .B2(n9087), .ZN(
        n5154) );
  INV_X1 U5761 ( .A(n5155), .ZN(n12821) );
  AOI22_X1 U5762 ( .A1(ram[730]), .A2(n5145), .B1(n12827), .B2(n9111), .ZN(
        n5155) );
  INV_X1 U5763 ( .A(n5156), .ZN(n12822) );
  AOI22_X1 U5764 ( .A1(ram[731]), .A2(n5145), .B1(n12827), .B2(n9135), .ZN(
        n5156) );
  INV_X1 U5765 ( .A(n5157), .ZN(n12823) );
  AOI22_X1 U5766 ( .A1(ram[732]), .A2(n5145), .B1(n12827), .B2(n9159), .ZN(
        n5157) );
  INV_X1 U5767 ( .A(n5158), .ZN(n12824) );
  AOI22_X1 U5768 ( .A1(ram[733]), .A2(n5145), .B1(n12827), .B2(n9183), .ZN(
        n5158) );
  INV_X1 U5769 ( .A(n5159), .ZN(n12825) );
  AOI22_X1 U5770 ( .A1(ram[734]), .A2(n5145), .B1(n12827), .B2(n9207), .ZN(
        n5159) );
  INV_X1 U5771 ( .A(n5160), .ZN(n12826) );
  AOI22_X1 U5772 ( .A1(ram[735]), .A2(n5145), .B1(n12827), .B2(n9231), .ZN(
        n5160) );
  INV_X1 U5773 ( .A(n5178), .ZN(n12777) );
  AOI22_X1 U5774 ( .A1(ram[752]), .A2(n5179), .B1(n12793), .B2(n8871), .ZN(
        n5178) );
  INV_X1 U5775 ( .A(n5180), .ZN(n12778) );
  AOI22_X1 U5776 ( .A1(ram[753]), .A2(n5179), .B1(n12793), .B2(n8895), .ZN(
        n5180) );
  INV_X1 U5777 ( .A(n5181), .ZN(n12779) );
  AOI22_X1 U5778 ( .A1(ram[754]), .A2(n5179), .B1(n12793), .B2(n8919), .ZN(
        n5181) );
  INV_X1 U5779 ( .A(n5182), .ZN(n12780) );
  AOI22_X1 U5780 ( .A1(ram[755]), .A2(n5179), .B1(n12793), .B2(n8943), .ZN(
        n5182) );
  INV_X1 U5781 ( .A(n5183), .ZN(n12781) );
  AOI22_X1 U5782 ( .A1(ram[756]), .A2(n5179), .B1(n12793), .B2(n8967), .ZN(
        n5183) );
  INV_X1 U5783 ( .A(n5184), .ZN(n12782) );
  AOI22_X1 U5784 ( .A1(ram[757]), .A2(n5179), .B1(n12793), .B2(n8991), .ZN(
        n5184) );
  INV_X1 U5785 ( .A(n5185), .ZN(n12783) );
  AOI22_X1 U5786 ( .A1(ram[758]), .A2(n5179), .B1(n12793), .B2(n9015), .ZN(
        n5185) );
  INV_X1 U5787 ( .A(n5186), .ZN(n12784) );
  AOI22_X1 U5788 ( .A1(ram[759]), .A2(n5179), .B1(n12793), .B2(n9039), .ZN(
        n5186) );
  INV_X1 U5789 ( .A(n5187), .ZN(n12785) );
  AOI22_X1 U5790 ( .A1(ram[760]), .A2(n5179), .B1(n12793), .B2(n9063), .ZN(
        n5187) );
  INV_X1 U5791 ( .A(n5188), .ZN(n12786) );
  AOI22_X1 U5792 ( .A1(ram[761]), .A2(n5179), .B1(n12793), .B2(n9087), .ZN(
        n5188) );
  INV_X1 U5793 ( .A(n5189), .ZN(n12787) );
  AOI22_X1 U5794 ( .A1(ram[762]), .A2(n5179), .B1(n12793), .B2(n9111), .ZN(
        n5189) );
  INV_X1 U5795 ( .A(n5190), .ZN(n12788) );
  AOI22_X1 U5796 ( .A1(ram[763]), .A2(n5179), .B1(n12793), .B2(n9135), .ZN(
        n5190) );
  INV_X1 U5797 ( .A(n5191), .ZN(n12789) );
  AOI22_X1 U5798 ( .A1(ram[764]), .A2(n5179), .B1(n12793), .B2(n9159), .ZN(
        n5191) );
  INV_X1 U5799 ( .A(n5192), .ZN(n12790) );
  AOI22_X1 U5800 ( .A1(ram[765]), .A2(n5179), .B1(n12793), .B2(n9183), .ZN(
        n5192) );
  INV_X1 U5801 ( .A(n5193), .ZN(n12791) );
  AOI22_X1 U5802 ( .A1(ram[766]), .A2(n5179), .B1(n12793), .B2(n9207), .ZN(
        n5193) );
  INV_X1 U5803 ( .A(n5194), .ZN(n12792) );
  AOI22_X1 U5804 ( .A1(ram[767]), .A2(n5179), .B1(n12793), .B2(n9231), .ZN(
        n5194) );
  INV_X1 U5805 ( .A(n5214), .ZN(n12743) );
  AOI22_X1 U5806 ( .A1(ram[784]), .A2(n5215), .B1(n12759), .B2(n8871), .ZN(
        n5214) );
  INV_X1 U5807 ( .A(n5216), .ZN(n12744) );
  AOI22_X1 U5808 ( .A1(ram[785]), .A2(n5215), .B1(n12759), .B2(n8895), .ZN(
        n5216) );
  INV_X1 U5809 ( .A(n5217), .ZN(n12745) );
  AOI22_X1 U5810 ( .A1(ram[786]), .A2(n5215), .B1(n12759), .B2(n8919), .ZN(
        n5217) );
  INV_X1 U5811 ( .A(n5218), .ZN(n12746) );
  AOI22_X1 U5812 ( .A1(ram[787]), .A2(n5215), .B1(n12759), .B2(n8943), .ZN(
        n5218) );
  INV_X1 U5813 ( .A(n5219), .ZN(n12747) );
  AOI22_X1 U5814 ( .A1(ram[788]), .A2(n5215), .B1(n12759), .B2(n8967), .ZN(
        n5219) );
  INV_X1 U5815 ( .A(n5220), .ZN(n12748) );
  AOI22_X1 U5816 ( .A1(ram[789]), .A2(n5215), .B1(n12759), .B2(n8991), .ZN(
        n5220) );
  INV_X1 U5817 ( .A(n5221), .ZN(n12749) );
  AOI22_X1 U5818 ( .A1(ram[790]), .A2(n5215), .B1(n12759), .B2(n9015), .ZN(
        n5221) );
  INV_X1 U5819 ( .A(n5222), .ZN(n12750) );
  AOI22_X1 U5820 ( .A1(ram[791]), .A2(n5215), .B1(n12759), .B2(n9039), .ZN(
        n5222) );
  INV_X1 U5821 ( .A(n5223), .ZN(n12751) );
  AOI22_X1 U5822 ( .A1(ram[792]), .A2(n5215), .B1(n12759), .B2(n9063), .ZN(
        n5223) );
  INV_X1 U5823 ( .A(n5224), .ZN(n12752) );
  AOI22_X1 U5824 ( .A1(ram[793]), .A2(n5215), .B1(n12759), .B2(n9087), .ZN(
        n5224) );
  INV_X1 U5825 ( .A(n5225), .ZN(n12753) );
  AOI22_X1 U5826 ( .A1(ram[794]), .A2(n5215), .B1(n12759), .B2(n9111), .ZN(
        n5225) );
  INV_X1 U5827 ( .A(n5226), .ZN(n12754) );
  AOI22_X1 U5828 ( .A1(ram[795]), .A2(n5215), .B1(n12759), .B2(n9135), .ZN(
        n5226) );
  INV_X1 U5829 ( .A(n5227), .ZN(n12755) );
  AOI22_X1 U5830 ( .A1(ram[796]), .A2(n5215), .B1(n12759), .B2(n9159), .ZN(
        n5227) );
  INV_X1 U5831 ( .A(n5228), .ZN(n12756) );
  AOI22_X1 U5832 ( .A1(ram[797]), .A2(n5215), .B1(n12759), .B2(n9183), .ZN(
        n5228) );
  INV_X1 U5833 ( .A(n5229), .ZN(n12757) );
  AOI22_X1 U5834 ( .A1(ram[798]), .A2(n5215), .B1(n12759), .B2(n9207), .ZN(
        n5229) );
  INV_X1 U5835 ( .A(n5230), .ZN(n12758) );
  AOI22_X1 U5836 ( .A1(ram[799]), .A2(n5215), .B1(n12759), .B2(n9231), .ZN(
        n5230) );
  INV_X1 U5837 ( .A(n5248), .ZN(n12709) );
  AOI22_X1 U5838 ( .A1(ram[816]), .A2(n5249), .B1(n12725), .B2(n8871), .ZN(
        n5248) );
  INV_X1 U5839 ( .A(n5250), .ZN(n12710) );
  AOI22_X1 U5840 ( .A1(ram[817]), .A2(n5249), .B1(n12725), .B2(n8895), .ZN(
        n5250) );
  INV_X1 U5841 ( .A(n5251), .ZN(n12711) );
  AOI22_X1 U5842 ( .A1(ram[818]), .A2(n5249), .B1(n12725), .B2(n8919), .ZN(
        n5251) );
  INV_X1 U5843 ( .A(n5252), .ZN(n12712) );
  AOI22_X1 U5844 ( .A1(ram[819]), .A2(n5249), .B1(n12725), .B2(n8943), .ZN(
        n5252) );
  INV_X1 U5845 ( .A(n5253), .ZN(n12713) );
  AOI22_X1 U5846 ( .A1(ram[820]), .A2(n5249), .B1(n12725), .B2(n8967), .ZN(
        n5253) );
  INV_X1 U5847 ( .A(n5254), .ZN(n12714) );
  AOI22_X1 U5848 ( .A1(ram[821]), .A2(n5249), .B1(n12725), .B2(n8991), .ZN(
        n5254) );
  INV_X1 U5849 ( .A(n5255), .ZN(n12715) );
  AOI22_X1 U5850 ( .A1(ram[822]), .A2(n5249), .B1(n12725), .B2(n9015), .ZN(
        n5255) );
  INV_X1 U5851 ( .A(n5256), .ZN(n12716) );
  AOI22_X1 U5852 ( .A1(ram[823]), .A2(n5249), .B1(n12725), .B2(n9039), .ZN(
        n5256) );
  INV_X1 U5853 ( .A(n5257), .ZN(n12717) );
  AOI22_X1 U5854 ( .A1(ram[824]), .A2(n5249), .B1(n12725), .B2(n9063), .ZN(
        n5257) );
  INV_X1 U5855 ( .A(n5258), .ZN(n12718) );
  AOI22_X1 U5856 ( .A1(ram[825]), .A2(n5249), .B1(n12725), .B2(n9087), .ZN(
        n5258) );
  INV_X1 U5857 ( .A(n5259), .ZN(n12719) );
  AOI22_X1 U5858 ( .A1(ram[826]), .A2(n5249), .B1(n12725), .B2(n9111), .ZN(
        n5259) );
  INV_X1 U5859 ( .A(n5260), .ZN(n12720) );
  AOI22_X1 U5860 ( .A1(ram[827]), .A2(n5249), .B1(n12725), .B2(n9135), .ZN(
        n5260) );
  INV_X1 U5861 ( .A(n5261), .ZN(n12721) );
  AOI22_X1 U5862 ( .A1(ram[828]), .A2(n5249), .B1(n12725), .B2(n9159), .ZN(
        n5261) );
  INV_X1 U5863 ( .A(n5262), .ZN(n12722) );
  AOI22_X1 U5864 ( .A1(ram[829]), .A2(n5249), .B1(n12725), .B2(n9183), .ZN(
        n5262) );
  INV_X1 U5865 ( .A(n5263), .ZN(n12723) );
  AOI22_X1 U5866 ( .A1(ram[830]), .A2(n5249), .B1(n12725), .B2(n9207), .ZN(
        n5263) );
  INV_X1 U5867 ( .A(n5264), .ZN(n12724) );
  AOI22_X1 U5868 ( .A1(ram[831]), .A2(n5249), .B1(n12725), .B2(n9231), .ZN(
        n5264) );
  INV_X1 U5869 ( .A(n5282), .ZN(n12675) );
  AOI22_X1 U5870 ( .A1(ram[848]), .A2(n5283), .B1(n12691), .B2(n8870), .ZN(
        n5282) );
  INV_X1 U5871 ( .A(n5284), .ZN(n12676) );
  AOI22_X1 U5872 ( .A1(ram[849]), .A2(n5283), .B1(n12691), .B2(n8894), .ZN(
        n5284) );
  INV_X1 U5873 ( .A(n5285), .ZN(n12677) );
  AOI22_X1 U5874 ( .A1(ram[850]), .A2(n5283), .B1(n12691), .B2(n8918), .ZN(
        n5285) );
  INV_X1 U5875 ( .A(n5286), .ZN(n12678) );
  AOI22_X1 U5876 ( .A1(ram[851]), .A2(n5283), .B1(n12691), .B2(n8942), .ZN(
        n5286) );
  INV_X1 U5877 ( .A(n5287), .ZN(n12679) );
  AOI22_X1 U5878 ( .A1(ram[852]), .A2(n5283), .B1(n12691), .B2(n8966), .ZN(
        n5287) );
  INV_X1 U5879 ( .A(n5288), .ZN(n12680) );
  AOI22_X1 U5880 ( .A1(ram[853]), .A2(n5283), .B1(n12691), .B2(n8990), .ZN(
        n5288) );
  INV_X1 U5881 ( .A(n5289), .ZN(n12681) );
  AOI22_X1 U5882 ( .A1(ram[854]), .A2(n5283), .B1(n12691), .B2(n9014), .ZN(
        n5289) );
  INV_X1 U5883 ( .A(n5290), .ZN(n12682) );
  AOI22_X1 U5884 ( .A1(ram[855]), .A2(n5283), .B1(n12691), .B2(n9038), .ZN(
        n5290) );
  INV_X1 U5885 ( .A(n5291), .ZN(n12683) );
  AOI22_X1 U5886 ( .A1(ram[856]), .A2(n5283), .B1(n12691), .B2(n9062), .ZN(
        n5291) );
  INV_X1 U5887 ( .A(n5292), .ZN(n12684) );
  AOI22_X1 U5888 ( .A1(ram[857]), .A2(n5283), .B1(n12691), .B2(n9086), .ZN(
        n5292) );
  INV_X1 U5889 ( .A(n5293), .ZN(n12685) );
  AOI22_X1 U5890 ( .A1(ram[858]), .A2(n5283), .B1(n12691), .B2(n9110), .ZN(
        n5293) );
  INV_X1 U5891 ( .A(n5294), .ZN(n12686) );
  AOI22_X1 U5892 ( .A1(ram[859]), .A2(n5283), .B1(n12691), .B2(n9134), .ZN(
        n5294) );
  INV_X1 U5893 ( .A(n5295), .ZN(n12687) );
  AOI22_X1 U5894 ( .A1(ram[860]), .A2(n5283), .B1(n12691), .B2(n9158), .ZN(
        n5295) );
  INV_X1 U5895 ( .A(n5296), .ZN(n12688) );
  AOI22_X1 U5896 ( .A1(ram[861]), .A2(n5283), .B1(n12691), .B2(n9182), .ZN(
        n5296) );
  INV_X1 U5897 ( .A(n5297), .ZN(n12689) );
  AOI22_X1 U5898 ( .A1(ram[862]), .A2(n5283), .B1(n12691), .B2(n9206), .ZN(
        n5297) );
  INV_X1 U5899 ( .A(n5298), .ZN(n12690) );
  AOI22_X1 U5900 ( .A1(ram[863]), .A2(n5283), .B1(n12691), .B2(n9230), .ZN(
        n5298) );
  INV_X1 U5901 ( .A(n5316), .ZN(n12641) );
  AOI22_X1 U5902 ( .A1(ram[880]), .A2(n5317), .B1(n12657), .B2(n8870), .ZN(
        n5316) );
  INV_X1 U5903 ( .A(n5318), .ZN(n12642) );
  AOI22_X1 U5904 ( .A1(ram[881]), .A2(n5317), .B1(n12657), .B2(n8894), .ZN(
        n5318) );
  INV_X1 U5905 ( .A(n5319), .ZN(n12643) );
  AOI22_X1 U5906 ( .A1(ram[882]), .A2(n5317), .B1(n12657), .B2(n8918), .ZN(
        n5319) );
  INV_X1 U5907 ( .A(n5320), .ZN(n12644) );
  AOI22_X1 U5908 ( .A1(ram[883]), .A2(n5317), .B1(n12657), .B2(n8942), .ZN(
        n5320) );
  INV_X1 U5909 ( .A(n5321), .ZN(n12645) );
  AOI22_X1 U5910 ( .A1(ram[884]), .A2(n5317), .B1(n12657), .B2(n8966), .ZN(
        n5321) );
  INV_X1 U5911 ( .A(n5322), .ZN(n12646) );
  AOI22_X1 U5912 ( .A1(ram[885]), .A2(n5317), .B1(n12657), .B2(n8990), .ZN(
        n5322) );
  INV_X1 U5913 ( .A(n5323), .ZN(n12647) );
  AOI22_X1 U5914 ( .A1(ram[886]), .A2(n5317), .B1(n12657), .B2(n9014), .ZN(
        n5323) );
  INV_X1 U5915 ( .A(n5324), .ZN(n12648) );
  AOI22_X1 U5916 ( .A1(ram[887]), .A2(n5317), .B1(n12657), .B2(n9038), .ZN(
        n5324) );
  INV_X1 U5917 ( .A(n5325), .ZN(n12649) );
  AOI22_X1 U5918 ( .A1(ram[888]), .A2(n5317), .B1(n12657), .B2(n9062), .ZN(
        n5325) );
  INV_X1 U5919 ( .A(n5326), .ZN(n12650) );
  AOI22_X1 U5920 ( .A1(ram[889]), .A2(n5317), .B1(n12657), .B2(n9086), .ZN(
        n5326) );
  INV_X1 U5921 ( .A(n5327), .ZN(n12651) );
  AOI22_X1 U5922 ( .A1(ram[890]), .A2(n5317), .B1(n12657), .B2(n9110), .ZN(
        n5327) );
  INV_X1 U5923 ( .A(n5328), .ZN(n12652) );
  AOI22_X1 U5924 ( .A1(ram[891]), .A2(n5317), .B1(n12657), .B2(n9134), .ZN(
        n5328) );
  INV_X1 U5925 ( .A(n5329), .ZN(n12653) );
  AOI22_X1 U5926 ( .A1(ram[892]), .A2(n5317), .B1(n12657), .B2(n9158), .ZN(
        n5329) );
  INV_X1 U5927 ( .A(n5330), .ZN(n12654) );
  AOI22_X1 U5928 ( .A1(ram[893]), .A2(n5317), .B1(n12657), .B2(n9182), .ZN(
        n5330) );
  INV_X1 U5929 ( .A(n5331), .ZN(n12655) );
  AOI22_X1 U5930 ( .A1(ram[894]), .A2(n5317), .B1(n12657), .B2(n9206), .ZN(
        n5331) );
  INV_X1 U5931 ( .A(n5332), .ZN(n12656) );
  AOI22_X1 U5932 ( .A1(ram[895]), .A2(n5317), .B1(n12657), .B2(n9230), .ZN(
        n5332) );
  INV_X1 U5933 ( .A(n5350), .ZN(n12607) );
  AOI22_X1 U5934 ( .A1(ram[912]), .A2(n5351), .B1(n12623), .B2(n8870), .ZN(
        n5350) );
  INV_X1 U5935 ( .A(n5352), .ZN(n12608) );
  AOI22_X1 U5936 ( .A1(ram[913]), .A2(n5351), .B1(n12623), .B2(n8894), .ZN(
        n5352) );
  INV_X1 U5937 ( .A(n5353), .ZN(n12609) );
  AOI22_X1 U5938 ( .A1(ram[914]), .A2(n5351), .B1(n12623), .B2(n8918), .ZN(
        n5353) );
  INV_X1 U5939 ( .A(n5354), .ZN(n12610) );
  AOI22_X1 U5940 ( .A1(ram[915]), .A2(n5351), .B1(n12623), .B2(n8942), .ZN(
        n5354) );
  INV_X1 U5941 ( .A(n5355), .ZN(n12611) );
  AOI22_X1 U5942 ( .A1(ram[916]), .A2(n5351), .B1(n12623), .B2(n8966), .ZN(
        n5355) );
  INV_X1 U5943 ( .A(n5356), .ZN(n12612) );
  AOI22_X1 U5944 ( .A1(ram[917]), .A2(n5351), .B1(n12623), .B2(n8990), .ZN(
        n5356) );
  INV_X1 U5945 ( .A(n5357), .ZN(n12613) );
  AOI22_X1 U5946 ( .A1(ram[918]), .A2(n5351), .B1(n12623), .B2(n9014), .ZN(
        n5357) );
  INV_X1 U5947 ( .A(n5358), .ZN(n12614) );
  AOI22_X1 U5948 ( .A1(ram[919]), .A2(n5351), .B1(n12623), .B2(n9038), .ZN(
        n5358) );
  INV_X1 U5949 ( .A(n5359), .ZN(n12615) );
  AOI22_X1 U5950 ( .A1(ram[920]), .A2(n5351), .B1(n12623), .B2(n9062), .ZN(
        n5359) );
  INV_X1 U5951 ( .A(n5360), .ZN(n12616) );
  AOI22_X1 U5952 ( .A1(ram[921]), .A2(n5351), .B1(n12623), .B2(n9086), .ZN(
        n5360) );
  INV_X1 U5953 ( .A(n5361), .ZN(n12617) );
  AOI22_X1 U5954 ( .A1(ram[922]), .A2(n5351), .B1(n12623), .B2(n9110), .ZN(
        n5361) );
  INV_X1 U5955 ( .A(n5362), .ZN(n12618) );
  AOI22_X1 U5956 ( .A1(ram[923]), .A2(n5351), .B1(n12623), .B2(n9134), .ZN(
        n5362) );
  INV_X1 U5957 ( .A(n5363), .ZN(n12619) );
  AOI22_X1 U5958 ( .A1(ram[924]), .A2(n5351), .B1(n12623), .B2(n9158), .ZN(
        n5363) );
  INV_X1 U5959 ( .A(n5364), .ZN(n12620) );
  AOI22_X1 U5960 ( .A1(ram[925]), .A2(n5351), .B1(n12623), .B2(n9182), .ZN(
        n5364) );
  INV_X1 U5961 ( .A(n5365), .ZN(n12621) );
  AOI22_X1 U5962 ( .A1(ram[926]), .A2(n5351), .B1(n12623), .B2(n9206), .ZN(
        n5365) );
  INV_X1 U5963 ( .A(n5366), .ZN(n12622) );
  AOI22_X1 U5964 ( .A1(ram[927]), .A2(n5351), .B1(n12623), .B2(n9230), .ZN(
        n5366) );
  INV_X1 U5965 ( .A(n5384), .ZN(n12573) );
  AOI22_X1 U5966 ( .A1(ram[944]), .A2(n5385), .B1(n12589), .B2(n8870), .ZN(
        n5384) );
  INV_X1 U5967 ( .A(n5386), .ZN(n12574) );
  AOI22_X1 U5968 ( .A1(ram[945]), .A2(n5385), .B1(n12589), .B2(n8894), .ZN(
        n5386) );
  INV_X1 U5969 ( .A(n5387), .ZN(n12575) );
  AOI22_X1 U5970 ( .A1(ram[946]), .A2(n5385), .B1(n12589), .B2(n8918), .ZN(
        n5387) );
  INV_X1 U5971 ( .A(n5388), .ZN(n12576) );
  AOI22_X1 U5972 ( .A1(ram[947]), .A2(n5385), .B1(n12589), .B2(n8942), .ZN(
        n5388) );
  INV_X1 U5973 ( .A(n5389), .ZN(n12577) );
  AOI22_X1 U5974 ( .A1(ram[948]), .A2(n5385), .B1(n12589), .B2(n8966), .ZN(
        n5389) );
  INV_X1 U5975 ( .A(n5390), .ZN(n12578) );
  AOI22_X1 U5976 ( .A1(ram[949]), .A2(n5385), .B1(n12589), .B2(n8990), .ZN(
        n5390) );
  INV_X1 U5977 ( .A(n5391), .ZN(n12579) );
  AOI22_X1 U5978 ( .A1(ram[950]), .A2(n5385), .B1(n12589), .B2(n9014), .ZN(
        n5391) );
  INV_X1 U5979 ( .A(n5392), .ZN(n12580) );
  AOI22_X1 U5980 ( .A1(ram[951]), .A2(n5385), .B1(n12589), .B2(n9038), .ZN(
        n5392) );
  INV_X1 U5981 ( .A(n5393), .ZN(n12581) );
  AOI22_X1 U5982 ( .A1(ram[952]), .A2(n5385), .B1(n12589), .B2(n9062), .ZN(
        n5393) );
  INV_X1 U5983 ( .A(n5394), .ZN(n12582) );
  AOI22_X1 U5984 ( .A1(ram[953]), .A2(n5385), .B1(n12589), .B2(n9086), .ZN(
        n5394) );
  INV_X1 U5985 ( .A(n5395), .ZN(n12583) );
  AOI22_X1 U5986 ( .A1(ram[954]), .A2(n5385), .B1(n12589), .B2(n9110), .ZN(
        n5395) );
  INV_X1 U5987 ( .A(n5396), .ZN(n12584) );
  AOI22_X1 U5988 ( .A1(ram[955]), .A2(n5385), .B1(n12589), .B2(n9134), .ZN(
        n5396) );
  INV_X1 U5989 ( .A(n5397), .ZN(n12585) );
  AOI22_X1 U5990 ( .A1(ram[956]), .A2(n5385), .B1(n12589), .B2(n9158), .ZN(
        n5397) );
  INV_X1 U5991 ( .A(n5398), .ZN(n12586) );
  AOI22_X1 U5992 ( .A1(ram[957]), .A2(n5385), .B1(n12589), .B2(n9182), .ZN(
        n5398) );
  INV_X1 U5993 ( .A(n5399), .ZN(n12587) );
  AOI22_X1 U5994 ( .A1(ram[958]), .A2(n5385), .B1(n12589), .B2(n9206), .ZN(
        n5399) );
  INV_X1 U5995 ( .A(n5400), .ZN(n12588) );
  AOI22_X1 U5996 ( .A1(ram[959]), .A2(n5385), .B1(n12589), .B2(n9230), .ZN(
        n5400) );
  INV_X1 U5997 ( .A(n5418), .ZN(n12539) );
  AOI22_X1 U5998 ( .A1(ram[976]), .A2(n5419), .B1(n12555), .B2(n8870), .ZN(
        n5418) );
  INV_X1 U5999 ( .A(n5420), .ZN(n12540) );
  AOI22_X1 U6000 ( .A1(ram[977]), .A2(n5419), .B1(n12555), .B2(n8894), .ZN(
        n5420) );
  INV_X1 U6001 ( .A(n5421), .ZN(n12541) );
  AOI22_X1 U6002 ( .A1(ram[978]), .A2(n5419), .B1(n12555), .B2(n8918), .ZN(
        n5421) );
  INV_X1 U6003 ( .A(n5422), .ZN(n12542) );
  AOI22_X1 U6004 ( .A1(ram[979]), .A2(n5419), .B1(n12555), .B2(n8942), .ZN(
        n5422) );
  INV_X1 U6005 ( .A(n5423), .ZN(n12543) );
  AOI22_X1 U6006 ( .A1(ram[980]), .A2(n5419), .B1(n12555), .B2(n8966), .ZN(
        n5423) );
  INV_X1 U6007 ( .A(n5424), .ZN(n12544) );
  AOI22_X1 U6008 ( .A1(ram[981]), .A2(n5419), .B1(n12555), .B2(n8990), .ZN(
        n5424) );
  INV_X1 U6009 ( .A(n5425), .ZN(n12545) );
  AOI22_X1 U6010 ( .A1(ram[982]), .A2(n5419), .B1(n12555), .B2(n9014), .ZN(
        n5425) );
  INV_X1 U6011 ( .A(n5426), .ZN(n12546) );
  AOI22_X1 U6012 ( .A1(ram[983]), .A2(n5419), .B1(n12555), .B2(n9038), .ZN(
        n5426) );
  INV_X1 U6013 ( .A(n5427), .ZN(n12547) );
  AOI22_X1 U6014 ( .A1(ram[984]), .A2(n5419), .B1(n12555), .B2(n9062), .ZN(
        n5427) );
  INV_X1 U6015 ( .A(n5428), .ZN(n12548) );
  AOI22_X1 U6016 ( .A1(ram[985]), .A2(n5419), .B1(n12555), .B2(n9086), .ZN(
        n5428) );
  INV_X1 U6017 ( .A(n5429), .ZN(n12549) );
  AOI22_X1 U6018 ( .A1(ram[986]), .A2(n5419), .B1(n12555), .B2(n9110), .ZN(
        n5429) );
  INV_X1 U6019 ( .A(n5430), .ZN(n12550) );
  AOI22_X1 U6020 ( .A1(ram[987]), .A2(n5419), .B1(n12555), .B2(n9134), .ZN(
        n5430) );
  INV_X1 U6021 ( .A(n5431), .ZN(n12551) );
  AOI22_X1 U6022 ( .A1(ram[988]), .A2(n5419), .B1(n12555), .B2(n9158), .ZN(
        n5431) );
  INV_X1 U6023 ( .A(n5432), .ZN(n12552) );
  AOI22_X1 U6024 ( .A1(ram[989]), .A2(n5419), .B1(n12555), .B2(n9182), .ZN(
        n5432) );
  INV_X1 U6025 ( .A(n5433), .ZN(n12553) );
  AOI22_X1 U6026 ( .A1(ram[990]), .A2(n5419), .B1(n12555), .B2(n9206), .ZN(
        n5433) );
  INV_X1 U6027 ( .A(n5434), .ZN(n12554) );
  AOI22_X1 U6028 ( .A1(ram[991]), .A2(n5419), .B1(n12555), .B2(n9230), .ZN(
        n5434) );
  INV_X1 U6029 ( .A(n5452), .ZN(n12505) );
  AOI22_X1 U6030 ( .A1(ram[1008]), .A2(n5453), .B1(n12521), .B2(n8870), .ZN(
        n5452) );
  INV_X1 U6031 ( .A(n5454), .ZN(n12506) );
  AOI22_X1 U6032 ( .A1(ram[1009]), .A2(n5453), .B1(n12521), .B2(n8894), .ZN(
        n5454) );
  INV_X1 U6033 ( .A(n5455), .ZN(n12507) );
  AOI22_X1 U6034 ( .A1(ram[1010]), .A2(n5453), .B1(n12521), .B2(n8918), .ZN(
        n5455) );
  INV_X1 U6035 ( .A(n5456), .ZN(n12508) );
  AOI22_X1 U6036 ( .A1(ram[1011]), .A2(n5453), .B1(n12521), .B2(n8942), .ZN(
        n5456) );
  INV_X1 U6037 ( .A(n5457), .ZN(n12509) );
  AOI22_X1 U6038 ( .A1(ram[1012]), .A2(n5453), .B1(n12521), .B2(n8966), .ZN(
        n5457) );
  INV_X1 U6039 ( .A(n5458), .ZN(n12510) );
  AOI22_X1 U6040 ( .A1(ram[1013]), .A2(n5453), .B1(n12521), .B2(n8990), .ZN(
        n5458) );
  INV_X1 U6041 ( .A(n5459), .ZN(n12511) );
  AOI22_X1 U6042 ( .A1(ram[1014]), .A2(n5453), .B1(n12521), .B2(n9014), .ZN(
        n5459) );
  INV_X1 U6043 ( .A(n5460), .ZN(n12512) );
  AOI22_X1 U6044 ( .A1(ram[1015]), .A2(n5453), .B1(n12521), .B2(n9038), .ZN(
        n5460) );
  INV_X1 U6045 ( .A(n5461), .ZN(n12513) );
  AOI22_X1 U6046 ( .A1(ram[1016]), .A2(n5453), .B1(n12521), .B2(n9062), .ZN(
        n5461) );
  INV_X1 U6047 ( .A(n5462), .ZN(n12514) );
  AOI22_X1 U6048 ( .A1(ram[1017]), .A2(n5453), .B1(n12521), .B2(n9086), .ZN(
        n5462) );
  INV_X1 U6049 ( .A(n5463), .ZN(n12515) );
  AOI22_X1 U6050 ( .A1(ram[1018]), .A2(n5453), .B1(n12521), .B2(n9110), .ZN(
        n5463) );
  INV_X1 U6051 ( .A(n5464), .ZN(n12516) );
  AOI22_X1 U6052 ( .A1(ram[1019]), .A2(n5453), .B1(n12521), .B2(n9134), .ZN(
        n5464) );
  INV_X1 U6053 ( .A(n5465), .ZN(n12517) );
  AOI22_X1 U6054 ( .A1(ram[1020]), .A2(n5453), .B1(n12521), .B2(n9158), .ZN(
        n5465) );
  INV_X1 U6055 ( .A(n5466), .ZN(n12518) );
  AOI22_X1 U6056 ( .A1(ram[1021]), .A2(n5453), .B1(n12521), .B2(n9182), .ZN(
        n5466) );
  INV_X1 U6057 ( .A(n5467), .ZN(n12519) );
  AOI22_X1 U6058 ( .A1(ram[1022]), .A2(n5453), .B1(n12521), .B2(n9206), .ZN(
        n5467) );
  INV_X1 U6059 ( .A(n5468), .ZN(n12520) );
  AOI22_X1 U6060 ( .A1(ram[1023]), .A2(n5453), .B1(n12521), .B2(n9230), .ZN(
        n5468) );
  INV_X1 U6061 ( .A(n5488), .ZN(n12471) );
  AOI22_X1 U6062 ( .A1(ram[1040]), .A2(n5489), .B1(n12487), .B2(n8869), .ZN(
        n5488) );
  INV_X1 U6063 ( .A(n5490), .ZN(n12472) );
  AOI22_X1 U6064 ( .A1(ram[1041]), .A2(n5489), .B1(n12487), .B2(n8893), .ZN(
        n5490) );
  INV_X1 U6065 ( .A(n5491), .ZN(n12473) );
  AOI22_X1 U6066 ( .A1(ram[1042]), .A2(n5489), .B1(n12487), .B2(n8917), .ZN(
        n5491) );
  INV_X1 U6067 ( .A(n5492), .ZN(n12474) );
  AOI22_X1 U6068 ( .A1(ram[1043]), .A2(n5489), .B1(n12487), .B2(n8941), .ZN(
        n5492) );
  INV_X1 U6069 ( .A(n5493), .ZN(n12475) );
  AOI22_X1 U6070 ( .A1(ram[1044]), .A2(n5489), .B1(n12487), .B2(n8965), .ZN(
        n5493) );
  INV_X1 U6071 ( .A(n5494), .ZN(n12476) );
  AOI22_X1 U6072 ( .A1(ram[1045]), .A2(n5489), .B1(n12487), .B2(n8989), .ZN(
        n5494) );
  INV_X1 U6073 ( .A(n5495), .ZN(n12477) );
  AOI22_X1 U6074 ( .A1(ram[1046]), .A2(n5489), .B1(n12487), .B2(n9013), .ZN(
        n5495) );
  INV_X1 U6075 ( .A(n5496), .ZN(n12478) );
  AOI22_X1 U6076 ( .A1(ram[1047]), .A2(n5489), .B1(n12487), .B2(n9037), .ZN(
        n5496) );
  INV_X1 U6077 ( .A(n5497), .ZN(n12479) );
  AOI22_X1 U6078 ( .A1(ram[1048]), .A2(n5489), .B1(n12487), .B2(n9061), .ZN(
        n5497) );
  INV_X1 U6079 ( .A(n5498), .ZN(n12480) );
  AOI22_X1 U6080 ( .A1(ram[1049]), .A2(n5489), .B1(n12487), .B2(n9085), .ZN(
        n5498) );
  INV_X1 U6081 ( .A(n5499), .ZN(n12481) );
  AOI22_X1 U6082 ( .A1(ram[1050]), .A2(n5489), .B1(n12487), .B2(n9109), .ZN(
        n5499) );
  INV_X1 U6083 ( .A(n5500), .ZN(n12482) );
  AOI22_X1 U6084 ( .A1(ram[1051]), .A2(n5489), .B1(n12487), .B2(n9133), .ZN(
        n5500) );
  INV_X1 U6085 ( .A(n5501), .ZN(n12483) );
  AOI22_X1 U6086 ( .A1(ram[1052]), .A2(n5489), .B1(n12487), .B2(n9157), .ZN(
        n5501) );
  INV_X1 U6087 ( .A(n5502), .ZN(n12484) );
  AOI22_X1 U6088 ( .A1(ram[1053]), .A2(n5489), .B1(n12487), .B2(n9181), .ZN(
        n5502) );
  INV_X1 U6089 ( .A(n5503), .ZN(n12485) );
  AOI22_X1 U6090 ( .A1(ram[1054]), .A2(n5489), .B1(n12487), .B2(n9205), .ZN(
        n5503) );
  INV_X1 U6091 ( .A(n5504), .ZN(n12486) );
  AOI22_X1 U6092 ( .A1(ram[1055]), .A2(n5489), .B1(n12487), .B2(n9229), .ZN(
        n5504) );
  INV_X1 U6093 ( .A(n5522), .ZN(n12437) );
  AOI22_X1 U6094 ( .A1(ram[1072]), .A2(n5523), .B1(n12453), .B2(n8869), .ZN(
        n5522) );
  INV_X1 U6095 ( .A(n5524), .ZN(n12438) );
  AOI22_X1 U6096 ( .A1(ram[1073]), .A2(n5523), .B1(n12453), .B2(n8893), .ZN(
        n5524) );
  INV_X1 U6097 ( .A(n5525), .ZN(n12439) );
  AOI22_X1 U6098 ( .A1(ram[1074]), .A2(n5523), .B1(n12453), .B2(n8917), .ZN(
        n5525) );
  INV_X1 U6099 ( .A(n5526), .ZN(n12440) );
  AOI22_X1 U6100 ( .A1(ram[1075]), .A2(n5523), .B1(n12453), .B2(n8941), .ZN(
        n5526) );
  INV_X1 U6101 ( .A(n5527), .ZN(n12441) );
  AOI22_X1 U6102 ( .A1(ram[1076]), .A2(n5523), .B1(n12453), .B2(n8965), .ZN(
        n5527) );
  INV_X1 U6103 ( .A(n5528), .ZN(n12442) );
  AOI22_X1 U6104 ( .A1(ram[1077]), .A2(n5523), .B1(n12453), .B2(n8989), .ZN(
        n5528) );
  INV_X1 U6105 ( .A(n5529), .ZN(n12443) );
  AOI22_X1 U6106 ( .A1(ram[1078]), .A2(n5523), .B1(n12453), .B2(n9013), .ZN(
        n5529) );
  INV_X1 U6107 ( .A(n5530), .ZN(n12444) );
  AOI22_X1 U6108 ( .A1(ram[1079]), .A2(n5523), .B1(n12453), .B2(n9037), .ZN(
        n5530) );
  INV_X1 U6109 ( .A(n5531), .ZN(n12445) );
  AOI22_X1 U6110 ( .A1(ram[1080]), .A2(n5523), .B1(n12453), .B2(n9061), .ZN(
        n5531) );
  INV_X1 U6111 ( .A(n5532), .ZN(n12446) );
  AOI22_X1 U6112 ( .A1(ram[1081]), .A2(n5523), .B1(n12453), .B2(n9085), .ZN(
        n5532) );
  INV_X1 U6113 ( .A(n5533), .ZN(n12447) );
  AOI22_X1 U6114 ( .A1(ram[1082]), .A2(n5523), .B1(n12453), .B2(n9109), .ZN(
        n5533) );
  INV_X1 U6115 ( .A(n5534), .ZN(n12448) );
  AOI22_X1 U6116 ( .A1(ram[1083]), .A2(n5523), .B1(n12453), .B2(n9133), .ZN(
        n5534) );
  INV_X1 U6117 ( .A(n5535), .ZN(n12449) );
  AOI22_X1 U6118 ( .A1(ram[1084]), .A2(n5523), .B1(n12453), .B2(n9157), .ZN(
        n5535) );
  INV_X1 U6119 ( .A(n5536), .ZN(n12450) );
  AOI22_X1 U6120 ( .A1(ram[1085]), .A2(n5523), .B1(n12453), .B2(n9181), .ZN(
        n5536) );
  INV_X1 U6121 ( .A(n5537), .ZN(n12451) );
  AOI22_X1 U6122 ( .A1(ram[1086]), .A2(n5523), .B1(n12453), .B2(n9205), .ZN(
        n5537) );
  INV_X1 U6123 ( .A(n5538), .ZN(n12452) );
  AOI22_X1 U6124 ( .A1(ram[1087]), .A2(n5523), .B1(n12453), .B2(n9229), .ZN(
        n5538) );
  INV_X1 U6125 ( .A(n5556), .ZN(n12403) );
  AOI22_X1 U6126 ( .A1(ram[1104]), .A2(n5557), .B1(n12419), .B2(n8869), .ZN(
        n5556) );
  INV_X1 U6127 ( .A(n5558), .ZN(n12404) );
  AOI22_X1 U6128 ( .A1(ram[1105]), .A2(n5557), .B1(n12419), .B2(n8893), .ZN(
        n5558) );
  INV_X1 U6129 ( .A(n5559), .ZN(n12405) );
  AOI22_X1 U6130 ( .A1(ram[1106]), .A2(n5557), .B1(n12419), .B2(n8917), .ZN(
        n5559) );
  INV_X1 U6131 ( .A(n5560), .ZN(n12406) );
  AOI22_X1 U6132 ( .A1(ram[1107]), .A2(n5557), .B1(n12419), .B2(n8941), .ZN(
        n5560) );
  INV_X1 U6133 ( .A(n5561), .ZN(n12407) );
  AOI22_X1 U6134 ( .A1(ram[1108]), .A2(n5557), .B1(n12419), .B2(n8965), .ZN(
        n5561) );
  INV_X1 U6135 ( .A(n5562), .ZN(n12408) );
  AOI22_X1 U6136 ( .A1(ram[1109]), .A2(n5557), .B1(n12419), .B2(n8989), .ZN(
        n5562) );
  INV_X1 U6137 ( .A(n5563), .ZN(n12409) );
  AOI22_X1 U6138 ( .A1(ram[1110]), .A2(n5557), .B1(n12419), .B2(n9013), .ZN(
        n5563) );
  INV_X1 U6139 ( .A(n5564), .ZN(n12410) );
  AOI22_X1 U6140 ( .A1(ram[1111]), .A2(n5557), .B1(n12419), .B2(n9037), .ZN(
        n5564) );
  INV_X1 U6141 ( .A(n5565), .ZN(n12411) );
  AOI22_X1 U6142 ( .A1(ram[1112]), .A2(n5557), .B1(n12419), .B2(n9061), .ZN(
        n5565) );
  INV_X1 U6143 ( .A(n5566), .ZN(n12412) );
  AOI22_X1 U6144 ( .A1(ram[1113]), .A2(n5557), .B1(n12419), .B2(n9085), .ZN(
        n5566) );
  INV_X1 U6145 ( .A(n5567), .ZN(n12413) );
  AOI22_X1 U6146 ( .A1(ram[1114]), .A2(n5557), .B1(n12419), .B2(n9109), .ZN(
        n5567) );
  INV_X1 U6147 ( .A(n5568), .ZN(n12414) );
  AOI22_X1 U6148 ( .A1(ram[1115]), .A2(n5557), .B1(n12419), .B2(n9133), .ZN(
        n5568) );
  INV_X1 U6149 ( .A(n5569), .ZN(n12415) );
  AOI22_X1 U6150 ( .A1(ram[1116]), .A2(n5557), .B1(n12419), .B2(n9157), .ZN(
        n5569) );
  INV_X1 U6151 ( .A(n5570), .ZN(n12416) );
  AOI22_X1 U6152 ( .A1(ram[1117]), .A2(n5557), .B1(n12419), .B2(n9181), .ZN(
        n5570) );
  INV_X1 U6153 ( .A(n5571), .ZN(n12417) );
  AOI22_X1 U6154 ( .A1(ram[1118]), .A2(n5557), .B1(n12419), .B2(n9205), .ZN(
        n5571) );
  INV_X1 U6155 ( .A(n5572), .ZN(n12418) );
  AOI22_X1 U6156 ( .A1(ram[1119]), .A2(n5557), .B1(n12419), .B2(n9229), .ZN(
        n5572) );
  INV_X1 U6157 ( .A(n5590), .ZN(n12369) );
  AOI22_X1 U6158 ( .A1(ram[1136]), .A2(n5591), .B1(n12385), .B2(n8869), .ZN(
        n5590) );
  INV_X1 U6159 ( .A(n5592), .ZN(n12370) );
  AOI22_X1 U6160 ( .A1(ram[1137]), .A2(n5591), .B1(n12385), .B2(n8893), .ZN(
        n5592) );
  INV_X1 U6161 ( .A(n5593), .ZN(n12371) );
  AOI22_X1 U6162 ( .A1(ram[1138]), .A2(n5591), .B1(n12385), .B2(n8917), .ZN(
        n5593) );
  INV_X1 U6163 ( .A(n5594), .ZN(n12372) );
  AOI22_X1 U6164 ( .A1(ram[1139]), .A2(n5591), .B1(n12385), .B2(n8941), .ZN(
        n5594) );
  INV_X1 U6165 ( .A(n5595), .ZN(n12373) );
  AOI22_X1 U6166 ( .A1(ram[1140]), .A2(n5591), .B1(n12385), .B2(n8965), .ZN(
        n5595) );
  INV_X1 U6167 ( .A(n5596), .ZN(n12374) );
  AOI22_X1 U6168 ( .A1(ram[1141]), .A2(n5591), .B1(n12385), .B2(n8989), .ZN(
        n5596) );
  INV_X1 U6169 ( .A(n5597), .ZN(n12375) );
  AOI22_X1 U6170 ( .A1(ram[1142]), .A2(n5591), .B1(n12385), .B2(n9013), .ZN(
        n5597) );
  INV_X1 U6171 ( .A(n5598), .ZN(n12376) );
  AOI22_X1 U6172 ( .A1(ram[1143]), .A2(n5591), .B1(n12385), .B2(n9037), .ZN(
        n5598) );
  INV_X1 U6173 ( .A(n5599), .ZN(n12377) );
  AOI22_X1 U6174 ( .A1(ram[1144]), .A2(n5591), .B1(n12385), .B2(n9061), .ZN(
        n5599) );
  INV_X1 U6175 ( .A(n5600), .ZN(n12378) );
  AOI22_X1 U6176 ( .A1(ram[1145]), .A2(n5591), .B1(n12385), .B2(n9085), .ZN(
        n5600) );
  INV_X1 U6177 ( .A(n5601), .ZN(n12379) );
  AOI22_X1 U6178 ( .A1(ram[1146]), .A2(n5591), .B1(n12385), .B2(n9109), .ZN(
        n5601) );
  INV_X1 U6179 ( .A(n5602), .ZN(n12380) );
  AOI22_X1 U6180 ( .A1(ram[1147]), .A2(n5591), .B1(n12385), .B2(n9133), .ZN(
        n5602) );
  INV_X1 U6181 ( .A(n5603), .ZN(n12381) );
  AOI22_X1 U6182 ( .A1(ram[1148]), .A2(n5591), .B1(n12385), .B2(n9157), .ZN(
        n5603) );
  INV_X1 U6183 ( .A(n5604), .ZN(n12382) );
  AOI22_X1 U6184 ( .A1(ram[1149]), .A2(n5591), .B1(n12385), .B2(n9181), .ZN(
        n5604) );
  INV_X1 U6185 ( .A(n5605), .ZN(n12383) );
  AOI22_X1 U6186 ( .A1(ram[1150]), .A2(n5591), .B1(n12385), .B2(n9205), .ZN(
        n5605) );
  INV_X1 U6187 ( .A(n5606), .ZN(n12384) );
  AOI22_X1 U6188 ( .A1(ram[1151]), .A2(n5591), .B1(n12385), .B2(n9229), .ZN(
        n5606) );
  INV_X1 U6189 ( .A(n5624), .ZN(n12335) );
  AOI22_X1 U6190 ( .A1(ram[1168]), .A2(n5625), .B1(n12351), .B2(n8869), .ZN(
        n5624) );
  INV_X1 U6191 ( .A(n5626), .ZN(n12336) );
  AOI22_X1 U6192 ( .A1(ram[1169]), .A2(n5625), .B1(n12351), .B2(n8893), .ZN(
        n5626) );
  INV_X1 U6193 ( .A(n5627), .ZN(n12337) );
  AOI22_X1 U6194 ( .A1(ram[1170]), .A2(n5625), .B1(n12351), .B2(n8917), .ZN(
        n5627) );
  INV_X1 U6195 ( .A(n5628), .ZN(n12338) );
  AOI22_X1 U6196 ( .A1(ram[1171]), .A2(n5625), .B1(n12351), .B2(n8941), .ZN(
        n5628) );
  INV_X1 U6197 ( .A(n5629), .ZN(n12339) );
  AOI22_X1 U6198 ( .A1(ram[1172]), .A2(n5625), .B1(n12351), .B2(n8965), .ZN(
        n5629) );
  INV_X1 U6199 ( .A(n5630), .ZN(n12340) );
  AOI22_X1 U6200 ( .A1(ram[1173]), .A2(n5625), .B1(n12351), .B2(n8989), .ZN(
        n5630) );
  INV_X1 U6201 ( .A(n5631), .ZN(n12341) );
  AOI22_X1 U6202 ( .A1(ram[1174]), .A2(n5625), .B1(n12351), .B2(n9013), .ZN(
        n5631) );
  INV_X1 U6203 ( .A(n5632), .ZN(n12342) );
  AOI22_X1 U6204 ( .A1(ram[1175]), .A2(n5625), .B1(n12351), .B2(n9037), .ZN(
        n5632) );
  INV_X1 U6205 ( .A(n5633), .ZN(n12343) );
  AOI22_X1 U6206 ( .A1(ram[1176]), .A2(n5625), .B1(n12351), .B2(n9061), .ZN(
        n5633) );
  INV_X1 U6207 ( .A(n5634), .ZN(n12344) );
  AOI22_X1 U6208 ( .A1(ram[1177]), .A2(n5625), .B1(n12351), .B2(n9085), .ZN(
        n5634) );
  INV_X1 U6209 ( .A(n5635), .ZN(n12345) );
  AOI22_X1 U6210 ( .A1(ram[1178]), .A2(n5625), .B1(n12351), .B2(n9109), .ZN(
        n5635) );
  INV_X1 U6211 ( .A(n5636), .ZN(n12346) );
  AOI22_X1 U6212 ( .A1(ram[1179]), .A2(n5625), .B1(n12351), .B2(n9133), .ZN(
        n5636) );
  INV_X1 U6213 ( .A(n5637), .ZN(n12347) );
  AOI22_X1 U6214 ( .A1(ram[1180]), .A2(n5625), .B1(n12351), .B2(n9157), .ZN(
        n5637) );
  INV_X1 U6215 ( .A(n5638), .ZN(n12348) );
  AOI22_X1 U6216 ( .A1(ram[1181]), .A2(n5625), .B1(n12351), .B2(n9181), .ZN(
        n5638) );
  INV_X1 U6217 ( .A(n5639), .ZN(n12349) );
  AOI22_X1 U6218 ( .A1(ram[1182]), .A2(n5625), .B1(n12351), .B2(n9205), .ZN(
        n5639) );
  INV_X1 U6219 ( .A(n5640), .ZN(n12350) );
  AOI22_X1 U6220 ( .A1(ram[1183]), .A2(n5625), .B1(n12351), .B2(n9229), .ZN(
        n5640) );
  INV_X1 U6221 ( .A(n5658), .ZN(n12301) );
  AOI22_X1 U6222 ( .A1(ram[1200]), .A2(n5659), .B1(n12317), .B2(n8869), .ZN(
        n5658) );
  INV_X1 U6223 ( .A(n5660), .ZN(n12302) );
  AOI22_X1 U6224 ( .A1(ram[1201]), .A2(n5659), .B1(n12317), .B2(n8893), .ZN(
        n5660) );
  INV_X1 U6225 ( .A(n5661), .ZN(n12303) );
  AOI22_X1 U6226 ( .A1(ram[1202]), .A2(n5659), .B1(n12317), .B2(n8917), .ZN(
        n5661) );
  INV_X1 U6227 ( .A(n5662), .ZN(n12304) );
  AOI22_X1 U6228 ( .A1(ram[1203]), .A2(n5659), .B1(n12317), .B2(n8941), .ZN(
        n5662) );
  INV_X1 U6229 ( .A(n5663), .ZN(n12305) );
  AOI22_X1 U6230 ( .A1(ram[1204]), .A2(n5659), .B1(n12317), .B2(n8965), .ZN(
        n5663) );
  INV_X1 U6231 ( .A(n5664), .ZN(n12306) );
  AOI22_X1 U6232 ( .A1(ram[1205]), .A2(n5659), .B1(n12317), .B2(n8989), .ZN(
        n5664) );
  INV_X1 U6233 ( .A(n5665), .ZN(n12307) );
  AOI22_X1 U6234 ( .A1(ram[1206]), .A2(n5659), .B1(n12317), .B2(n9013), .ZN(
        n5665) );
  INV_X1 U6235 ( .A(n5666), .ZN(n12308) );
  AOI22_X1 U6236 ( .A1(ram[1207]), .A2(n5659), .B1(n12317), .B2(n9037), .ZN(
        n5666) );
  INV_X1 U6237 ( .A(n5667), .ZN(n12309) );
  AOI22_X1 U6238 ( .A1(ram[1208]), .A2(n5659), .B1(n12317), .B2(n9061), .ZN(
        n5667) );
  INV_X1 U6239 ( .A(n5668), .ZN(n12310) );
  AOI22_X1 U6240 ( .A1(ram[1209]), .A2(n5659), .B1(n12317), .B2(n9085), .ZN(
        n5668) );
  INV_X1 U6241 ( .A(n5669), .ZN(n12311) );
  AOI22_X1 U6242 ( .A1(ram[1210]), .A2(n5659), .B1(n12317), .B2(n9109), .ZN(
        n5669) );
  INV_X1 U6243 ( .A(n5670), .ZN(n12312) );
  AOI22_X1 U6244 ( .A1(ram[1211]), .A2(n5659), .B1(n12317), .B2(n9133), .ZN(
        n5670) );
  INV_X1 U6245 ( .A(n5671), .ZN(n12313) );
  AOI22_X1 U6246 ( .A1(ram[1212]), .A2(n5659), .B1(n12317), .B2(n9157), .ZN(
        n5671) );
  INV_X1 U6247 ( .A(n5672), .ZN(n12314) );
  AOI22_X1 U6248 ( .A1(ram[1213]), .A2(n5659), .B1(n12317), .B2(n9181), .ZN(
        n5672) );
  INV_X1 U6249 ( .A(n5673), .ZN(n12315) );
  AOI22_X1 U6250 ( .A1(ram[1214]), .A2(n5659), .B1(n12317), .B2(n9205), .ZN(
        n5673) );
  INV_X1 U6251 ( .A(n5674), .ZN(n12316) );
  AOI22_X1 U6252 ( .A1(ram[1215]), .A2(n5659), .B1(n12317), .B2(n9229), .ZN(
        n5674) );
  INV_X1 U6253 ( .A(n5692), .ZN(n12267) );
  AOI22_X1 U6254 ( .A1(ram[1232]), .A2(n5693), .B1(n12283), .B2(n8868), .ZN(
        n5692) );
  INV_X1 U6255 ( .A(n5694), .ZN(n12268) );
  AOI22_X1 U6256 ( .A1(ram[1233]), .A2(n5693), .B1(n12283), .B2(n8892), .ZN(
        n5694) );
  INV_X1 U6257 ( .A(n5695), .ZN(n12269) );
  AOI22_X1 U6258 ( .A1(ram[1234]), .A2(n5693), .B1(n12283), .B2(n8916), .ZN(
        n5695) );
  INV_X1 U6259 ( .A(n5696), .ZN(n12270) );
  AOI22_X1 U6260 ( .A1(ram[1235]), .A2(n5693), .B1(n12283), .B2(n8940), .ZN(
        n5696) );
  INV_X1 U6261 ( .A(n5697), .ZN(n12271) );
  AOI22_X1 U6262 ( .A1(ram[1236]), .A2(n5693), .B1(n12283), .B2(n8964), .ZN(
        n5697) );
  INV_X1 U6263 ( .A(n5698), .ZN(n12272) );
  AOI22_X1 U6264 ( .A1(ram[1237]), .A2(n5693), .B1(n12283), .B2(n8988), .ZN(
        n5698) );
  INV_X1 U6265 ( .A(n5699), .ZN(n12273) );
  AOI22_X1 U6266 ( .A1(ram[1238]), .A2(n5693), .B1(n12283), .B2(n9012), .ZN(
        n5699) );
  INV_X1 U6267 ( .A(n5700), .ZN(n12274) );
  AOI22_X1 U6268 ( .A1(ram[1239]), .A2(n5693), .B1(n12283), .B2(n9036), .ZN(
        n5700) );
  INV_X1 U6269 ( .A(n5701), .ZN(n12275) );
  AOI22_X1 U6270 ( .A1(ram[1240]), .A2(n5693), .B1(n12283), .B2(n9060), .ZN(
        n5701) );
  INV_X1 U6271 ( .A(n5702), .ZN(n12276) );
  AOI22_X1 U6272 ( .A1(ram[1241]), .A2(n5693), .B1(n12283), .B2(n9084), .ZN(
        n5702) );
  INV_X1 U6273 ( .A(n5703), .ZN(n12277) );
  AOI22_X1 U6274 ( .A1(ram[1242]), .A2(n5693), .B1(n12283), .B2(n9108), .ZN(
        n5703) );
  INV_X1 U6275 ( .A(n5704), .ZN(n12278) );
  AOI22_X1 U6276 ( .A1(ram[1243]), .A2(n5693), .B1(n12283), .B2(n9132), .ZN(
        n5704) );
  INV_X1 U6277 ( .A(n5705), .ZN(n12279) );
  AOI22_X1 U6278 ( .A1(ram[1244]), .A2(n5693), .B1(n12283), .B2(n9156), .ZN(
        n5705) );
  INV_X1 U6279 ( .A(n5706), .ZN(n12280) );
  AOI22_X1 U6280 ( .A1(ram[1245]), .A2(n5693), .B1(n12283), .B2(n9180), .ZN(
        n5706) );
  INV_X1 U6281 ( .A(n5707), .ZN(n12281) );
  AOI22_X1 U6282 ( .A1(ram[1246]), .A2(n5693), .B1(n12283), .B2(n9204), .ZN(
        n5707) );
  INV_X1 U6283 ( .A(n5708), .ZN(n12282) );
  AOI22_X1 U6284 ( .A1(ram[1247]), .A2(n5693), .B1(n12283), .B2(n9228), .ZN(
        n5708) );
  INV_X1 U6285 ( .A(n5726), .ZN(n12233) );
  AOI22_X1 U6286 ( .A1(ram[1264]), .A2(n5727), .B1(n12249), .B2(n8868), .ZN(
        n5726) );
  INV_X1 U6287 ( .A(n5728), .ZN(n12234) );
  AOI22_X1 U6288 ( .A1(ram[1265]), .A2(n5727), .B1(n12249), .B2(n8892), .ZN(
        n5728) );
  INV_X1 U6289 ( .A(n5729), .ZN(n12235) );
  AOI22_X1 U6290 ( .A1(ram[1266]), .A2(n5727), .B1(n12249), .B2(n8916), .ZN(
        n5729) );
  INV_X1 U6291 ( .A(n5730), .ZN(n12236) );
  AOI22_X1 U6292 ( .A1(ram[1267]), .A2(n5727), .B1(n12249), .B2(n8940), .ZN(
        n5730) );
  INV_X1 U6293 ( .A(n5731), .ZN(n12237) );
  AOI22_X1 U6294 ( .A1(ram[1268]), .A2(n5727), .B1(n12249), .B2(n8964), .ZN(
        n5731) );
  INV_X1 U6295 ( .A(n5732), .ZN(n12238) );
  AOI22_X1 U6296 ( .A1(ram[1269]), .A2(n5727), .B1(n12249), .B2(n8988), .ZN(
        n5732) );
  INV_X1 U6297 ( .A(n5733), .ZN(n12239) );
  AOI22_X1 U6298 ( .A1(ram[1270]), .A2(n5727), .B1(n12249), .B2(n9012), .ZN(
        n5733) );
  INV_X1 U6299 ( .A(n5734), .ZN(n12240) );
  AOI22_X1 U6300 ( .A1(ram[1271]), .A2(n5727), .B1(n12249), .B2(n9036), .ZN(
        n5734) );
  INV_X1 U6301 ( .A(n5735), .ZN(n12241) );
  AOI22_X1 U6302 ( .A1(ram[1272]), .A2(n5727), .B1(n12249), .B2(n9060), .ZN(
        n5735) );
  INV_X1 U6303 ( .A(n5736), .ZN(n12242) );
  AOI22_X1 U6304 ( .A1(ram[1273]), .A2(n5727), .B1(n12249), .B2(n9084), .ZN(
        n5736) );
  INV_X1 U6305 ( .A(n5737), .ZN(n12243) );
  AOI22_X1 U6306 ( .A1(ram[1274]), .A2(n5727), .B1(n12249), .B2(n9108), .ZN(
        n5737) );
  INV_X1 U6307 ( .A(n5738), .ZN(n12244) );
  AOI22_X1 U6308 ( .A1(ram[1275]), .A2(n5727), .B1(n12249), .B2(n9132), .ZN(
        n5738) );
  INV_X1 U6309 ( .A(n5739), .ZN(n12245) );
  AOI22_X1 U6310 ( .A1(ram[1276]), .A2(n5727), .B1(n12249), .B2(n9156), .ZN(
        n5739) );
  INV_X1 U6311 ( .A(n5740), .ZN(n12246) );
  AOI22_X1 U6312 ( .A1(ram[1277]), .A2(n5727), .B1(n12249), .B2(n9180), .ZN(
        n5740) );
  INV_X1 U6313 ( .A(n5741), .ZN(n12247) );
  AOI22_X1 U6314 ( .A1(ram[1278]), .A2(n5727), .B1(n12249), .B2(n9204), .ZN(
        n5741) );
  INV_X1 U6315 ( .A(n5742), .ZN(n12248) );
  AOI22_X1 U6316 ( .A1(ram[1279]), .A2(n5727), .B1(n12249), .B2(n9228), .ZN(
        n5742) );
  INV_X1 U6317 ( .A(n5762), .ZN(n12199) );
  AOI22_X1 U6318 ( .A1(ram[1296]), .A2(n5763), .B1(n12215), .B2(n8868), .ZN(
        n5762) );
  INV_X1 U6319 ( .A(n5764), .ZN(n12200) );
  AOI22_X1 U6320 ( .A1(ram[1297]), .A2(n5763), .B1(n12215), .B2(n8892), .ZN(
        n5764) );
  INV_X1 U6321 ( .A(n5765), .ZN(n12201) );
  AOI22_X1 U6322 ( .A1(ram[1298]), .A2(n5763), .B1(n12215), .B2(n8916), .ZN(
        n5765) );
  INV_X1 U6323 ( .A(n5766), .ZN(n12202) );
  AOI22_X1 U6324 ( .A1(ram[1299]), .A2(n5763), .B1(n12215), .B2(n8940), .ZN(
        n5766) );
  INV_X1 U6325 ( .A(n5767), .ZN(n12203) );
  AOI22_X1 U6326 ( .A1(ram[1300]), .A2(n5763), .B1(n12215), .B2(n8964), .ZN(
        n5767) );
  INV_X1 U6327 ( .A(n5768), .ZN(n12204) );
  AOI22_X1 U6328 ( .A1(ram[1301]), .A2(n5763), .B1(n12215), .B2(n8988), .ZN(
        n5768) );
  INV_X1 U6329 ( .A(n5769), .ZN(n12205) );
  AOI22_X1 U6330 ( .A1(ram[1302]), .A2(n5763), .B1(n12215), .B2(n9012), .ZN(
        n5769) );
  INV_X1 U6331 ( .A(n5770), .ZN(n12206) );
  AOI22_X1 U6332 ( .A1(ram[1303]), .A2(n5763), .B1(n12215), .B2(n9036), .ZN(
        n5770) );
  INV_X1 U6333 ( .A(n5771), .ZN(n12207) );
  AOI22_X1 U6334 ( .A1(ram[1304]), .A2(n5763), .B1(n12215), .B2(n9060), .ZN(
        n5771) );
  INV_X1 U6335 ( .A(n5772), .ZN(n12208) );
  AOI22_X1 U6336 ( .A1(ram[1305]), .A2(n5763), .B1(n12215), .B2(n9084), .ZN(
        n5772) );
  INV_X1 U6337 ( .A(n5773), .ZN(n12209) );
  AOI22_X1 U6338 ( .A1(ram[1306]), .A2(n5763), .B1(n12215), .B2(n9108), .ZN(
        n5773) );
  INV_X1 U6339 ( .A(n5774), .ZN(n12210) );
  AOI22_X1 U6340 ( .A1(ram[1307]), .A2(n5763), .B1(n12215), .B2(n9132), .ZN(
        n5774) );
  INV_X1 U6341 ( .A(n5775), .ZN(n12211) );
  AOI22_X1 U6342 ( .A1(ram[1308]), .A2(n5763), .B1(n12215), .B2(n9156), .ZN(
        n5775) );
  INV_X1 U6343 ( .A(n5776), .ZN(n12212) );
  AOI22_X1 U6344 ( .A1(ram[1309]), .A2(n5763), .B1(n12215), .B2(n9180), .ZN(
        n5776) );
  INV_X1 U6345 ( .A(n5777), .ZN(n12213) );
  AOI22_X1 U6346 ( .A1(ram[1310]), .A2(n5763), .B1(n12215), .B2(n9204), .ZN(
        n5777) );
  INV_X1 U6347 ( .A(n5778), .ZN(n12214) );
  AOI22_X1 U6348 ( .A1(ram[1311]), .A2(n5763), .B1(n12215), .B2(n9228), .ZN(
        n5778) );
  INV_X1 U6349 ( .A(n5796), .ZN(n12165) );
  AOI22_X1 U6350 ( .A1(ram[1328]), .A2(n5797), .B1(n12181), .B2(n8868), .ZN(
        n5796) );
  INV_X1 U6351 ( .A(n5798), .ZN(n12166) );
  AOI22_X1 U6352 ( .A1(ram[1329]), .A2(n5797), .B1(n12181), .B2(n8892), .ZN(
        n5798) );
  INV_X1 U6353 ( .A(n5799), .ZN(n12167) );
  AOI22_X1 U6354 ( .A1(ram[1330]), .A2(n5797), .B1(n12181), .B2(n8916), .ZN(
        n5799) );
  INV_X1 U6355 ( .A(n5800), .ZN(n12168) );
  AOI22_X1 U6356 ( .A1(ram[1331]), .A2(n5797), .B1(n12181), .B2(n8940), .ZN(
        n5800) );
  INV_X1 U6357 ( .A(n5801), .ZN(n12169) );
  AOI22_X1 U6358 ( .A1(ram[1332]), .A2(n5797), .B1(n12181), .B2(n8964), .ZN(
        n5801) );
  INV_X1 U6359 ( .A(n5802), .ZN(n12170) );
  AOI22_X1 U6360 ( .A1(ram[1333]), .A2(n5797), .B1(n12181), .B2(n8988), .ZN(
        n5802) );
  INV_X1 U6361 ( .A(n5803), .ZN(n12171) );
  AOI22_X1 U6362 ( .A1(ram[1334]), .A2(n5797), .B1(n12181), .B2(n9012), .ZN(
        n5803) );
  INV_X1 U6363 ( .A(n5804), .ZN(n12172) );
  AOI22_X1 U6364 ( .A1(ram[1335]), .A2(n5797), .B1(n12181), .B2(n9036), .ZN(
        n5804) );
  INV_X1 U6365 ( .A(n5805), .ZN(n12173) );
  AOI22_X1 U6366 ( .A1(ram[1336]), .A2(n5797), .B1(n12181), .B2(n9060), .ZN(
        n5805) );
  INV_X1 U6367 ( .A(n5806), .ZN(n12174) );
  AOI22_X1 U6368 ( .A1(ram[1337]), .A2(n5797), .B1(n12181), .B2(n9084), .ZN(
        n5806) );
  INV_X1 U6369 ( .A(n5807), .ZN(n12175) );
  AOI22_X1 U6370 ( .A1(ram[1338]), .A2(n5797), .B1(n12181), .B2(n9108), .ZN(
        n5807) );
  INV_X1 U6371 ( .A(n5808), .ZN(n12176) );
  AOI22_X1 U6372 ( .A1(ram[1339]), .A2(n5797), .B1(n12181), .B2(n9132), .ZN(
        n5808) );
  INV_X1 U6373 ( .A(n5809), .ZN(n12177) );
  AOI22_X1 U6374 ( .A1(ram[1340]), .A2(n5797), .B1(n12181), .B2(n9156), .ZN(
        n5809) );
  INV_X1 U6375 ( .A(n5810), .ZN(n12178) );
  AOI22_X1 U6376 ( .A1(ram[1341]), .A2(n5797), .B1(n12181), .B2(n9180), .ZN(
        n5810) );
  INV_X1 U6377 ( .A(n5811), .ZN(n12179) );
  AOI22_X1 U6378 ( .A1(ram[1342]), .A2(n5797), .B1(n12181), .B2(n9204), .ZN(
        n5811) );
  INV_X1 U6379 ( .A(n5812), .ZN(n12180) );
  AOI22_X1 U6380 ( .A1(ram[1343]), .A2(n5797), .B1(n12181), .B2(n9228), .ZN(
        n5812) );
  INV_X1 U6381 ( .A(n5830), .ZN(n12131) );
  AOI22_X1 U6382 ( .A1(ram[1360]), .A2(n5831), .B1(n12147), .B2(n8868), .ZN(
        n5830) );
  INV_X1 U6383 ( .A(n5832), .ZN(n12132) );
  AOI22_X1 U6384 ( .A1(ram[1361]), .A2(n5831), .B1(n12147), .B2(n8892), .ZN(
        n5832) );
  INV_X1 U6385 ( .A(n5833), .ZN(n12133) );
  AOI22_X1 U6386 ( .A1(ram[1362]), .A2(n5831), .B1(n12147), .B2(n8916), .ZN(
        n5833) );
  INV_X1 U6387 ( .A(n5834), .ZN(n12134) );
  AOI22_X1 U6388 ( .A1(ram[1363]), .A2(n5831), .B1(n12147), .B2(n8940), .ZN(
        n5834) );
  INV_X1 U6389 ( .A(n5835), .ZN(n12135) );
  AOI22_X1 U6390 ( .A1(ram[1364]), .A2(n5831), .B1(n12147), .B2(n8964), .ZN(
        n5835) );
  INV_X1 U6391 ( .A(n5836), .ZN(n12136) );
  AOI22_X1 U6392 ( .A1(ram[1365]), .A2(n5831), .B1(n12147), .B2(n8988), .ZN(
        n5836) );
  INV_X1 U6393 ( .A(n5837), .ZN(n12137) );
  AOI22_X1 U6394 ( .A1(ram[1366]), .A2(n5831), .B1(n12147), .B2(n9012), .ZN(
        n5837) );
  INV_X1 U6395 ( .A(n5838), .ZN(n12138) );
  AOI22_X1 U6396 ( .A1(ram[1367]), .A2(n5831), .B1(n12147), .B2(n9036), .ZN(
        n5838) );
  INV_X1 U6397 ( .A(n5839), .ZN(n12139) );
  AOI22_X1 U6398 ( .A1(ram[1368]), .A2(n5831), .B1(n12147), .B2(n9060), .ZN(
        n5839) );
  INV_X1 U6399 ( .A(n5840), .ZN(n12140) );
  AOI22_X1 U6400 ( .A1(ram[1369]), .A2(n5831), .B1(n12147), .B2(n9084), .ZN(
        n5840) );
  INV_X1 U6401 ( .A(n5841), .ZN(n12141) );
  AOI22_X1 U6402 ( .A1(ram[1370]), .A2(n5831), .B1(n12147), .B2(n9108), .ZN(
        n5841) );
  INV_X1 U6403 ( .A(n5842), .ZN(n12142) );
  AOI22_X1 U6404 ( .A1(ram[1371]), .A2(n5831), .B1(n12147), .B2(n9132), .ZN(
        n5842) );
  INV_X1 U6405 ( .A(n5843), .ZN(n12143) );
  AOI22_X1 U6406 ( .A1(ram[1372]), .A2(n5831), .B1(n12147), .B2(n9156), .ZN(
        n5843) );
  INV_X1 U6407 ( .A(n5844), .ZN(n12144) );
  AOI22_X1 U6408 ( .A1(ram[1373]), .A2(n5831), .B1(n12147), .B2(n9180), .ZN(
        n5844) );
  INV_X1 U6409 ( .A(n5845), .ZN(n12145) );
  AOI22_X1 U6410 ( .A1(ram[1374]), .A2(n5831), .B1(n12147), .B2(n9204), .ZN(
        n5845) );
  INV_X1 U6411 ( .A(n5846), .ZN(n12146) );
  AOI22_X1 U6412 ( .A1(ram[1375]), .A2(n5831), .B1(n12147), .B2(n9228), .ZN(
        n5846) );
  INV_X1 U6413 ( .A(n5864), .ZN(n12097) );
  AOI22_X1 U6414 ( .A1(ram[1392]), .A2(n5865), .B1(n12113), .B2(n8868), .ZN(
        n5864) );
  INV_X1 U6415 ( .A(n5866), .ZN(n12098) );
  AOI22_X1 U6416 ( .A1(ram[1393]), .A2(n5865), .B1(n12113), .B2(n8892), .ZN(
        n5866) );
  INV_X1 U6417 ( .A(n5867), .ZN(n12099) );
  AOI22_X1 U6418 ( .A1(ram[1394]), .A2(n5865), .B1(n12113), .B2(n8916), .ZN(
        n5867) );
  INV_X1 U6419 ( .A(n5868), .ZN(n12100) );
  AOI22_X1 U6420 ( .A1(ram[1395]), .A2(n5865), .B1(n12113), .B2(n8940), .ZN(
        n5868) );
  INV_X1 U6421 ( .A(n5869), .ZN(n12101) );
  AOI22_X1 U6422 ( .A1(ram[1396]), .A2(n5865), .B1(n12113), .B2(n8964), .ZN(
        n5869) );
  INV_X1 U6423 ( .A(n5870), .ZN(n12102) );
  AOI22_X1 U6424 ( .A1(ram[1397]), .A2(n5865), .B1(n12113), .B2(n8988), .ZN(
        n5870) );
  INV_X1 U6425 ( .A(n5871), .ZN(n12103) );
  AOI22_X1 U6426 ( .A1(ram[1398]), .A2(n5865), .B1(n12113), .B2(n9012), .ZN(
        n5871) );
  INV_X1 U6427 ( .A(n5872), .ZN(n12104) );
  AOI22_X1 U6428 ( .A1(ram[1399]), .A2(n5865), .B1(n12113), .B2(n9036), .ZN(
        n5872) );
  INV_X1 U6429 ( .A(n5873), .ZN(n12105) );
  AOI22_X1 U6430 ( .A1(ram[1400]), .A2(n5865), .B1(n12113), .B2(n9060), .ZN(
        n5873) );
  INV_X1 U6431 ( .A(n5874), .ZN(n12106) );
  AOI22_X1 U6432 ( .A1(ram[1401]), .A2(n5865), .B1(n12113), .B2(n9084), .ZN(
        n5874) );
  INV_X1 U6433 ( .A(n5875), .ZN(n12107) );
  AOI22_X1 U6434 ( .A1(ram[1402]), .A2(n5865), .B1(n12113), .B2(n9108), .ZN(
        n5875) );
  INV_X1 U6435 ( .A(n5876), .ZN(n12108) );
  AOI22_X1 U6436 ( .A1(ram[1403]), .A2(n5865), .B1(n12113), .B2(n9132), .ZN(
        n5876) );
  INV_X1 U6437 ( .A(n5877), .ZN(n12109) );
  AOI22_X1 U6438 ( .A1(ram[1404]), .A2(n5865), .B1(n12113), .B2(n9156), .ZN(
        n5877) );
  INV_X1 U6439 ( .A(n5878), .ZN(n12110) );
  AOI22_X1 U6440 ( .A1(ram[1405]), .A2(n5865), .B1(n12113), .B2(n9180), .ZN(
        n5878) );
  INV_X1 U6441 ( .A(n5879), .ZN(n12111) );
  AOI22_X1 U6442 ( .A1(ram[1406]), .A2(n5865), .B1(n12113), .B2(n9204), .ZN(
        n5879) );
  INV_X1 U6443 ( .A(n5880), .ZN(n12112) );
  AOI22_X1 U6444 ( .A1(ram[1407]), .A2(n5865), .B1(n12113), .B2(n9228), .ZN(
        n5880) );
  INV_X1 U6445 ( .A(n5898), .ZN(n12063) );
  AOI22_X1 U6446 ( .A1(ram[1424]), .A2(n5899), .B1(n12079), .B2(n8867), .ZN(
        n5898) );
  INV_X1 U6447 ( .A(n5900), .ZN(n12064) );
  AOI22_X1 U6448 ( .A1(ram[1425]), .A2(n5899), .B1(n12079), .B2(n8891), .ZN(
        n5900) );
  INV_X1 U6449 ( .A(n5901), .ZN(n12065) );
  AOI22_X1 U6450 ( .A1(ram[1426]), .A2(n5899), .B1(n12079), .B2(n8915), .ZN(
        n5901) );
  INV_X1 U6451 ( .A(n5902), .ZN(n12066) );
  AOI22_X1 U6452 ( .A1(ram[1427]), .A2(n5899), .B1(n12079), .B2(n8939), .ZN(
        n5902) );
  INV_X1 U6453 ( .A(n5903), .ZN(n12067) );
  AOI22_X1 U6454 ( .A1(ram[1428]), .A2(n5899), .B1(n12079), .B2(n8963), .ZN(
        n5903) );
  INV_X1 U6455 ( .A(n5904), .ZN(n12068) );
  AOI22_X1 U6456 ( .A1(ram[1429]), .A2(n5899), .B1(n12079), .B2(n8987), .ZN(
        n5904) );
  INV_X1 U6457 ( .A(n5905), .ZN(n12069) );
  AOI22_X1 U6458 ( .A1(ram[1430]), .A2(n5899), .B1(n12079), .B2(n9011), .ZN(
        n5905) );
  INV_X1 U6459 ( .A(n5906), .ZN(n12070) );
  AOI22_X1 U6460 ( .A1(ram[1431]), .A2(n5899), .B1(n12079), .B2(n9035), .ZN(
        n5906) );
  INV_X1 U6461 ( .A(n5907), .ZN(n12071) );
  AOI22_X1 U6462 ( .A1(ram[1432]), .A2(n5899), .B1(n12079), .B2(n9059), .ZN(
        n5907) );
  INV_X1 U6463 ( .A(n5908), .ZN(n12072) );
  AOI22_X1 U6464 ( .A1(ram[1433]), .A2(n5899), .B1(n12079), .B2(n9083), .ZN(
        n5908) );
  INV_X1 U6465 ( .A(n5909), .ZN(n12073) );
  AOI22_X1 U6466 ( .A1(ram[1434]), .A2(n5899), .B1(n12079), .B2(n9107), .ZN(
        n5909) );
  INV_X1 U6467 ( .A(n5910), .ZN(n12074) );
  AOI22_X1 U6468 ( .A1(ram[1435]), .A2(n5899), .B1(n12079), .B2(n9131), .ZN(
        n5910) );
  INV_X1 U6469 ( .A(n5911), .ZN(n12075) );
  AOI22_X1 U6470 ( .A1(ram[1436]), .A2(n5899), .B1(n12079), .B2(n9155), .ZN(
        n5911) );
  INV_X1 U6471 ( .A(n5912), .ZN(n12076) );
  AOI22_X1 U6472 ( .A1(ram[1437]), .A2(n5899), .B1(n12079), .B2(n9179), .ZN(
        n5912) );
  INV_X1 U6473 ( .A(n5913), .ZN(n12077) );
  AOI22_X1 U6474 ( .A1(ram[1438]), .A2(n5899), .B1(n12079), .B2(n9203), .ZN(
        n5913) );
  INV_X1 U6475 ( .A(n5914), .ZN(n12078) );
  AOI22_X1 U6476 ( .A1(ram[1439]), .A2(n5899), .B1(n12079), .B2(n9227), .ZN(
        n5914) );
  INV_X1 U6477 ( .A(n5932), .ZN(n12029) );
  AOI22_X1 U6478 ( .A1(ram[1456]), .A2(n5933), .B1(n12045), .B2(n8867), .ZN(
        n5932) );
  INV_X1 U6479 ( .A(n5934), .ZN(n12030) );
  AOI22_X1 U6480 ( .A1(ram[1457]), .A2(n5933), .B1(n12045), .B2(n8891), .ZN(
        n5934) );
  INV_X1 U6481 ( .A(n5935), .ZN(n12031) );
  AOI22_X1 U6482 ( .A1(ram[1458]), .A2(n5933), .B1(n12045), .B2(n8915), .ZN(
        n5935) );
  INV_X1 U6483 ( .A(n5936), .ZN(n12032) );
  AOI22_X1 U6484 ( .A1(ram[1459]), .A2(n5933), .B1(n12045), .B2(n8939), .ZN(
        n5936) );
  INV_X1 U6485 ( .A(n5937), .ZN(n12033) );
  AOI22_X1 U6486 ( .A1(ram[1460]), .A2(n5933), .B1(n12045), .B2(n8963), .ZN(
        n5937) );
  INV_X1 U6487 ( .A(n5938), .ZN(n12034) );
  AOI22_X1 U6488 ( .A1(ram[1461]), .A2(n5933), .B1(n12045), .B2(n8987), .ZN(
        n5938) );
  INV_X1 U6489 ( .A(n5939), .ZN(n12035) );
  AOI22_X1 U6490 ( .A1(ram[1462]), .A2(n5933), .B1(n12045), .B2(n9011), .ZN(
        n5939) );
  INV_X1 U6491 ( .A(n5940), .ZN(n12036) );
  AOI22_X1 U6492 ( .A1(ram[1463]), .A2(n5933), .B1(n12045), .B2(n9035), .ZN(
        n5940) );
  INV_X1 U6493 ( .A(n5941), .ZN(n12037) );
  AOI22_X1 U6494 ( .A1(ram[1464]), .A2(n5933), .B1(n12045), .B2(n9059), .ZN(
        n5941) );
  INV_X1 U6495 ( .A(n5942), .ZN(n12038) );
  AOI22_X1 U6496 ( .A1(ram[1465]), .A2(n5933), .B1(n12045), .B2(n9083), .ZN(
        n5942) );
  INV_X1 U6497 ( .A(n5943), .ZN(n12039) );
  AOI22_X1 U6498 ( .A1(ram[1466]), .A2(n5933), .B1(n12045), .B2(n9107), .ZN(
        n5943) );
  INV_X1 U6499 ( .A(n5944), .ZN(n12040) );
  AOI22_X1 U6500 ( .A1(ram[1467]), .A2(n5933), .B1(n12045), .B2(n9131), .ZN(
        n5944) );
  INV_X1 U6501 ( .A(n5945), .ZN(n12041) );
  AOI22_X1 U6502 ( .A1(ram[1468]), .A2(n5933), .B1(n12045), .B2(n9155), .ZN(
        n5945) );
  INV_X1 U6503 ( .A(n5946), .ZN(n12042) );
  AOI22_X1 U6504 ( .A1(ram[1469]), .A2(n5933), .B1(n12045), .B2(n9179), .ZN(
        n5946) );
  INV_X1 U6505 ( .A(n5947), .ZN(n12043) );
  AOI22_X1 U6506 ( .A1(ram[1470]), .A2(n5933), .B1(n12045), .B2(n9203), .ZN(
        n5947) );
  INV_X1 U6507 ( .A(n5948), .ZN(n12044) );
  AOI22_X1 U6508 ( .A1(ram[1471]), .A2(n5933), .B1(n12045), .B2(n9227), .ZN(
        n5948) );
  INV_X1 U6509 ( .A(n5966), .ZN(n11995) );
  AOI22_X1 U6510 ( .A1(ram[1488]), .A2(n5967), .B1(n12011), .B2(n8867), .ZN(
        n5966) );
  INV_X1 U6511 ( .A(n5968), .ZN(n11996) );
  AOI22_X1 U6512 ( .A1(ram[1489]), .A2(n5967), .B1(n12011), .B2(n8891), .ZN(
        n5968) );
  INV_X1 U6513 ( .A(n5969), .ZN(n11997) );
  AOI22_X1 U6514 ( .A1(ram[1490]), .A2(n5967), .B1(n12011), .B2(n8915), .ZN(
        n5969) );
  INV_X1 U6515 ( .A(n5970), .ZN(n11998) );
  AOI22_X1 U6516 ( .A1(ram[1491]), .A2(n5967), .B1(n12011), .B2(n8939), .ZN(
        n5970) );
  INV_X1 U6517 ( .A(n5971), .ZN(n11999) );
  AOI22_X1 U6518 ( .A1(ram[1492]), .A2(n5967), .B1(n12011), .B2(n8963), .ZN(
        n5971) );
  INV_X1 U6519 ( .A(n5972), .ZN(n12000) );
  AOI22_X1 U6520 ( .A1(ram[1493]), .A2(n5967), .B1(n12011), .B2(n8987), .ZN(
        n5972) );
  INV_X1 U6521 ( .A(n5973), .ZN(n12001) );
  AOI22_X1 U6522 ( .A1(ram[1494]), .A2(n5967), .B1(n12011), .B2(n9011), .ZN(
        n5973) );
  INV_X1 U6523 ( .A(n5974), .ZN(n12002) );
  AOI22_X1 U6524 ( .A1(ram[1495]), .A2(n5967), .B1(n12011), .B2(n9035), .ZN(
        n5974) );
  INV_X1 U6525 ( .A(n5975), .ZN(n12003) );
  AOI22_X1 U6526 ( .A1(ram[1496]), .A2(n5967), .B1(n12011), .B2(n9059), .ZN(
        n5975) );
  INV_X1 U6527 ( .A(n5976), .ZN(n12004) );
  AOI22_X1 U6528 ( .A1(ram[1497]), .A2(n5967), .B1(n12011), .B2(n9083), .ZN(
        n5976) );
  INV_X1 U6529 ( .A(n5977), .ZN(n12005) );
  AOI22_X1 U6530 ( .A1(ram[1498]), .A2(n5967), .B1(n12011), .B2(n9107), .ZN(
        n5977) );
  INV_X1 U6531 ( .A(n5978), .ZN(n12006) );
  AOI22_X1 U6532 ( .A1(ram[1499]), .A2(n5967), .B1(n12011), .B2(n9131), .ZN(
        n5978) );
  INV_X1 U6533 ( .A(n5979), .ZN(n12007) );
  AOI22_X1 U6534 ( .A1(ram[1500]), .A2(n5967), .B1(n12011), .B2(n9155), .ZN(
        n5979) );
  INV_X1 U6535 ( .A(n5980), .ZN(n12008) );
  AOI22_X1 U6536 ( .A1(ram[1501]), .A2(n5967), .B1(n12011), .B2(n9179), .ZN(
        n5980) );
  INV_X1 U6537 ( .A(n5981), .ZN(n12009) );
  AOI22_X1 U6538 ( .A1(ram[1502]), .A2(n5967), .B1(n12011), .B2(n9203), .ZN(
        n5981) );
  INV_X1 U6539 ( .A(n5982), .ZN(n12010) );
  AOI22_X1 U6540 ( .A1(ram[1503]), .A2(n5967), .B1(n12011), .B2(n9227), .ZN(
        n5982) );
  INV_X1 U6541 ( .A(n6000), .ZN(n11961) );
  AOI22_X1 U6542 ( .A1(ram[1520]), .A2(n6001), .B1(n11977), .B2(n8867), .ZN(
        n6000) );
  INV_X1 U6543 ( .A(n6002), .ZN(n11962) );
  AOI22_X1 U6544 ( .A1(ram[1521]), .A2(n6001), .B1(n11977), .B2(n8891), .ZN(
        n6002) );
  INV_X1 U6545 ( .A(n6003), .ZN(n11963) );
  AOI22_X1 U6546 ( .A1(ram[1522]), .A2(n6001), .B1(n11977), .B2(n8915), .ZN(
        n6003) );
  INV_X1 U6547 ( .A(n6004), .ZN(n11964) );
  AOI22_X1 U6548 ( .A1(ram[1523]), .A2(n6001), .B1(n11977), .B2(n8939), .ZN(
        n6004) );
  INV_X1 U6549 ( .A(n6005), .ZN(n11965) );
  AOI22_X1 U6550 ( .A1(ram[1524]), .A2(n6001), .B1(n11977), .B2(n8963), .ZN(
        n6005) );
  INV_X1 U6551 ( .A(n6006), .ZN(n11966) );
  AOI22_X1 U6552 ( .A1(ram[1525]), .A2(n6001), .B1(n11977), .B2(n8987), .ZN(
        n6006) );
  INV_X1 U6553 ( .A(n6007), .ZN(n11967) );
  AOI22_X1 U6554 ( .A1(ram[1526]), .A2(n6001), .B1(n11977), .B2(n9011), .ZN(
        n6007) );
  INV_X1 U6555 ( .A(n6008), .ZN(n11968) );
  AOI22_X1 U6556 ( .A1(ram[1527]), .A2(n6001), .B1(n11977), .B2(n9035), .ZN(
        n6008) );
  INV_X1 U6557 ( .A(n6009), .ZN(n11969) );
  AOI22_X1 U6558 ( .A1(ram[1528]), .A2(n6001), .B1(n11977), .B2(n9059), .ZN(
        n6009) );
  INV_X1 U6559 ( .A(n6010), .ZN(n11970) );
  AOI22_X1 U6560 ( .A1(ram[1529]), .A2(n6001), .B1(n11977), .B2(n9083), .ZN(
        n6010) );
  INV_X1 U6561 ( .A(n6011), .ZN(n11971) );
  AOI22_X1 U6562 ( .A1(ram[1530]), .A2(n6001), .B1(n11977), .B2(n9107), .ZN(
        n6011) );
  INV_X1 U6563 ( .A(n6012), .ZN(n11972) );
  AOI22_X1 U6564 ( .A1(ram[1531]), .A2(n6001), .B1(n11977), .B2(n9131), .ZN(
        n6012) );
  INV_X1 U6565 ( .A(n6013), .ZN(n11973) );
  AOI22_X1 U6566 ( .A1(ram[1532]), .A2(n6001), .B1(n11977), .B2(n9155), .ZN(
        n6013) );
  INV_X1 U6567 ( .A(n6014), .ZN(n11974) );
  AOI22_X1 U6568 ( .A1(ram[1533]), .A2(n6001), .B1(n11977), .B2(n9179), .ZN(
        n6014) );
  INV_X1 U6569 ( .A(n6015), .ZN(n11975) );
  AOI22_X1 U6570 ( .A1(ram[1534]), .A2(n6001), .B1(n11977), .B2(n9203), .ZN(
        n6015) );
  INV_X1 U6571 ( .A(n6016), .ZN(n11976) );
  AOI22_X1 U6572 ( .A1(ram[1535]), .A2(n6001), .B1(n11977), .B2(n9227), .ZN(
        n6016) );
  INV_X1 U6573 ( .A(n6035), .ZN(n11927) );
  AOI22_X1 U6574 ( .A1(ram[1552]), .A2(n6036), .B1(n11943), .B2(n8867), .ZN(
        n6035) );
  INV_X1 U6575 ( .A(n6037), .ZN(n11928) );
  AOI22_X1 U6576 ( .A1(ram[1553]), .A2(n6036), .B1(n11943), .B2(n8891), .ZN(
        n6037) );
  INV_X1 U6577 ( .A(n6038), .ZN(n11929) );
  AOI22_X1 U6578 ( .A1(ram[1554]), .A2(n6036), .B1(n11943), .B2(n8915), .ZN(
        n6038) );
  INV_X1 U6579 ( .A(n6039), .ZN(n11930) );
  AOI22_X1 U6580 ( .A1(ram[1555]), .A2(n6036), .B1(n11943), .B2(n8939), .ZN(
        n6039) );
  INV_X1 U6581 ( .A(n6040), .ZN(n11931) );
  AOI22_X1 U6582 ( .A1(ram[1556]), .A2(n6036), .B1(n11943), .B2(n8963), .ZN(
        n6040) );
  INV_X1 U6583 ( .A(n6041), .ZN(n11932) );
  AOI22_X1 U6584 ( .A1(ram[1557]), .A2(n6036), .B1(n11943), .B2(n8987), .ZN(
        n6041) );
  INV_X1 U6585 ( .A(n6042), .ZN(n11933) );
  AOI22_X1 U6586 ( .A1(ram[1558]), .A2(n6036), .B1(n11943), .B2(n9011), .ZN(
        n6042) );
  INV_X1 U6587 ( .A(n6043), .ZN(n11934) );
  AOI22_X1 U6588 ( .A1(ram[1559]), .A2(n6036), .B1(n11943), .B2(n9035), .ZN(
        n6043) );
  INV_X1 U6589 ( .A(n6044), .ZN(n11935) );
  AOI22_X1 U6590 ( .A1(ram[1560]), .A2(n6036), .B1(n11943), .B2(n9059), .ZN(
        n6044) );
  INV_X1 U6591 ( .A(n6045), .ZN(n11936) );
  AOI22_X1 U6592 ( .A1(ram[1561]), .A2(n6036), .B1(n11943), .B2(n9083), .ZN(
        n6045) );
  INV_X1 U6593 ( .A(n6046), .ZN(n11937) );
  AOI22_X1 U6594 ( .A1(ram[1562]), .A2(n6036), .B1(n11943), .B2(n9107), .ZN(
        n6046) );
  INV_X1 U6595 ( .A(n6047), .ZN(n11938) );
  AOI22_X1 U6596 ( .A1(ram[1563]), .A2(n6036), .B1(n11943), .B2(n9131), .ZN(
        n6047) );
  INV_X1 U6597 ( .A(n6048), .ZN(n11939) );
  AOI22_X1 U6598 ( .A1(ram[1564]), .A2(n6036), .B1(n11943), .B2(n9155), .ZN(
        n6048) );
  INV_X1 U6599 ( .A(n6049), .ZN(n11940) );
  AOI22_X1 U6600 ( .A1(ram[1565]), .A2(n6036), .B1(n11943), .B2(n9179), .ZN(
        n6049) );
  INV_X1 U6601 ( .A(n6050), .ZN(n11941) );
  AOI22_X1 U6602 ( .A1(ram[1566]), .A2(n6036), .B1(n11943), .B2(n9203), .ZN(
        n6050) );
  INV_X1 U6603 ( .A(n6051), .ZN(n11942) );
  AOI22_X1 U6604 ( .A1(ram[1567]), .A2(n6036), .B1(n11943), .B2(n9227), .ZN(
        n6051) );
  INV_X1 U6605 ( .A(n6069), .ZN(n11893) );
  AOI22_X1 U6606 ( .A1(ram[1584]), .A2(n6070), .B1(n11909), .B2(n8867), .ZN(
        n6069) );
  INV_X1 U6607 ( .A(n6071), .ZN(n11894) );
  AOI22_X1 U6608 ( .A1(ram[1585]), .A2(n6070), .B1(n11909), .B2(n8891), .ZN(
        n6071) );
  INV_X1 U6609 ( .A(n6072), .ZN(n11895) );
  AOI22_X1 U6610 ( .A1(ram[1586]), .A2(n6070), .B1(n11909), .B2(n8915), .ZN(
        n6072) );
  INV_X1 U6611 ( .A(n6073), .ZN(n11896) );
  AOI22_X1 U6612 ( .A1(ram[1587]), .A2(n6070), .B1(n11909), .B2(n8939), .ZN(
        n6073) );
  INV_X1 U6613 ( .A(n6074), .ZN(n11897) );
  AOI22_X1 U6614 ( .A1(ram[1588]), .A2(n6070), .B1(n11909), .B2(n8963), .ZN(
        n6074) );
  INV_X1 U6615 ( .A(n6075), .ZN(n11898) );
  AOI22_X1 U6616 ( .A1(ram[1589]), .A2(n6070), .B1(n11909), .B2(n8987), .ZN(
        n6075) );
  INV_X1 U6617 ( .A(n6076), .ZN(n11899) );
  AOI22_X1 U6618 ( .A1(ram[1590]), .A2(n6070), .B1(n11909), .B2(n9011), .ZN(
        n6076) );
  INV_X1 U6619 ( .A(n6077), .ZN(n11900) );
  AOI22_X1 U6620 ( .A1(ram[1591]), .A2(n6070), .B1(n11909), .B2(n9035), .ZN(
        n6077) );
  INV_X1 U6621 ( .A(n6078), .ZN(n11901) );
  AOI22_X1 U6622 ( .A1(ram[1592]), .A2(n6070), .B1(n11909), .B2(n9059), .ZN(
        n6078) );
  INV_X1 U6623 ( .A(n6079), .ZN(n11902) );
  AOI22_X1 U6624 ( .A1(ram[1593]), .A2(n6070), .B1(n11909), .B2(n9083), .ZN(
        n6079) );
  INV_X1 U6625 ( .A(n6080), .ZN(n11903) );
  AOI22_X1 U6626 ( .A1(ram[1594]), .A2(n6070), .B1(n11909), .B2(n9107), .ZN(
        n6080) );
  INV_X1 U6627 ( .A(n6081), .ZN(n11904) );
  AOI22_X1 U6628 ( .A1(ram[1595]), .A2(n6070), .B1(n11909), .B2(n9131), .ZN(
        n6081) );
  INV_X1 U6629 ( .A(n6082), .ZN(n11905) );
  AOI22_X1 U6630 ( .A1(ram[1596]), .A2(n6070), .B1(n11909), .B2(n9155), .ZN(
        n6082) );
  INV_X1 U6631 ( .A(n6083), .ZN(n11906) );
  AOI22_X1 U6632 ( .A1(ram[1597]), .A2(n6070), .B1(n11909), .B2(n9179), .ZN(
        n6083) );
  INV_X1 U6633 ( .A(n6084), .ZN(n11907) );
  AOI22_X1 U6634 ( .A1(ram[1598]), .A2(n6070), .B1(n11909), .B2(n9203), .ZN(
        n6084) );
  INV_X1 U6635 ( .A(n6085), .ZN(n11908) );
  AOI22_X1 U6636 ( .A1(ram[1599]), .A2(n6070), .B1(n11909), .B2(n9227), .ZN(
        n6085) );
  INV_X1 U6637 ( .A(n6103), .ZN(n11859) );
  AOI22_X1 U6638 ( .A1(ram[1616]), .A2(n6104), .B1(n11875), .B2(n8866), .ZN(
        n6103) );
  INV_X1 U6639 ( .A(n6105), .ZN(n11860) );
  AOI22_X1 U6640 ( .A1(ram[1617]), .A2(n6104), .B1(n11875), .B2(n8890), .ZN(
        n6105) );
  INV_X1 U6641 ( .A(n6106), .ZN(n11861) );
  AOI22_X1 U6642 ( .A1(ram[1618]), .A2(n6104), .B1(n11875), .B2(n8914), .ZN(
        n6106) );
  INV_X1 U6643 ( .A(n6107), .ZN(n11862) );
  AOI22_X1 U6644 ( .A1(ram[1619]), .A2(n6104), .B1(n11875), .B2(n8938), .ZN(
        n6107) );
  INV_X1 U6645 ( .A(n6108), .ZN(n11863) );
  AOI22_X1 U6646 ( .A1(ram[1620]), .A2(n6104), .B1(n11875), .B2(n8962), .ZN(
        n6108) );
  INV_X1 U6647 ( .A(n6109), .ZN(n11864) );
  AOI22_X1 U6648 ( .A1(ram[1621]), .A2(n6104), .B1(n11875), .B2(n8986), .ZN(
        n6109) );
  INV_X1 U6649 ( .A(n6110), .ZN(n11865) );
  AOI22_X1 U6650 ( .A1(ram[1622]), .A2(n6104), .B1(n11875), .B2(n9010), .ZN(
        n6110) );
  INV_X1 U6651 ( .A(n6111), .ZN(n11866) );
  AOI22_X1 U6652 ( .A1(ram[1623]), .A2(n6104), .B1(n11875), .B2(n9034), .ZN(
        n6111) );
  INV_X1 U6653 ( .A(n6112), .ZN(n11867) );
  AOI22_X1 U6654 ( .A1(ram[1624]), .A2(n6104), .B1(n11875), .B2(n9058), .ZN(
        n6112) );
  INV_X1 U6655 ( .A(n6113), .ZN(n11868) );
  AOI22_X1 U6656 ( .A1(ram[1625]), .A2(n6104), .B1(n11875), .B2(n9082), .ZN(
        n6113) );
  INV_X1 U6657 ( .A(n6114), .ZN(n11869) );
  AOI22_X1 U6658 ( .A1(ram[1626]), .A2(n6104), .B1(n11875), .B2(n9106), .ZN(
        n6114) );
  INV_X1 U6659 ( .A(n6115), .ZN(n11870) );
  AOI22_X1 U6660 ( .A1(ram[1627]), .A2(n6104), .B1(n11875), .B2(n9130), .ZN(
        n6115) );
  INV_X1 U6661 ( .A(n6116), .ZN(n11871) );
  AOI22_X1 U6662 ( .A1(ram[1628]), .A2(n6104), .B1(n11875), .B2(n9154), .ZN(
        n6116) );
  INV_X1 U6663 ( .A(n6117), .ZN(n11872) );
  AOI22_X1 U6664 ( .A1(ram[1629]), .A2(n6104), .B1(n11875), .B2(n9178), .ZN(
        n6117) );
  INV_X1 U6665 ( .A(n6118), .ZN(n11873) );
  AOI22_X1 U6666 ( .A1(ram[1630]), .A2(n6104), .B1(n11875), .B2(n9202), .ZN(
        n6118) );
  INV_X1 U6667 ( .A(n6119), .ZN(n11874) );
  AOI22_X1 U6668 ( .A1(ram[1631]), .A2(n6104), .B1(n11875), .B2(n9226), .ZN(
        n6119) );
  INV_X1 U6669 ( .A(n6137), .ZN(n11825) );
  AOI22_X1 U6670 ( .A1(ram[1648]), .A2(n6138), .B1(n11841), .B2(n8866), .ZN(
        n6137) );
  INV_X1 U6671 ( .A(n6139), .ZN(n11826) );
  AOI22_X1 U6672 ( .A1(ram[1649]), .A2(n6138), .B1(n11841), .B2(n8890), .ZN(
        n6139) );
  INV_X1 U6673 ( .A(n6140), .ZN(n11827) );
  AOI22_X1 U6674 ( .A1(ram[1650]), .A2(n6138), .B1(n11841), .B2(n8914), .ZN(
        n6140) );
  INV_X1 U6675 ( .A(n6141), .ZN(n11828) );
  AOI22_X1 U6676 ( .A1(ram[1651]), .A2(n6138), .B1(n11841), .B2(n8938), .ZN(
        n6141) );
  INV_X1 U6677 ( .A(n6142), .ZN(n11829) );
  AOI22_X1 U6678 ( .A1(ram[1652]), .A2(n6138), .B1(n11841), .B2(n8962), .ZN(
        n6142) );
  INV_X1 U6679 ( .A(n6143), .ZN(n11830) );
  AOI22_X1 U6680 ( .A1(ram[1653]), .A2(n6138), .B1(n11841), .B2(n8986), .ZN(
        n6143) );
  INV_X1 U6681 ( .A(n6144), .ZN(n11831) );
  AOI22_X1 U6682 ( .A1(ram[1654]), .A2(n6138), .B1(n11841), .B2(n9010), .ZN(
        n6144) );
  INV_X1 U6683 ( .A(n6145), .ZN(n11832) );
  AOI22_X1 U6684 ( .A1(ram[1655]), .A2(n6138), .B1(n11841), .B2(n9034), .ZN(
        n6145) );
  INV_X1 U6685 ( .A(n6146), .ZN(n11833) );
  AOI22_X1 U6686 ( .A1(ram[1656]), .A2(n6138), .B1(n11841), .B2(n9058), .ZN(
        n6146) );
  INV_X1 U6687 ( .A(n6147), .ZN(n11834) );
  AOI22_X1 U6688 ( .A1(ram[1657]), .A2(n6138), .B1(n11841), .B2(n9082), .ZN(
        n6147) );
  INV_X1 U6689 ( .A(n6148), .ZN(n11835) );
  AOI22_X1 U6690 ( .A1(ram[1658]), .A2(n6138), .B1(n11841), .B2(n9106), .ZN(
        n6148) );
  INV_X1 U6691 ( .A(n6149), .ZN(n11836) );
  AOI22_X1 U6692 ( .A1(ram[1659]), .A2(n6138), .B1(n11841), .B2(n9130), .ZN(
        n6149) );
  INV_X1 U6693 ( .A(n6150), .ZN(n11837) );
  AOI22_X1 U6694 ( .A1(ram[1660]), .A2(n6138), .B1(n11841), .B2(n9154), .ZN(
        n6150) );
  INV_X1 U6695 ( .A(n6151), .ZN(n11838) );
  AOI22_X1 U6696 ( .A1(ram[1661]), .A2(n6138), .B1(n11841), .B2(n9178), .ZN(
        n6151) );
  INV_X1 U6697 ( .A(n6152), .ZN(n11839) );
  AOI22_X1 U6698 ( .A1(ram[1662]), .A2(n6138), .B1(n11841), .B2(n9202), .ZN(
        n6152) );
  INV_X1 U6699 ( .A(n6153), .ZN(n11840) );
  AOI22_X1 U6700 ( .A1(ram[1663]), .A2(n6138), .B1(n11841), .B2(n9226), .ZN(
        n6153) );
  INV_X1 U6701 ( .A(n6171), .ZN(n11791) );
  AOI22_X1 U6702 ( .A1(ram[1680]), .A2(n6172), .B1(n11807), .B2(n8866), .ZN(
        n6171) );
  INV_X1 U6703 ( .A(n6173), .ZN(n11792) );
  AOI22_X1 U6704 ( .A1(ram[1681]), .A2(n6172), .B1(n11807), .B2(n8890), .ZN(
        n6173) );
  INV_X1 U6705 ( .A(n6174), .ZN(n11793) );
  AOI22_X1 U6706 ( .A1(ram[1682]), .A2(n6172), .B1(n11807), .B2(n8914), .ZN(
        n6174) );
  INV_X1 U6707 ( .A(n6175), .ZN(n11794) );
  AOI22_X1 U6708 ( .A1(ram[1683]), .A2(n6172), .B1(n11807), .B2(n8938), .ZN(
        n6175) );
  INV_X1 U6709 ( .A(n6176), .ZN(n11795) );
  AOI22_X1 U6710 ( .A1(ram[1684]), .A2(n6172), .B1(n11807), .B2(n8962), .ZN(
        n6176) );
  INV_X1 U6711 ( .A(n6177), .ZN(n11796) );
  AOI22_X1 U6712 ( .A1(ram[1685]), .A2(n6172), .B1(n11807), .B2(n8986), .ZN(
        n6177) );
  INV_X1 U6713 ( .A(n6178), .ZN(n11797) );
  AOI22_X1 U6714 ( .A1(ram[1686]), .A2(n6172), .B1(n11807), .B2(n9010), .ZN(
        n6178) );
  INV_X1 U6715 ( .A(n6179), .ZN(n11798) );
  AOI22_X1 U6716 ( .A1(ram[1687]), .A2(n6172), .B1(n11807), .B2(n9034), .ZN(
        n6179) );
  INV_X1 U6717 ( .A(n6180), .ZN(n11799) );
  AOI22_X1 U6718 ( .A1(ram[1688]), .A2(n6172), .B1(n11807), .B2(n9058), .ZN(
        n6180) );
  INV_X1 U6719 ( .A(n6181), .ZN(n11800) );
  AOI22_X1 U6720 ( .A1(ram[1689]), .A2(n6172), .B1(n11807), .B2(n9082), .ZN(
        n6181) );
  INV_X1 U6721 ( .A(n6182), .ZN(n11801) );
  AOI22_X1 U6722 ( .A1(ram[1690]), .A2(n6172), .B1(n11807), .B2(n9106), .ZN(
        n6182) );
  INV_X1 U6723 ( .A(n6183), .ZN(n11802) );
  AOI22_X1 U6724 ( .A1(ram[1691]), .A2(n6172), .B1(n11807), .B2(n9130), .ZN(
        n6183) );
  INV_X1 U6725 ( .A(n6184), .ZN(n11803) );
  AOI22_X1 U6726 ( .A1(ram[1692]), .A2(n6172), .B1(n11807), .B2(n9154), .ZN(
        n6184) );
  INV_X1 U6727 ( .A(n6185), .ZN(n11804) );
  AOI22_X1 U6728 ( .A1(ram[1693]), .A2(n6172), .B1(n11807), .B2(n9178), .ZN(
        n6185) );
  INV_X1 U6729 ( .A(n6186), .ZN(n11805) );
  AOI22_X1 U6730 ( .A1(ram[1694]), .A2(n6172), .B1(n11807), .B2(n9202), .ZN(
        n6186) );
  INV_X1 U6731 ( .A(n6187), .ZN(n11806) );
  AOI22_X1 U6732 ( .A1(ram[1695]), .A2(n6172), .B1(n11807), .B2(n9226), .ZN(
        n6187) );
  INV_X1 U6733 ( .A(n6205), .ZN(n11757) );
  AOI22_X1 U6734 ( .A1(ram[1712]), .A2(n6206), .B1(n11773), .B2(n8866), .ZN(
        n6205) );
  INV_X1 U6735 ( .A(n6207), .ZN(n11758) );
  AOI22_X1 U6736 ( .A1(ram[1713]), .A2(n6206), .B1(n11773), .B2(n8890), .ZN(
        n6207) );
  INV_X1 U6737 ( .A(n6208), .ZN(n11759) );
  AOI22_X1 U6738 ( .A1(ram[1714]), .A2(n6206), .B1(n11773), .B2(n8914), .ZN(
        n6208) );
  INV_X1 U6739 ( .A(n6209), .ZN(n11760) );
  AOI22_X1 U6740 ( .A1(ram[1715]), .A2(n6206), .B1(n11773), .B2(n8938), .ZN(
        n6209) );
  INV_X1 U6741 ( .A(n6210), .ZN(n11761) );
  AOI22_X1 U6742 ( .A1(ram[1716]), .A2(n6206), .B1(n11773), .B2(n8962), .ZN(
        n6210) );
  INV_X1 U6743 ( .A(n6211), .ZN(n11762) );
  AOI22_X1 U6744 ( .A1(ram[1717]), .A2(n6206), .B1(n11773), .B2(n8986), .ZN(
        n6211) );
  INV_X1 U6745 ( .A(n6212), .ZN(n11763) );
  AOI22_X1 U6746 ( .A1(ram[1718]), .A2(n6206), .B1(n11773), .B2(n9010), .ZN(
        n6212) );
  INV_X1 U6747 ( .A(n6213), .ZN(n11764) );
  AOI22_X1 U6748 ( .A1(ram[1719]), .A2(n6206), .B1(n11773), .B2(n9034), .ZN(
        n6213) );
  INV_X1 U6749 ( .A(n6214), .ZN(n11765) );
  AOI22_X1 U6750 ( .A1(ram[1720]), .A2(n6206), .B1(n11773), .B2(n9058), .ZN(
        n6214) );
  INV_X1 U6751 ( .A(n6215), .ZN(n11766) );
  AOI22_X1 U6752 ( .A1(ram[1721]), .A2(n6206), .B1(n11773), .B2(n9082), .ZN(
        n6215) );
  INV_X1 U6753 ( .A(n6216), .ZN(n11767) );
  AOI22_X1 U6754 ( .A1(ram[1722]), .A2(n6206), .B1(n11773), .B2(n9106), .ZN(
        n6216) );
  INV_X1 U6755 ( .A(n6217), .ZN(n11768) );
  AOI22_X1 U6756 ( .A1(ram[1723]), .A2(n6206), .B1(n11773), .B2(n9130), .ZN(
        n6217) );
  INV_X1 U6757 ( .A(n6218), .ZN(n11769) );
  AOI22_X1 U6758 ( .A1(ram[1724]), .A2(n6206), .B1(n11773), .B2(n9154), .ZN(
        n6218) );
  INV_X1 U6759 ( .A(n6219), .ZN(n11770) );
  AOI22_X1 U6760 ( .A1(ram[1725]), .A2(n6206), .B1(n11773), .B2(n9178), .ZN(
        n6219) );
  INV_X1 U6761 ( .A(n6220), .ZN(n11771) );
  AOI22_X1 U6762 ( .A1(ram[1726]), .A2(n6206), .B1(n11773), .B2(n9202), .ZN(
        n6220) );
  INV_X1 U6763 ( .A(n6221), .ZN(n11772) );
  AOI22_X1 U6764 ( .A1(ram[1727]), .A2(n6206), .B1(n11773), .B2(n9226), .ZN(
        n6221) );
  INV_X1 U6765 ( .A(n6239), .ZN(n11723) );
  AOI22_X1 U6766 ( .A1(ram[1744]), .A2(n6240), .B1(n11739), .B2(n8866), .ZN(
        n6239) );
  INV_X1 U6767 ( .A(n6241), .ZN(n11724) );
  AOI22_X1 U6768 ( .A1(ram[1745]), .A2(n6240), .B1(n11739), .B2(n8890), .ZN(
        n6241) );
  INV_X1 U6769 ( .A(n6242), .ZN(n11725) );
  AOI22_X1 U6770 ( .A1(ram[1746]), .A2(n6240), .B1(n11739), .B2(n8914), .ZN(
        n6242) );
  INV_X1 U6771 ( .A(n6243), .ZN(n11726) );
  AOI22_X1 U6772 ( .A1(ram[1747]), .A2(n6240), .B1(n11739), .B2(n8938), .ZN(
        n6243) );
  INV_X1 U6773 ( .A(n6244), .ZN(n11727) );
  AOI22_X1 U6774 ( .A1(ram[1748]), .A2(n6240), .B1(n11739), .B2(n8962), .ZN(
        n6244) );
  INV_X1 U6775 ( .A(n6245), .ZN(n11728) );
  AOI22_X1 U6776 ( .A1(ram[1749]), .A2(n6240), .B1(n11739), .B2(n8986), .ZN(
        n6245) );
  INV_X1 U6777 ( .A(n6246), .ZN(n11729) );
  AOI22_X1 U6778 ( .A1(ram[1750]), .A2(n6240), .B1(n11739), .B2(n9010), .ZN(
        n6246) );
  INV_X1 U6779 ( .A(n6247), .ZN(n11730) );
  AOI22_X1 U6780 ( .A1(ram[1751]), .A2(n6240), .B1(n11739), .B2(n9034), .ZN(
        n6247) );
  INV_X1 U6781 ( .A(n6248), .ZN(n11731) );
  AOI22_X1 U6782 ( .A1(ram[1752]), .A2(n6240), .B1(n11739), .B2(n9058), .ZN(
        n6248) );
  INV_X1 U6783 ( .A(n6249), .ZN(n11732) );
  AOI22_X1 U6784 ( .A1(ram[1753]), .A2(n6240), .B1(n11739), .B2(n9082), .ZN(
        n6249) );
  INV_X1 U6785 ( .A(n6250), .ZN(n11733) );
  AOI22_X1 U6786 ( .A1(ram[1754]), .A2(n6240), .B1(n11739), .B2(n9106), .ZN(
        n6250) );
  INV_X1 U6787 ( .A(n6251), .ZN(n11734) );
  AOI22_X1 U6788 ( .A1(ram[1755]), .A2(n6240), .B1(n11739), .B2(n9130), .ZN(
        n6251) );
  INV_X1 U6789 ( .A(n6252), .ZN(n11735) );
  AOI22_X1 U6790 ( .A1(ram[1756]), .A2(n6240), .B1(n11739), .B2(n9154), .ZN(
        n6252) );
  INV_X1 U6791 ( .A(n6253), .ZN(n11736) );
  AOI22_X1 U6792 ( .A1(ram[1757]), .A2(n6240), .B1(n11739), .B2(n9178), .ZN(
        n6253) );
  INV_X1 U6793 ( .A(n6254), .ZN(n11737) );
  AOI22_X1 U6794 ( .A1(ram[1758]), .A2(n6240), .B1(n11739), .B2(n9202), .ZN(
        n6254) );
  INV_X1 U6795 ( .A(n6255), .ZN(n11738) );
  AOI22_X1 U6796 ( .A1(ram[1759]), .A2(n6240), .B1(n11739), .B2(n9226), .ZN(
        n6255) );
  INV_X1 U6797 ( .A(n6273), .ZN(n11689) );
  AOI22_X1 U6798 ( .A1(ram[1776]), .A2(n6274), .B1(n11705), .B2(n8866), .ZN(
        n6273) );
  INV_X1 U6799 ( .A(n6275), .ZN(n11690) );
  AOI22_X1 U6800 ( .A1(ram[1777]), .A2(n6274), .B1(n11705), .B2(n8890), .ZN(
        n6275) );
  INV_X1 U6801 ( .A(n6276), .ZN(n11691) );
  AOI22_X1 U6802 ( .A1(ram[1778]), .A2(n6274), .B1(n11705), .B2(n8914), .ZN(
        n6276) );
  INV_X1 U6803 ( .A(n6277), .ZN(n11692) );
  AOI22_X1 U6804 ( .A1(ram[1779]), .A2(n6274), .B1(n11705), .B2(n8938), .ZN(
        n6277) );
  INV_X1 U6805 ( .A(n6278), .ZN(n11693) );
  AOI22_X1 U6806 ( .A1(ram[1780]), .A2(n6274), .B1(n11705), .B2(n8962), .ZN(
        n6278) );
  INV_X1 U6807 ( .A(n6279), .ZN(n11694) );
  AOI22_X1 U6808 ( .A1(ram[1781]), .A2(n6274), .B1(n11705), .B2(n8986), .ZN(
        n6279) );
  INV_X1 U6809 ( .A(n6280), .ZN(n11695) );
  AOI22_X1 U6810 ( .A1(ram[1782]), .A2(n6274), .B1(n11705), .B2(n9010), .ZN(
        n6280) );
  INV_X1 U6811 ( .A(n6281), .ZN(n11696) );
  AOI22_X1 U6812 ( .A1(ram[1783]), .A2(n6274), .B1(n11705), .B2(n9034), .ZN(
        n6281) );
  INV_X1 U6813 ( .A(n6282), .ZN(n11697) );
  AOI22_X1 U6814 ( .A1(ram[1784]), .A2(n6274), .B1(n11705), .B2(n9058), .ZN(
        n6282) );
  INV_X1 U6815 ( .A(n6283), .ZN(n11698) );
  AOI22_X1 U6816 ( .A1(ram[1785]), .A2(n6274), .B1(n11705), .B2(n9082), .ZN(
        n6283) );
  INV_X1 U6817 ( .A(n6284), .ZN(n11699) );
  AOI22_X1 U6818 ( .A1(ram[1786]), .A2(n6274), .B1(n11705), .B2(n9106), .ZN(
        n6284) );
  INV_X1 U6819 ( .A(n6285), .ZN(n11700) );
  AOI22_X1 U6820 ( .A1(ram[1787]), .A2(n6274), .B1(n11705), .B2(n9130), .ZN(
        n6285) );
  INV_X1 U6821 ( .A(n6286), .ZN(n11701) );
  AOI22_X1 U6822 ( .A1(ram[1788]), .A2(n6274), .B1(n11705), .B2(n9154), .ZN(
        n6286) );
  INV_X1 U6823 ( .A(n6287), .ZN(n11702) );
  AOI22_X1 U6824 ( .A1(ram[1789]), .A2(n6274), .B1(n11705), .B2(n9178), .ZN(
        n6287) );
  INV_X1 U6825 ( .A(n6288), .ZN(n11703) );
  AOI22_X1 U6826 ( .A1(ram[1790]), .A2(n6274), .B1(n11705), .B2(n9202), .ZN(
        n6288) );
  INV_X1 U6827 ( .A(n6289), .ZN(n11704) );
  AOI22_X1 U6828 ( .A1(ram[1791]), .A2(n6274), .B1(n11705), .B2(n9226), .ZN(
        n6289) );
  INV_X1 U6829 ( .A(n6308), .ZN(n11655) );
  AOI22_X1 U6830 ( .A1(ram[1808]), .A2(n6309), .B1(n11671), .B2(n8865), .ZN(
        n6308) );
  INV_X1 U6831 ( .A(n6310), .ZN(n11656) );
  AOI22_X1 U6832 ( .A1(ram[1809]), .A2(n6309), .B1(n11671), .B2(n8889), .ZN(
        n6310) );
  INV_X1 U6833 ( .A(n6311), .ZN(n11657) );
  AOI22_X1 U6834 ( .A1(ram[1810]), .A2(n6309), .B1(n11671), .B2(n8913), .ZN(
        n6311) );
  INV_X1 U6835 ( .A(n6312), .ZN(n11658) );
  AOI22_X1 U6836 ( .A1(ram[1811]), .A2(n6309), .B1(n11671), .B2(n8937), .ZN(
        n6312) );
  INV_X1 U6837 ( .A(n6313), .ZN(n11659) );
  AOI22_X1 U6838 ( .A1(ram[1812]), .A2(n6309), .B1(n11671), .B2(n8961), .ZN(
        n6313) );
  INV_X1 U6839 ( .A(n6314), .ZN(n11660) );
  AOI22_X1 U6840 ( .A1(ram[1813]), .A2(n6309), .B1(n11671), .B2(n8985), .ZN(
        n6314) );
  INV_X1 U6841 ( .A(n6315), .ZN(n11661) );
  AOI22_X1 U6842 ( .A1(ram[1814]), .A2(n6309), .B1(n11671), .B2(n9009), .ZN(
        n6315) );
  INV_X1 U6843 ( .A(n6316), .ZN(n11662) );
  AOI22_X1 U6844 ( .A1(ram[1815]), .A2(n6309), .B1(n11671), .B2(n9033), .ZN(
        n6316) );
  INV_X1 U6845 ( .A(n6317), .ZN(n11663) );
  AOI22_X1 U6846 ( .A1(ram[1816]), .A2(n6309), .B1(n11671), .B2(n9057), .ZN(
        n6317) );
  INV_X1 U6847 ( .A(n6318), .ZN(n11664) );
  AOI22_X1 U6848 ( .A1(ram[1817]), .A2(n6309), .B1(n11671), .B2(n9081), .ZN(
        n6318) );
  INV_X1 U6849 ( .A(n6319), .ZN(n11665) );
  AOI22_X1 U6850 ( .A1(ram[1818]), .A2(n6309), .B1(n11671), .B2(n9105), .ZN(
        n6319) );
  INV_X1 U6851 ( .A(n6320), .ZN(n11666) );
  AOI22_X1 U6852 ( .A1(ram[1819]), .A2(n6309), .B1(n11671), .B2(n9129), .ZN(
        n6320) );
  INV_X1 U6853 ( .A(n6321), .ZN(n11667) );
  AOI22_X1 U6854 ( .A1(ram[1820]), .A2(n6309), .B1(n11671), .B2(n9153), .ZN(
        n6321) );
  INV_X1 U6855 ( .A(n6322), .ZN(n11668) );
  AOI22_X1 U6856 ( .A1(ram[1821]), .A2(n6309), .B1(n11671), .B2(n9177), .ZN(
        n6322) );
  INV_X1 U6857 ( .A(n6323), .ZN(n11669) );
  AOI22_X1 U6858 ( .A1(ram[1822]), .A2(n6309), .B1(n11671), .B2(n9201), .ZN(
        n6323) );
  INV_X1 U6859 ( .A(n6324), .ZN(n11670) );
  AOI22_X1 U6860 ( .A1(ram[1823]), .A2(n6309), .B1(n11671), .B2(n9225), .ZN(
        n6324) );
  INV_X1 U6861 ( .A(n6342), .ZN(n11621) );
  AOI22_X1 U6862 ( .A1(ram[1840]), .A2(n6343), .B1(n11637), .B2(n8865), .ZN(
        n6342) );
  INV_X1 U6863 ( .A(n6344), .ZN(n11622) );
  AOI22_X1 U6864 ( .A1(ram[1841]), .A2(n6343), .B1(n11637), .B2(n8889), .ZN(
        n6344) );
  INV_X1 U6865 ( .A(n6345), .ZN(n11623) );
  AOI22_X1 U6866 ( .A1(ram[1842]), .A2(n6343), .B1(n11637), .B2(n8913), .ZN(
        n6345) );
  INV_X1 U6867 ( .A(n6346), .ZN(n11624) );
  AOI22_X1 U6868 ( .A1(ram[1843]), .A2(n6343), .B1(n11637), .B2(n8937), .ZN(
        n6346) );
  INV_X1 U6869 ( .A(n6347), .ZN(n11625) );
  AOI22_X1 U6870 ( .A1(ram[1844]), .A2(n6343), .B1(n11637), .B2(n8961), .ZN(
        n6347) );
  INV_X1 U6871 ( .A(n6348), .ZN(n11626) );
  AOI22_X1 U6872 ( .A1(ram[1845]), .A2(n6343), .B1(n11637), .B2(n8985), .ZN(
        n6348) );
  INV_X1 U6873 ( .A(n6349), .ZN(n11627) );
  AOI22_X1 U6874 ( .A1(ram[1846]), .A2(n6343), .B1(n11637), .B2(n9009), .ZN(
        n6349) );
  INV_X1 U6875 ( .A(n6350), .ZN(n11628) );
  AOI22_X1 U6876 ( .A1(ram[1847]), .A2(n6343), .B1(n11637), .B2(n9033), .ZN(
        n6350) );
  INV_X1 U6877 ( .A(n6351), .ZN(n11629) );
  AOI22_X1 U6878 ( .A1(ram[1848]), .A2(n6343), .B1(n11637), .B2(n9057), .ZN(
        n6351) );
  INV_X1 U6879 ( .A(n6352), .ZN(n11630) );
  AOI22_X1 U6880 ( .A1(ram[1849]), .A2(n6343), .B1(n11637), .B2(n9081), .ZN(
        n6352) );
  INV_X1 U6881 ( .A(n6353), .ZN(n11631) );
  AOI22_X1 U6882 ( .A1(ram[1850]), .A2(n6343), .B1(n11637), .B2(n9105), .ZN(
        n6353) );
  INV_X1 U6883 ( .A(n6354), .ZN(n11632) );
  AOI22_X1 U6884 ( .A1(ram[1851]), .A2(n6343), .B1(n11637), .B2(n9129), .ZN(
        n6354) );
  INV_X1 U6885 ( .A(n6355), .ZN(n11633) );
  AOI22_X1 U6886 ( .A1(ram[1852]), .A2(n6343), .B1(n11637), .B2(n9153), .ZN(
        n6355) );
  INV_X1 U6887 ( .A(n6356), .ZN(n11634) );
  AOI22_X1 U6888 ( .A1(ram[1853]), .A2(n6343), .B1(n11637), .B2(n9177), .ZN(
        n6356) );
  INV_X1 U6889 ( .A(n6357), .ZN(n11635) );
  AOI22_X1 U6890 ( .A1(ram[1854]), .A2(n6343), .B1(n11637), .B2(n9201), .ZN(
        n6357) );
  INV_X1 U6891 ( .A(n6358), .ZN(n11636) );
  AOI22_X1 U6892 ( .A1(ram[1855]), .A2(n6343), .B1(n11637), .B2(n9225), .ZN(
        n6358) );
  INV_X1 U6893 ( .A(n6376), .ZN(n11587) );
  AOI22_X1 U6894 ( .A1(ram[1872]), .A2(n6377), .B1(n11603), .B2(n8865), .ZN(
        n6376) );
  INV_X1 U6895 ( .A(n6378), .ZN(n11588) );
  AOI22_X1 U6896 ( .A1(ram[1873]), .A2(n6377), .B1(n11603), .B2(n8889), .ZN(
        n6378) );
  INV_X1 U6897 ( .A(n6379), .ZN(n11589) );
  AOI22_X1 U6898 ( .A1(ram[1874]), .A2(n6377), .B1(n11603), .B2(n8913), .ZN(
        n6379) );
  INV_X1 U6899 ( .A(n6380), .ZN(n11590) );
  AOI22_X1 U6900 ( .A1(ram[1875]), .A2(n6377), .B1(n11603), .B2(n8937), .ZN(
        n6380) );
  INV_X1 U6901 ( .A(n6381), .ZN(n11591) );
  AOI22_X1 U6902 ( .A1(ram[1876]), .A2(n6377), .B1(n11603), .B2(n8961), .ZN(
        n6381) );
  INV_X1 U6903 ( .A(n6382), .ZN(n11592) );
  AOI22_X1 U6904 ( .A1(ram[1877]), .A2(n6377), .B1(n11603), .B2(n8985), .ZN(
        n6382) );
  INV_X1 U6905 ( .A(n6383), .ZN(n11593) );
  AOI22_X1 U6906 ( .A1(ram[1878]), .A2(n6377), .B1(n11603), .B2(n9009), .ZN(
        n6383) );
  INV_X1 U6907 ( .A(n6384), .ZN(n11594) );
  AOI22_X1 U6908 ( .A1(ram[1879]), .A2(n6377), .B1(n11603), .B2(n9033), .ZN(
        n6384) );
  INV_X1 U6909 ( .A(n6385), .ZN(n11595) );
  AOI22_X1 U6910 ( .A1(ram[1880]), .A2(n6377), .B1(n11603), .B2(n9057), .ZN(
        n6385) );
  INV_X1 U6911 ( .A(n6386), .ZN(n11596) );
  AOI22_X1 U6912 ( .A1(ram[1881]), .A2(n6377), .B1(n11603), .B2(n9081), .ZN(
        n6386) );
  INV_X1 U6913 ( .A(n6387), .ZN(n11597) );
  AOI22_X1 U6914 ( .A1(ram[1882]), .A2(n6377), .B1(n11603), .B2(n9105), .ZN(
        n6387) );
  INV_X1 U6915 ( .A(n6388), .ZN(n11598) );
  AOI22_X1 U6916 ( .A1(ram[1883]), .A2(n6377), .B1(n11603), .B2(n9129), .ZN(
        n6388) );
  INV_X1 U6917 ( .A(n6389), .ZN(n11599) );
  AOI22_X1 U6918 ( .A1(ram[1884]), .A2(n6377), .B1(n11603), .B2(n9153), .ZN(
        n6389) );
  INV_X1 U6919 ( .A(n6390), .ZN(n11600) );
  AOI22_X1 U6920 ( .A1(ram[1885]), .A2(n6377), .B1(n11603), .B2(n9177), .ZN(
        n6390) );
  INV_X1 U6921 ( .A(n6391), .ZN(n11601) );
  AOI22_X1 U6922 ( .A1(ram[1886]), .A2(n6377), .B1(n11603), .B2(n9201), .ZN(
        n6391) );
  INV_X1 U6923 ( .A(n6392), .ZN(n11602) );
  AOI22_X1 U6924 ( .A1(ram[1887]), .A2(n6377), .B1(n11603), .B2(n9225), .ZN(
        n6392) );
  INV_X1 U6925 ( .A(n6410), .ZN(n11553) );
  AOI22_X1 U6926 ( .A1(ram[1904]), .A2(n6411), .B1(n11569), .B2(n8865), .ZN(
        n6410) );
  INV_X1 U6927 ( .A(n6412), .ZN(n11554) );
  AOI22_X1 U6928 ( .A1(ram[1905]), .A2(n6411), .B1(n11569), .B2(n8889), .ZN(
        n6412) );
  INV_X1 U6929 ( .A(n6413), .ZN(n11555) );
  AOI22_X1 U6930 ( .A1(ram[1906]), .A2(n6411), .B1(n11569), .B2(n8913), .ZN(
        n6413) );
  INV_X1 U6931 ( .A(n6414), .ZN(n11556) );
  AOI22_X1 U6932 ( .A1(ram[1907]), .A2(n6411), .B1(n11569), .B2(n8937), .ZN(
        n6414) );
  INV_X1 U6933 ( .A(n6415), .ZN(n11557) );
  AOI22_X1 U6934 ( .A1(ram[1908]), .A2(n6411), .B1(n11569), .B2(n8961), .ZN(
        n6415) );
  INV_X1 U6935 ( .A(n6416), .ZN(n11558) );
  AOI22_X1 U6936 ( .A1(ram[1909]), .A2(n6411), .B1(n11569), .B2(n8985), .ZN(
        n6416) );
  INV_X1 U6937 ( .A(n6417), .ZN(n11559) );
  AOI22_X1 U6938 ( .A1(ram[1910]), .A2(n6411), .B1(n11569), .B2(n9009), .ZN(
        n6417) );
  INV_X1 U6939 ( .A(n6418), .ZN(n11560) );
  AOI22_X1 U6940 ( .A1(ram[1911]), .A2(n6411), .B1(n11569), .B2(n9033), .ZN(
        n6418) );
  INV_X1 U6941 ( .A(n6419), .ZN(n11561) );
  AOI22_X1 U6942 ( .A1(ram[1912]), .A2(n6411), .B1(n11569), .B2(n9057), .ZN(
        n6419) );
  INV_X1 U6943 ( .A(n6420), .ZN(n11562) );
  AOI22_X1 U6944 ( .A1(ram[1913]), .A2(n6411), .B1(n11569), .B2(n9081), .ZN(
        n6420) );
  INV_X1 U6945 ( .A(n6421), .ZN(n11563) );
  AOI22_X1 U6946 ( .A1(ram[1914]), .A2(n6411), .B1(n11569), .B2(n9105), .ZN(
        n6421) );
  INV_X1 U6947 ( .A(n6422), .ZN(n11564) );
  AOI22_X1 U6948 ( .A1(ram[1915]), .A2(n6411), .B1(n11569), .B2(n9129), .ZN(
        n6422) );
  INV_X1 U6949 ( .A(n6423), .ZN(n11565) );
  AOI22_X1 U6950 ( .A1(ram[1916]), .A2(n6411), .B1(n11569), .B2(n9153), .ZN(
        n6423) );
  INV_X1 U6951 ( .A(n6424), .ZN(n11566) );
  AOI22_X1 U6952 ( .A1(ram[1917]), .A2(n6411), .B1(n11569), .B2(n9177), .ZN(
        n6424) );
  INV_X1 U6953 ( .A(n6425), .ZN(n11567) );
  AOI22_X1 U6954 ( .A1(ram[1918]), .A2(n6411), .B1(n11569), .B2(n9201), .ZN(
        n6425) );
  INV_X1 U6955 ( .A(n6426), .ZN(n11568) );
  AOI22_X1 U6956 ( .A1(ram[1919]), .A2(n6411), .B1(n11569), .B2(n9225), .ZN(
        n6426) );
  INV_X1 U6957 ( .A(n6444), .ZN(n11519) );
  AOI22_X1 U6958 ( .A1(ram[1936]), .A2(n6445), .B1(n11535), .B2(n8865), .ZN(
        n6444) );
  INV_X1 U6959 ( .A(n6446), .ZN(n11520) );
  AOI22_X1 U6960 ( .A1(ram[1937]), .A2(n6445), .B1(n11535), .B2(n8889), .ZN(
        n6446) );
  INV_X1 U6961 ( .A(n6447), .ZN(n11521) );
  AOI22_X1 U6962 ( .A1(ram[1938]), .A2(n6445), .B1(n11535), .B2(n8913), .ZN(
        n6447) );
  INV_X1 U6963 ( .A(n6448), .ZN(n11522) );
  AOI22_X1 U6964 ( .A1(ram[1939]), .A2(n6445), .B1(n11535), .B2(n8937), .ZN(
        n6448) );
  INV_X1 U6965 ( .A(n6449), .ZN(n11523) );
  AOI22_X1 U6966 ( .A1(ram[1940]), .A2(n6445), .B1(n11535), .B2(n8961), .ZN(
        n6449) );
  INV_X1 U6967 ( .A(n6450), .ZN(n11524) );
  AOI22_X1 U6968 ( .A1(ram[1941]), .A2(n6445), .B1(n11535), .B2(n8985), .ZN(
        n6450) );
  INV_X1 U6969 ( .A(n6451), .ZN(n11525) );
  AOI22_X1 U6970 ( .A1(ram[1942]), .A2(n6445), .B1(n11535), .B2(n9009), .ZN(
        n6451) );
  INV_X1 U6971 ( .A(n6452), .ZN(n11526) );
  AOI22_X1 U6972 ( .A1(ram[1943]), .A2(n6445), .B1(n11535), .B2(n9033), .ZN(
        n6452) );
  INV_X1 U6973 ( .A(n6453), .ZN(n11527) );
  AOI22_X1 U6974 ( .A1(ram[1944]), .A2(n6445), .B1(n11535), .B2(n9057), .ZN(
        n6453) );
  INV_X1 U6975 ( .A(n6454), .ZN(n11528) );
  AOI22_X1 U6976 ( .A1(ram[1945]), .A2(n6445), .B1(n11535), .B2(n9081), .ZN(
        n6454) );
  INV_X1 U6977 ( .A(n6455), .ZN(n11529) );
  AOI22_X1 U6978 ( .A1(ram[1946]), .A2(n6445), .B1(n11535), .B2(n9105), .ZN(
        n6455) );
  INV_X1 U6979 ( .A(n6456), .ZN(n11530) );
  AOI22_X1 U6980 ( .A1(ram[1947]), .A2(n6445), .B1(n11535), .B2(n9129), .ZN(
        n6456) );
  INV_X1 U6981 ( .A(n6457), .ZN(n11531) );
  AOI22_X1 U6982 ( .A1(ram[1948]), .A2(n6445), .B1(n11535), .B2(n9153), .ZN(
        n6457) );
  INV_X1 U6983 ( .A(n6458), .ZN(n11532) );
  AOI22_X1 U6984 ( .A1(ram[1949]), .A2(n6445), .B1(n11535), .B2(n9177), .ZN(
        n6458) );
  INV_X1 U6985 ( .A(n6459), .ZN(n11533) );
  AOI22_X1 U6986 ( .A1(ram[1950]), .A2(n6445), .B1(n11535), .B2(n9201), .ZN(
        n6459) );
  INV_X1 U6987 ( .A(n6460), .ZN(n11534) );
  AOI22_X1 U6988 ( .A1(ram[1951]), .A2(n6445), .B1(n11535), .B2(n9225), .ZN(
        n6460) );
  INV_X1 U6989 ( .A(n6478), .ZN(n11485) );
  AOI22_X1 U6990 ( .A1(ram[1968]), .A2(n6479), .B1(n11501), .B2(n8865), .ZN(
        n6478) );
  INV_X1 U6991 ( .A(n6480), .ZN(n11486) );
  AOI22_X1 U6992 ( .A1(ram[1969]), .A2(n6479), .B1(n11501), .B2(n8889), .ZN(
        n6480) );
  INV_X1 U6993 ( .A(n6481), .ZN(n11487) );
  AOI22_X1 U6994 ( .A1(ram[1970]), .A2(n6479), .B1(n11501), .B2(n8913), .ZN(
        n6481) );
  INV_X1 U6995 ( .A(n6482), .ZN(n11488) );
  AOI22_X1 U6996 ( .A1(ram[1971]), .A2(n6479), .B1(n11501), .B2(n8937), .ZN(
        n6482) );
  INV_X1 U6997 ( .A(n6483), .ZN(n11489) );
  AOI22_X1 U6998 ( .A1(ram[1972]), .A2(n6479), .B1(n11501), .B2(n8961), .ZN(
        n6483) );
  INV_X1 U6999 ( .A(n6484), .ZN(n11490) );
  AOI22_X1 U7000 ( .A1(ram[1973]), .A2(n6479), .B1(n11501), .B2(n8985), .ZN(
        n6484) );
  INV_X1 U7001 ( .A(n6485), .ZN(n11491) );
  AOI22_X1 U7002 ( .A1(ram[1974]), .A2(n6479), .B1(n11501), .B2(n9009), .ZN(
        n6485) );
  INV_X1 U7003 ( .A(n6486), .ZN(n11492) );
  AOI22_X1 U7004 ( .A1(ram[1975]), .A2(n6479), .B1(n11501), .B2(n9033), .ZN(
        n6486) );
  INV_X1 U7005 ( .A(n6487), .ZN(n11493) );
  AOI22_X1 U7006 ( .A1(ram[1976]), .A2(n6479), .B1(n11501), .B2(n9057), .ZN(
        n6487) );
  INV_X1 U7007 ( .A(n6488), .ZN(n11494) );
  AOI22_X1 U7008 ( .A1(ram[1977]), .A2(n6479), .B1(n11501), .B2(n9081), .ZN(
        n6488) );
  INV_X1 U7009 ( .A(n6489), .ZN(n11495) );
  AOI22_X1 U7010 ( .A1(ram[1978]), .A2(n6479), .B1(n11501), .B2(n9105), .ZN(
        n6489) );
  INV_X1 U7011 ( .A(n6490), .ZN(n11496) );
  AOI22_X1 U7012 ( .A1(ram[1979]), .A2(n6479), .B1(n11501), .B2(n9129), .ZN(
        n6490) );
  INV_X1 U7013 ( .A(n6491), .ZN(n11497) );
  AOI22_X1 U7014 ( .A1(ram[1980]), .A2(n6479), .B1(n11501), .B2(n9153), .ZN(
        n6491) );
  INV_X1 U7015 ( .A(n6492), .ZN(n11498) );
  AOI22_X1 U7016 ( .A1(ram[1981]), .A2(n6479), .B1(n11501), .B2(n9177), .ZN(
        n6492) );
  INV_X1 U7017 ( .A(n6493), .ZN(n11499) );
  AOI22_X1 U7018 ( .A1(ram[1982]), .A2(n6479), .B1(n11501), .B2(n9201), .ZN(
        n6493) );
  INV_X1 U7019 ( .A(n6494), .ZN(n11500) );
  AOI22_X1 U7020 ( .A1(ram[1983]), .A2(n6479), .B1(n11501), .B2(n9225), .ZN(
        n6494) );
  INV_X1 U7021 ( .A(n6512), .ZN(n11451) );
  AOI22_X1 U7022 ( .A1(ram[2000]), .A2(n6513), .B1(n11467), .B2(n8864), .ZN(
        n6512) );
  INV_X1 U7023 ( .A(n6514), .ZN(n11452) );
  AOI22_X1 U7024 ( .A1(ram[2001]), .A2(n6513), .B1(n11467), .B2(n8888), .ZN(
        n6514) );
  INV_X1 U7025 ( .A(n6515), .ZN(n11453) );
  AOI22_X1 U7026 ( .A1(ram[2002]), .A2(n6513), .B1(n11467), .B2(n8912), .ZN(
        n6515) );
  INV_X1 U7027 ( .A(n6516), .ZN(n11454) );
  AOI22_X1 U7028 ( .A1(ram[2003]), .A2(n6513), .B1(n11467), .B2(n8936), .ZN(
        n6516) );
  INV_X1 U7029 ( .A(n6517), .ZN(n11455) );
  AOI22_X1 U7030 ( .A1(ram[2004]), .A2(n6513), .B1(n11467), .B2(n8960), .ZN(
        n6517) );
  INV_X1 U7031 ( .A(n6518), .ZN(n11456) );
  AOI22_X1 U7032 ( .A1(ram[2005]), .A2(n6513), .B1(n11467), .B2(n8984), .ZN(
        n6518) );
  INV_X1 U7033 ( .A(n6519), .ZN(n11457) );
  AOI22_X1 U7034 ( .A1(ram[2006]), .A2(n6513), .B1(n11467), .B2(n9008), .ZN(
        n6519) );
  INV_X1 U7035 ( .A(n6520), .ZN(n11458) );
  AOI22_X1 U7036 ( .A1(ram[2007]), .A2(n6513), .B1(n11467), .B2(n9032), .ZN(
        n6520) );
  INV_X1 U7037 ( .A(n6521), .ZN(n11459) );
  AOI22_X1 U7038 ( .A1(ram[2008]), .A2(n6513), .B1(n11467), .B2(n9056), .ZN(
        n6521) );
  INV_X1 U7039 ( .A(n6522), .ZN(n11460) );
  AOI22_X1 U7040 ( .A1(ram[2009]), .A2(n6513), .B1(n11467), .B2(n9080), .ZN(
        n6522) );
  INV_X1 U7041 ( .A(n6523), .ZN(n11461) );
  AOI22_X1 U7042 ( .A1(ram[2010]), .A2(n6513), .B1(n11467), .B2(n9104), .ZN(
        n6523) );
  INV_X1 U7043 ( .A(n6524), .ZN(n11462) );
  AOI22_X1 U7044 ( .A1(ram[2011]), .A2(n6513), .B1(n11467), .B2(n9128), .ZN(
        n6524) );
  INV_X1 U7045 ( .A(n6525), .ZN(n11463) );
  AOI22_X1 U7046 ( .A1(ram[2012]), .A2(n6513), .B1(n11467), .B2(n9152), .ZN(
        n6525) );
  INV_X1 U7047 ( .A(n6526), .ZN(n11464) );
  AOI22_X1 U7048 ( .A1(ram[2013]), .A2(n6513), .B1(n11467), .B2(n9176), .ZN(
        n6526) );
  INV_X1 U7049 ( .A(n6527), .ZN(n11465) );
  AOI22_X1 U7050 ( .A1(ram[2014]), .A2(n6513), .B1(n11467), .B2(n9200), .ZN(
        n6527) );
  INV_X1 U7051 ( .A(n6528), .ZN(n11466) );
  AOI22_X1 U7052 ( .A1(ram[2015]), .A2(n6513), .B1(n11467), .B2(n9224), .ZN(
        n6528) );
  INV_X1 U7053 ( .A(n6546), .ZN(n11417) );
  AOI22_X1 U7054 ( .A1(ram[2032]), .A2(n6547), .B1(n11433), .B2(n8864), .ZN(
        n6546) );
  INV_X1 U7055 ( .A(n6548), .ZN(n11418) );
  AOI22_X1 U7056 ( .A1(ram[2033]), .A2(n6547), .B1(n11433), .B2(n8888), .ZN(
        n6548) );
  INV_X1 U7057 ( .A(n6549), .ZN(n11419) );
  AOI22_X1 U7058 ( .A1(ram[2034]), .A2(n6547), .B1(n11433), .B2(n8912), .ZN(
        n6549) );
  INV_X1 U7059 ( .A(n6550), .ZN(n11420) );
  AOI22_X1 U7060 ( .A1(ram[2035]), .A2(n6547), .B1(n11433), .B2(n8936), .ZN(
        n6550) );
  INV_X1 U7061 ( .A(n6551), .ZN(n11421) );
  AOI22_X1 U7062 ( .A1(ram[2036]), .A2(n6547), .B1(n11433), .B2(n8960), .ZN(
        n6551) );
  INV_X1 U7063 ( .A(n6552), .ZN(n11422) );
  AOI22_X1 U7064 ( .A1(ram[2037]), .A2(n6547), .B1(n11433), .B2(n8984), .ZN(
        n6552) );
  INV_X1 U7065 ( .A(n6553), .ZN(n11423) );
  AOI22_X1 U7066 ( .A1(ram[2038]), .A2(n6547), .B1(n11433), .B2(n9008), .ZN(
        n6553) );
  INV_X1 U7067 ( .A(n6554), .ZN(n11424) );
  AOI22_X1 U7068 ( .A1(ram[2039]), .A2(n6547), .B1(n11433), .B2(n9032), .ZN(
        n6554) );
  INV_X1 U7069 ( .A(n6555), .ZN(n11425) );
  AOI22_X1 U7070 ( .A1(ram[2040]), .A2(n6547), .B1(n11433), .B2(n9056), .ZN(
        n6555) );
  INV_X1 U7071 ( .A(n6556), .ZN(n11426) );
  AOI22_X1 U7072 ( .A1(ram[2041]), .A2(n6547), .B1(n11433), .B2(n9080), .ZN(
        n6556) );
  INV_X1 U7073 ( .A(n6557), .ZN(n11427) );
  AOI22_X1 U7074 ( .A1(ram[2042]), .A2(n6547), .B1(n11433), .B2(n9104), .ZN(
        n6557) );
  INV_X1 U7075 ( .A(n6558), .ZN(n11428) );
  AOI22_X1 U7076 ( .A1(ram[2043]), .A2(n6547), .B1(n11433), .B2(n9128), .ZN(
        n6558) );
  INV_X1 U7077 ( .A(n6559), .ZN(n11429) );
  AOI22_X1 U7078 ( .A1(ram[2044]), .A2(n6547), .B1(n11433), .B2(n9152), .ZN(
        n6559) );
  INV_X1 U7079 ( .A(n6560), .ZN(n11430) );
  AOI22_X1 U7080 ( .A1(ram[2045]), .A2(n6547), .B1(n11433), .B2(n9176), .ZN(
        n6560) );
  INV_X1 U7081 ( .A(n6561), .ZN(n11431) );
  AOI22_X1 U7082 ( .A1(ram[2046]), .A2(n6547), .B1(n11433), .B2(n9200), .ZN(
        n6561) );
  INV_X1 U7083 ( .A(n6562), .ZN(n11432) );
  AOI22_X1 U7084 ( .A1(ram[2047]), .A2(n6547), .B1(n11433), .B2(n9224), .ZN(
        n6562) );
  INV_X1 U7085 ( .A(n6581), .ZN(n11383) );
  AOI22_X1 U7086 ( .A1(ram[2064]), .A2(n6582), .B1(n11399), .B2(n8864), .ZN(
        n6581) );
  INV_X1 U7087 ( .A(n6583), .ZN(n11384) );
  AOI22_X1 U7088 ( .A1(ram[2065]), .A2(n6582), .B1(n11399), .B2(n8888), .ZN(
        n6583) );
  INV_X1 U7089 ( .A(n6584), .ZN(n11385) );
  AOI22_X1 U7090 ( .A1(ram[2066]), .A2(n6582), .B1(n11399), .B2(n8912), .ZN(
        n6584) );
  INV_X1 U7091 ( .A(n6585), .ZN(n11386) );
  AOI22_X1 U7092 ( .A1(ram[2067]), .A2(n6582), .B1(n11399), .B2(n8936), .ZN(
        n6585) );
  INV_X1 U7093 ( .A(n6586), .ZN(n11387) );
  AOI22_X1 U7094 ( .A1(ram[2068]), .A2(n6582), .B1(n11399), .B2(n8960), .ZN(
        n6586) );
  INV_X1 U7095 ( .A(n6587), .ZN(n11388) );
  AOI22_X1 U7096 ( .A1(ram[2069]), .A2(n6582), .B1(n11399), .B2(n8984), .ZN(
        n6587) );
  INV_X1 U7097 ( .A(n6588), .ZN(n11389) );
  AOI22_X1 U7098 ( .A1(ram[2070]), .A2(n6582), .B1(n11399), .B2(n9008), .ZN(
        n6588) );
  INV_X1 U7099 ( .A(n6589), .ZN(n11390) );
  AOI22_X1 U7100 ( .A1(ram[2071]), .A2(n6582), .B1(n11399), .B2(n9032), .ZN(
        n6589) );
  INV_X1 U7101 ( .A(n6590), .ZN(n11391) );
  AOI22_X1 U7102 ( .A1(ram[2072]), .A2(n6582), .B1(n11399), .B2(n9056), .ZN(
        n6590) );
  INV_X1 U7103 ( .A(n6591), .ZN(n11392) );
  AOI22_X1 U7104 ( .A1(ram[2073]), .A2(n6582), .B1(n11399), .B2(n9080), .ZN(
        n6591) );
  INV_X1 U7105 ( .A(n6592), .ZN(n11393) );
  AOI22_X1 U7106 ( .A1(ram[2074]), .A2(n6582), .B1(n11399), .B2(n9104), .ZN(
        n6592) );
  INV_X1 U7107 ( .A(n6593), .ZN(n11394) );
  AOI22_X1 U7108 ( .A1(ram[2075]), .A2(n6582), .B1(n11399), .B2(n9128), .ZN(
        n6593) );
  INV_X1 U7109 ( .A(n6594), .ZN(n11395) );
  AOI22_X1 U7110 ( .A1(ram[2076]), .A2(n6582), .B1(n11399), .B2(n9152), .ZN(
        n6594) );
  INV_X1 U7111 ( .A(n6595), .ZN(n11396) );
  AOI22_X1 U7112 ( .A1(ram[2077]), .A2(n6582), .B1(n11399), .B2(n9176), .ZN(
        n6595) );
  INV_X1 U7113 ( .A(n6596), .ZN(n11397) );
  AOI22_X1 U7114 ( .A1(ram[2078]), .A2(n6582), .B1(n11399), .B2(n9200), .ZN(
        n6596) );
  INV_X1 U7115 ( .A(n6597), .ZN(n11398) );
  AOI22_X1 U7116 ( .A1(ram[2079]), .A2(n6582), .B1(n11399), .B2(n9224), .ZN(
        n6597) );
  INV_X1 U7117 ( .A(n6615), .ZN(n11349) );
  AOI22_X1 U7118 ( .A1(ram[2096]), .A2(n6616), .B1(n11365), .B2(n8864), .ZN(
        n6615) );
  INV_X1 U7119 ( .A(n6617), .ZN(n11350) );
  AOI22_X1 U7120 ( .A1(ram[2097]), .A2(n6616), .B1(n11365), .B2(n8888), .ZN(
        n6617) );
  INV_X1 U7121 ( .A(n6618), .ZN(n11351) );
  AOI22_X1 U7122 ( .A1(ram[2098]), .A2(n6616), .B1(n11365), .B2(n8912), .ZN(
        n6618) );
  INV_X1 U7123 ( .A(n6619), .ZN(n11352) );
  AOI22_X1 U7124 ( .A1(ram[2099]), .A2(n6616), .B1(n11365), .B2(n8936), .ZN(
        n6619) );
  INV_X1 U7125 ( .A(n6620), .ZN(n11353) );
  AOI22_X1 U7126 ( .A1(ram[2100]), .A2(n6616), .B1(n11365), .B2(n8960), .ZN(
        n6620) );
  INV_X1 U7127 ( .A(n6621), .ZN(n11354) );
  AOI22_X1 U7128 ( .A1(ram[2101]), .A2(n6616), .B1(n11365), .B2(n8984), .ZN(
        n6621) );
  INV_X1 U7129 ( .A(n6622), .ZN(n11355) );
  AOI22_X1 U7130 ( .A1(ram[2102]), .A2(n6616), .B1(n11365), .B2(n9008), .ZN(
        n6622) );
  INV_X1 U7131 ( .A(n6623), .ZN(n11356) );
  AOI22_X1 U7132 ( .A1(ram[2103]), .A2(n6616), .B1(n11365), .B2(n9032), .ZN(
        n6623) );
  INV_X1 U7133 ( .A(n6624), .ZN(n11357) );
  AOI22_X1 U7134 ( .A1(ram[2104]), .A2(n6616), .B1(n11365), .B2(n9056), .ZN(
        n6624) );
  INV_X1 U7135 ( .A(n6625), .ZN(n11358) );
  AOI22_X1 U7136 ( .A1(ram[2105]), .A2(n6616), .B1(n11365), .B2(n9080), .ZN(
        n6625) );
  INV_X1 U7137 ( .A(n6626), .ZN(n11359) );
  AOI22_X1 U7138 ( .A1(ram[2106]), .A2(n6616), .B1(n11365), .B2(n9104), .ZN(
        n6626) );
  INV_X1 U7139 ( .A(n6627), .ZN(n11360) );
  AOI22_X1 U7140 ( .A1(ram[2107]), .A2(n6616), .B1(n11365), .B2(n9128), .ZN(
        n6627) );
  INV_X1 U7141 ( .A(n6628), .ZN(n11361) );
  AOI22_X1 U7142 ( .A1(ram[2108]), .A2(n6616), .B1(n11365), .B2(n9152), .ZN(
        n6628) );
  INV_X1 U7143 ( .A(n6629), .ZN(n11362) );
  AOI22_X1 U7144 ( .A1(ram[2109]), .A2(n6616), .B1(n11365), .B2(n9176), .ZN(
        n6629) );
  INV_X1 U7145 ( .A(n6630), .ZN(n11363) );
  AOI22_X1 U7146 ( .A1(ram[2110]), .A2(n6616), .B1(n11365), .B2(n9200), .ZN(
        n6630) );
  INV_X1 U7147 ( .A(n6631), .ZN(n11364) );
  AOI22_X1 U7148 ( .A1(ram[2111]), .A2(n6616), .B1(n11365), .B2(n9224), .ZN(
        n6631) );
  INV_X1 U7149 ( .A(n6649), .ZN(n11315) );
  AOI22_X1 U7150 ( .A1(ram[2128]), .A2(n6650), .B1(n11331), .B2(n8864), .ZN(
        n6649) );
  INV_X1 U7151 ( .A(n6651), .ZN(n11316) );
  AOI22_X1 U7152 ( .A1(ram[2129]), .A2(n6650), .B1(n11331), .B2(n8888), .ZN(
        n6651) );
  INV_X1 U7153 ( .A(n6652), .ZN(n11317) );
  AOI22_X1 U7154 ( .A1(ram[2130]), .A2(n6650), .B1(n11331), .B2(n8912), .ZN(
        n6652) );
  INV_X1 U7155 ( .A(n6653), .ZN(n11318) );
  AOI22_X1 U7156 ( .A1(ram[2131]), .A2(n6650), .B1(n11331), .B2(n8936), .ZN(
        n6653) );
  INV_X1 U7157 ( .A(n6654), .ZN(n11319) );
  AOI22_X1 U7158 ( .A1(ram[2132]), .A2(n6650), .B1(n11331), .B2(n8960), .ZN(
        n6654) );
  INV_X1 U7159 ( .A(n6655), .ZN(n11320) );
  AOI22_X1 U7160 ( .A1(ram[2133]), .A2(n6650), .B1(n11331), .B2(n8984), .ZN(
        n6655) );
  INV_X1 U7161 ( .A(n6656), .ZN(n11321) );
  AOI22_X1 U7162 ( .A1(ram[2134]), .A2(n6650), .B1(n11331), .B2(n9008), .ZN(
        n6656) );
  INV_X1 U7163 ( .A(n6657), .ZN(n11322) );
  AOI22_X1 U7164 ( .A1(ram[2135]), .A2(n6650), .B1(n11331), .B2(n9032), .ZN(
        n6657) );
  INV_X1 U7165 ( .A(n6658), .ZN(n11323) );
  AOI22_X1 U7166 ( .A1(ram[2136]), .A2(n6650), .B1(n11331), .B2(n9056), .ZN(
        n6658) );
  INV_X1 U7167 ( .A(n6659), .ZN(n11324) );
  AOI22_X1 U7168 ( .A1(ram[2137]), .A2(n6650), .B1(n11331), .B2(n9080), .ZN(
        n6659) );
  INV_X1 U7169 ( .A(n6660), .ZN(n11325) );
  AOI22_X1 U7170 ( .A1(ram[2138]), .A2(n6650), .B1(n11331), .B2(n9104), .ZN(
        n6660) );
  INV_X1 U7171 ( .A(n6661), .ZN(n11326) );
  AOI22_X1 U7172 ( .A1(ram[2139]), .A2(n6650), .B1(n11331), .B2(n9128), .ZN(
        n6661) );
  INV_X1 U7173 ( .A(n6662), .ZN(n11327) );
  AOI22_X1 U7174 ( .A1(ram[2140]), .A2(n6650), .B1(n11331), .B2(n9152), .ZN(
        n6662) );
  INV_X1 U7175 ( .A(n6663), .ZN(n11328) );
  AOI22_X1 U7176 ( .A1(ram[2141]), .A2(n6650), .B1(n11331), .B2(n9176), .ZN(
        n6663) );
  INV_X1 U7177 ( .A(n6664), .ZN(n11329) );
  AOI22_X1 U7178 ( .A1(ram[2142]), .A2(n6650), .B1(n11331), .B2(n9200), .ZN(
        n6664) );
  INV_X1 U7179 ( .A(n6665), .ZN(n11330) );
  AOI22_X1 U7180 ( .A1(ram[2143]), .A2(n6650), .B1(n11331), .B2(n9224), .ZN(
        n6665) );
  INV_X1 U7181 ( .A(n6683), .ZN(n11281) );
  AOI22_X1 U7182 ( .A1(ram[2160]), .A2(n6684), .B1(n11297), .B2(n8864), .ZN(
        n6683) );
  INV_X1 U7183 ( .A(n6685), .ZN(n11282) );
  AOI22_X1 U7184 ( .A1(ram[2161]), .A2(n6684), .B1(n11297), .B2(n8888), .ZN(
        n6685) );
  INV_X1 U7185 ( .A(n6686), .ZN(n11283) );
  AOI22_X1 U7186 ( .A1(ram[2162]), .A2(n6684), .B1(n11297), .B2(n8912), .ZN(
        n6686) );
  INV_X1 U7187 ( .A(n6687), .ZN(n11284) );
  AOI22_X1 U7188 ( .A1(ram[2163]), .A2(n6684), .B1(n11297), .B2(n8936), .ZN(
        n6687) );
  INV_X1 U7189 ( .A(n6688), .ZN(n11285) );
  AOI22_X1 U7190 ( .A1(ram[2164]), .A2(n6684), .B1(n11297), .B2(n8960), .ZN(
        n6688) );
  INV_X1 U7191 ( .A(n6689), .ZN(n11286) );
  AOI22_X1 U7192 ( .A1(ram[2165]), .A2(n6684), .B1(n11297), .B2(n8984), .ZN(
        n6689) );
  INV_X1 U7193 ( .A(n6690), .ZN(n11287) );
  AOI22_X1 U7194 ( .A1(ram[2166]), .A2(n6684), .B1(n11297), .B2(n9008), .ZN(
        n6690) );
  INV_X1 U7195 ( .A(n6691), .ZN(n11288) );
  AOI22_X1 U7196 ( .A1(ram[2167]), .A2(n6684), .B1(n11297), .B2(n9032), .ZN(
        n6691) );
  INV_X1 U7197 ( .A(n6692), .ZN(n11289) );
  AOI22_X1 U7198 ( .A1(ram[2168]), .A2(n6684), .B1(n11297), .B2(n9056), .ZN(
        n6692) );
  INV_X1 U7199 ( .A(n6693), .ZN(n11290) );
  AOI22_X1 U7200 ( .A1(ram[2169]), .A2(n6684), .B1(n11297), .B2(n9080), .ZN(
        n6693) );
  INV_X1 U7201 ( .A(n6694), .ZN(n11291) );
  AOI22_X1 U7202 ( .A1(ram[2170]), .A2(n6684), .B1(n11297), .B2(n9104), .ZN(
        n6694) );
  INV_X1 U7203 ( .A(n6695), .ZN(n11292) );
  AOI22_X1 U7204 ( .A1(ram[2171]), .A2(n6684), .B1(n11297), .B2(n9128), .ZN(
        n6695) );
  INV_X1 U7205 ( .A(n6696), .ZN(n11293) );
  AOI22_X1 U7206 ( .A1(ram[2172]), .A2(n6684), .B1(n11297), .B2(n9152), .ZN(
        n6696) );
  INV_X1 U7207 ( .A(n6697), .ZN(n11294) );
  AOI22_X1 U7208 ( .A1(ram[2173]), .A2(n6684), .B1(n11297), .B2(n9176), .ZN(
        n6697) );
  INV_X1 U7209 ( .A(n6698), .ZN(n11295) );
  AOI22_X1 U7210 ( .A1(ram[2174]), .A2(n6684), .B1(n11297), .B2(n9200), .ZN(
        n6698) );
  INV_X1 U7211 ( .A(n6699), .ZN(n11296) );
  AOI22_X1 U7212 ( .A1(ram[2175]), .A2(n6684), .B1(n11297), .B2(n9224), .ZN(
        n6699) );
  INV_X1 U7213 ( .A(n6717), .ZN(n11247) );
  AOI22_X1 U7214 ( .A1(ram[2192]), .A2(n6718), .B1(n11263), .B2(n8863), .ZN(
        n6717) );
  INV_X1 U7215 ( .A(n6719), .ZN(n11248) );
  AOI22_X1 U7216 ( .A1(ram[2193]), .A2(n6718), .B1(n11263), .B2(n8887), .ZN(
        n6719) );
  INV_X1 U7217 ( .A(n6720), .ZN(n11249) );
  AOI22_X1 U7218 ( .A1(ram[2194]), .A2(n6718), .B1(n11263), .B2(n8911), .ZN(
        n6720) );
  INV_X1 U7219 ( .A(n6721), .ZN(n11250) );
  AOI22_X1 U7220 ( .A1(ram[2195]), .A2(n6718), .B1(n11263), .B2(n8935), .ZN(
        n6721) );
  INV_X1 U7221 ( .A(n6722), .ZN(n11251) );
  AOI22_X1 U7222 ( .A1(ram[2196]), .A2(n6718), .B1(n11263), .B2(n8959), .ZN(
        n6722) );
  INV_X1 U7223 ( .A(n6723), .ZN(n11252) );
  AOI22_X1 U7224 ( .A1(ram[2197]), .A2(n6718), .B1(n11263), .B2(n8983), .ZN(
        n6723) );
  INV_X1 U7225 ( .A(n6724), .ZN(n11253) );
  AOI22_X1 U7226 ( .A1(ram[2198]), .A2(n6718), .B1(n11263), .B2(n9007), .ZN(
        n6724) );
  INV_X1 U7227 ( .A(n6725), .ZN(n11254) );
  AOI22_X1 U7228 ( .A1(ram[2199]), .A2(n6718), .B1(n11263), .B2(n9031), .ZN(
        n6725) );
  INV_X1 U7229 ( .A(n6726), .ZN(n11255) );
  AOI22_X1 U7230 ( .A1(ram[2200]), .A2(n6718), .B1(n11263), .B2(n9055), .ZN(
        n6726) );
  INV_X1 U7231 ( .A(n6727), .ZN(n11256) );
  AOI22_X1 U7232 ( .A1(ram[2201]), .A2(n6718), .B1(n11263), .B2(n9079), .ZN(
        n6727) );
  INV_X1 U7233 ( .A(n6728), .ZN(n11257) );
  AOI22_X1 U7234 ( .A1(ram[2202]), .A2(n6718), .B1(n11263), .B2(n9103), .ZN(
        n6728) );
  INV_X1 U7235 ( .A(n6729), .ZN(n11258) );
  AOI22_X1 U7236 ( .A1(ram[2203]), .A2(n6718), .B1(n11263), .B2(n9127), .ZN(
        n6729) );
  INV_X1 U7237 ( .A(n6730), .ZN(n11259) );
  AOI22_X1 U7238 ( .A1(ram[2204]), .A2(n6718), .B1(n11263), .B2(n9151), .ZN(
        n6730) );
  INV_X1 U7239 ( .A(n6731), .ZN(n11260) );
  AOI22_X1 U7240 ( .A1(ram[2205]), .A2(n6718), .B1(n11263), .B2(n9175), .ZN(
        n6731) );
  INV_X1 U7241 ( .A(n6732), .ZN(n11261) );
  AOI22_X1 U7242 ( .A1(ram[2206]), .A2(n6718), .B1(n11263), .B2(n9199), .ZN(
        n6732) );
  INV_X1 U7243 ( .A(n6733), .ZN(n11262) );
  AOI22_X1 U7244 ( .A1(ram[2207]), .A2(n6718), .B1(n11263), .B2(n9223), .ZN(
        n6733) );
  INV_X1 U7245 ( .A(n6751), .ZN(n11213) );
  AOI22_X1 U7246 ( .A1(ram[2224]), .A2(n6752), .B1(n11229), .B2(n8863), .ZN(
        n6751) );
  INV_X1 U7247 ( .A(n6753), .ZN(n11214) );
  AOI22_X1 U7248 ( .A1(ram[2225]), .A2(n6752), .B1(n11229), .B2(n8887), .ZN(
        n6753) );
  INV_X1 U7249 ( .A(n6754), .ZN(n11215) );
  AOI22_X1 U7250 ( .A1(ram[2226]), .A2(n6752), .B1(n11229), .B2(n8911), .ZN(
        n6754) );
  INV_X1 U7251 ( .A(n6755), .ZN(n11216) );
  AOI22_X1 U7252 ( .A1(ram[2227]), .A2(n6752), .B1(n11229), .B2(n8935), .ZN(
        n6755) );
  INV_X1 U7253 ( .A(n6756), .ZN(n11217) );
  AOI22_X1 U7254 ( .A1(ram[2228]), .A2(n6752), .B1(n11229), .B2(n8959), .ZN(
        n6756) );
  INV_X1 U7255 ( .A(n6757), .ZN(n11218) );
  AOI22_X1 U7256 ( .A1(ram[2229]), .A2(n6752), .B1(n11229), .B2(n8983), .ZN(
        n6757) );
  INV_X1 U7257 ( .A(n6758), .ZN(n11219) );
  AOI22_X1 U7258 ( .A1(ram[2230]), .A2(n6752), .B1(n11229), .B2(n9007), .ZN(
        n6758) );
  INV_X1 U7259 ( .A(n6759), .ZN(n11220) );
  AOI22_X1 U7260 ( .A1(ram[2231]), .A2(n6752), .B1(n11229), .B2(n9031), .ZN(
        n6759) );
  INV_X1 U7261 ( .A(n6760), .ZN(n11221) );
  AOI22_X1 U7262 ( .A1(ram[2232]), .A2(n6752), .B1(n11229), .B2(n9055), .ZN(
        n6760) );
  INV_X1 U7263 ( .A(n6761), .ZN(n11222) );
  AOI22_X1 U7264 ( .A1(ram[2233]), .A2(n6752), .B1(n11229), .B2(n9079), .ZN(
        n6761) );
  INV_X1 U7265 ( .A(n6762), .ZN(n11223) );
  AOI22_X1 U7266 ( .A1(ram[2234]), .A2(n6752), .B1(n11229), .B2(n9103), .ZN(
        n6762) );
  INV_X1 U7267 ( .A(n6763), .ZN(n11224) );
  AOI22_X1 U7268 ( .A1(ram[2235]), .A2(n6752), .B1(n11229), .B2(n9127), .ZN(
        n6763) );
  INV_X1 U7269 ( .A(n6764), .ZN(n11225) );
  AOI22_X1 U7270 ( .A1(ram[2236]), .A2(n6752), .B1(n11229), .B2(n9151), .ZN(
        n6764) );
  INV_X1 U7271 ( .A(n6765), .ZN(n11226) );
  AOI22_X1 U7272 ( .A1(ram[2237]), .A2(n6752), .B1(n11229), .B2(n9175), .ZN(
        n6765) );
  INV_X1 U7273 ( .A(n6766), .ZN(n11227) );
  AOI22_X1 U7274 ( .A1(ram[2238]), .A2(n6752), .B1(n11229), .B2(n9199), .ZN(
        n6766) );
  INV_X1 U7275 ( .A(n6767), .ZN(n11228) );
  AOI22_X1 U7276 ( .A1(ram[2239]), .A2(n6752), .B1(n11229), .B2(n9223), .ZN(
        n6767) );
  INV_X1 U7277 ( .A(n6785), .ZN(n11179) );
  AOI22_X1 U7278 ( .A1(ram[2256]), .A2(n6786), .B1(n11195), .B2(n8863), .ZN(
        n6785) );
  INV_X1 U7279 ( .A(n6787), .ZN(n11180) );
  AOI22_X1 U7280 ( .A1(ram[2257]), .A2(n6786), .B1(n11195), .B2(n8887), .ZN(
        n6787) );
  INV_X1 U7281 ( .A(n6788), .ZN(n11181) );
  AOI22_X1 U7282 ( .A1(ram[2258]), .A2(n6786), .B1(n11195), .B2(n8911), .ZN(
        n6788) );
  INV_X1 U7283 ( .A(n6789), .ZN(n11182) );
  AOI22_X1 U7284 ( .A1(ram[2259]), .A2(n6786), .B1(n11195), .B2(n8935), .ZN(
        n6789) );
  INV_X1 U7285 ( .A(n6790), .ZN(n11183) );
  AOI22_X1 U7286 ( .A1(ram[2260]), .A2(n6786), .B1(n11195), .B2(n8959), .ZN(
        n6790) );
  INV_X1 U7287 ( .A(n6791), .ZN(n11184) );
  AOI22_X1 U7288 ( .A1(ram[2261]), .A2(n6786), .B1(n11195), .B2(n8983), .ZN(
        n6791) );
  INV_X1 U7289 ( .A(n6792), .ZN(n11185) );
  AOI22_X1 U7290 ( .A1(ram[2262]), .A2(n6786), .B1(n11195), .B2(n9007), .ZN(
        n6792) );
  INV_X1 U7291 ( .A(n6793), .ZN(n11186) );
  AOI22_X1 U7292 ( .A1(ram[2263]), .A2(n6786), .B1(n11195), .B2(n9031), .ZN(
        n6793) );
  INV_X1 U7293 ( .A(n6794), .ZN(n11187) );
  AOI22_X1 U7294 ( .A1(ram[2264]), .A2(n6786), .B1(n11195), .B2(n9055), .ZN(
        n6794) );
  INV_X1 U7295 ( .A(n6795), .ZN(n11188) );
  AOI22_X1 U7296 ( .A1(ram[2265]), .A2(n6786), .B1(n11195), .B2(n9079), .ZN(
        n6795) );
  INV_X1 U7297 ( .A(n6796), .ZN(n11189) );
  AOI22_X1 U7298 ( .A1(ram[2266]), .A2(n6786), .B1(n11195), .B2(n9103), .ZN(
        n6796) );
  INV_X1 U7299 ( .A(n6797), .ZN(n11190) );
  AOI22_X1 U7300 ( .A1(ram[2267]), .A2(n6786), .B1(n11195), .B2(n9127), .ZN(
        n6797) );
  INV_X1 U7301 ( .A(n6798), .ZN(n11191) );
  AOI22_X1 U7302 ( .A1(ram[2268]), .A2(n6786), .B1(n11195), .B2(n9151), .ZN(
        n6798) );
  INV_X1 U7303 ( .A(n6799), .ZN(n11192) );
  AOI22_X1 U7304 ( .A1(ram[2269]), .A2(n6786), .B1(n11195), .B2(n9175), .ZN(
        n6799) );
  INV_X1 U7305 ( .A(n6800), .ZN(n11193) );
  AOI22_X1 U7306 ( .A1(ram[2270]), .A2(n6786), .B1(n11195), .B2(n9199), .ZN(
        n6800) );
  INV_X1 U7307 ( .A(n6801), .ZN(n11194) );
  AOI22_X1 U7308 ( .A1(ram[2271]), .A2(n6786), .B1(n11195), .B2(n9223), .ZN(
        n6801) );
  INV_X1 U7309 ( .A(n6819), .ZN(n11145) );
  AOI22_X1 U7310 ( .A1(ram[2288]), .A2(n6820), .B1(n11161), .B2(n8863), .ZN(
        n6819) );
  INV_X1 U7311 ( .A(n6821), .ZN(n11146) );
  AOI22_X1 U7312 ( .A1(ram[2289]), .A2(n6820), .B1(n11161), .B2(n8887), .ZN(
        n6821) );
  INV_X1 U7313 ( .A(n6822), .ZN(n11147) );
  AOI22_X1 U7314 ( .A1(ram[2290]), .A2(n6820), .B1(n11161), .B2(n8911), .ZN(
        n6822) );
  INV_X1 U7315 ( .A(n6823), .ZN(n11148) );
  AOI22_X1 U7316 ( .A1(ram[2291]), .A2(n6820), .B1(n11161), .B2(n8935), .ZN(
        n6823) );
  INV_X1 U7317 ( .A(n6824), .ZN(n11149) );
  AOI22_X1 U7318 ( .A1(ram[2292]), .A2(n6820), .B1(n11161), .B2(n8959), .ZN(
        n6824) );
  INV_X1 U7319 ( .A(n6825), .ZN(n11150) );
  AOI22_X1 U7320 ( .A1(ram[2293]), .A2(n6820), .B1(n11161), .B2(n8983), .ZN(
        n6825) );
  INV_X1 U7321 ( .A(n6826), .ZN(n11151) );
  AOI22_X1 U7322 ( .A1(ram[2294]), .A2(n6820), .B1(n11161), .B2(n9007), .ZN(
        n6826) );
  INV_X1 U7323 ( .A(n6827), .ZN(n11152) );
  AOI22_X1 U7324 ( .A1(ram[2295]), .A2(n6820), .B1(n11161), .B2(n9031), .ZN(
        n6827) );
  INV_X1 U7325 ( .A(n6828), .ZN(n11153) );
  AOI22_X1 U7326 ( .A1(ram[2296]), .A2(n6820), .B1(n11161), .B2(n9055), .ZN(
        n6828) );
  INV_X1 U7327 ( .A(n6829), .ZN(n11154) );
  AOI22_X1 U7328 ( .A1(ram[2297]), .A2(n6820), .B1(n11161), .B2(n9079), .ZN(
        n6829) );
  INV_X1 U7329 ( .A(n6830), .ZN(n11155) );
  AOI22_X1 U7330 ( .A1(ram[2298]), .A2(n6820), .B1(n11161), .B2(n9103), .ZN(
        n6830) );
  INV_X1 U7331 ( .A(n6831), .ZN(n11156) );
  AOI22_X1 U7332 ( .A1(ram[2299]), .A2(n6820), .B1(n11161), .B2(n9127), .ZN(
        n6831) );
  INV_X1 U7333 ( .A(n6832), .ZN(n11157) );
  AOI22_X1 U7334 ( .A1(ram[2300]), .A2(n6820), .B1(n11161), .B2(n9151), .ZN(
        n6832) );
  INV_X1 U7335 ( .A(n6833), .ZN(n11158) );
  AOI22_X1 U7336 ( .A1(ram[2301]), .A2(n6820), .B1(n11161), .B2(n9175), .ZN(
        n6833) );
  INV_X1 U7337 ( .A(n6834), .ZN(n11159) );
  AOI22_X1 U7338 ( .A1(ram[2302]), .A2(n6820), .B1(n11161), .B2(n9199), .ZN(
        n6834) );
  INV_X1 U7339 ( .A(n6835), .ZN(n11160) );
  AOI22_X1 U7340 ( .A1(ram[2303]), .A2(n6820), .B1(n11161), .B2(n9223), .ZN(
        n6835) );
  INV_X1 U7341 ( .A(n6855), .ZN(n11111) );
  AOI22_X1 U7342 ( .A1(ram[2320]), .A2(n6856), .B1(n11127), .B2(n8863), .ZN(
        n6855) );
  INV_X1 U7343 ( .A(n6857), .ZN(n11112) );
  AOI22_X1 U7344 ( .A1(ram[2321]), .A2(n6856), .B1(n11127), .B2(n8887), .ZN(
        n6857) );
  INV_X1 U7345 ( .A(n6858), .ZN(n11113) );
  AOI22_X1 U7346 ( .A1(ram[2322]), .A2(n6856), .B1(n11127), .B2(n8911), .ZN(
        n6858) );
  INV_X1 U7347 ( .A(n6859), .ZN(n11114) );
  AOI22_X1 U7348 ( .A1(ram[2323]), .A2(n6856), .B1(n11127), .B2(n8935), .ZN(
        n6859) );
  INV_X1 U7349 ( .A(n6860), .ZN(n11115) );
  AOI22_X1 U7350 ( .A1(ram[2324]), .A2(n6856), .B1(n11127), .B2(n8959), .ZN(
        n6860) );
  INV_X1 U7351 ( .A(n6861), .ZN(n11116) );
  AOI22_X1 U7352 ( .A1(ram[2325]), .A2(n6856), .B1(n11127), .B2(n8983), .ZN(
        n6861) );
  INV_X1 U7353 ( .A(n6862), .ZN(n11117) );
  AOI22_X1 U7354 ( .A1(ram[2326]), .A2(n6856), .B1(n11127), .B2(n9007), .ZN(
        n6862) );
  INV_X1 U7355 ( .A(n6863), .ZN(n11118) );
  AOI22_X1 U7356 ( .A1(ram[2327]), .A2(n6856), .B1(n11127), .B2(n9031), .ZN(
        n6863) );
  INV_X1 U7357 ( .A(n6864), .ZN(n11119) );
  AOI22_X1 U7358 ( .A1(ram[2328]), .A2(n6856), .B1(n11127), .B2(n9055), .ZN(
        n6864) );
  INV_X1 U7359 ( .A(n6865), .ZN(n11120) );
  AOI22_X1 U7360 ( .A1(ram[2329]), .A2(n6856), .B1(n11127), .B2(n9079), .ZN(
        n6865) );
  INV_X1 U7361 ( .A(n6866), .ZN(n11121) );
  AOI22_X1 U7362 ( .A1(ram[2330]), .A2(n6856), .B1(n11127), .B2(n9103), .ZN(
        n6866) );
  INV_X1 U7363 ( .A(n6867), .ZN(n11122) );
  AOI22_X1 U7364 ( .A1(ram[2331]), .A2(n6856), .B1(n11127), .B2(n9127), .ZN(
        n6867) );
  INV_X1 U7365 ( .A(n6868), .ZN(n11123) );
  AOI22_X1 U7366 ( .A1(ram[2332]), .A2(n6856), .B1(n11127), .B2(n9151), .ZN(
        n6868) );
  INV_X1 U7367 ( .A(n6869), .ZN(n11124) );
  AOI22_X1 U7368 ( .A1(ram[2333]), .A2(n6856), .B1(n11127), .B2(n9175), .ZN(
        n6869) );
  INV_X1 U7369 ( .A(n6870), .ZN(n11125) );
  AOI22_X1 U7370 ( .A1(ram[2334]), .A2(n6856), .B1(n11127), .B2(n9199), .ZN(
        n6870) );
  INV_X1 U7371 ( .A(n6871), .ZN(n11126) );
  AOI22_X1 U7372 ( .A1(ram[2335]), .A2(n6856), .B1(n11127), .B2(n9223), .ZN(
        n6871) );
  INV_X1 U7373 ( .A(n6889), .ZN(n11077) );
  AOI22_X1 U7374 ( .A1(ram[2352]), .A2(n6890), .B1(n11093), .B2(n8863), .ZN(
        n6889) );
  INV_X1 U7375 ( .A(n6891), .ZN(n11078) );
  AOI22_X1 U7376 ( .A1(ram[2353]), .A2(n6890), .B1(n11093), .B2(n8887), .ZN(
        n6891) );
  INV_X1 U7377 ( .A(n6892), .ZN(n11079) );
  AOI22_X1 U7378 ( .A1(ram[2354]), .A2(n6890), .B1(n11093), .B2(n8911), .ZN(
        n6892) );
  INV_X1 U7379 ( .A(n6893), .ZN(n11080) );
  AOI22_X1 U7380 ( .A1(ram[2355]), .A2(n6890), .B1(n11093), .B2(n8935), .ZN(
        n6893) );
  INV_X1 U7381 ( .A(n6894), .ZN(n11081) );
  AOI22_X1 U7382 ( .A1(ram[2356]), .A2(n6890), .B1(n11093), .B2(n8959), .ZN(
        n6894) );
  INV_X1 U7383 ( .A(n6895), .ZN(n11082) );
  AOI22_X1 U7384 ( .A1(ram[2357]), .A2(n6890), .B1(n11093), .B2(n8983), .ZN(
        n6895) );
  INV_X1 U7385 ( .A(n6896), .ZN(n11083) );
  AOI22_X1 U7386 ( .A1(ram[2358]), .A2(n6890), .B1(n11093), .B2(n9007), .ZN(
        n6896) );
  INV_X1 U7387 ( .A(n6897), .ZN(n11084) );
  AOI22_X1 U7388 ( .A1(ram[2359]), .A2(n6890), .B1(n11093), .B2(n9031), .ZN(
        n6897) );
  INV_X1 U7389 ( .A(n6898), .ZN(n11085) );
  AOI22_X1 U7390 ( .A1(ram[2360]), .A2(n6890), .B1(n11093), .B2(n9055), .ZN(
        n6898) );
  INV_X1 U7391 ( .A(n6899), .ZN(n11086) );
  AOI22_X1 U7392 ( .A1(ram[2361]), .A2(n6890), .B1(n11093), .B2(n9079), .ZN(
        n6899) );
  INV_X1 U7393 ( .A(n6900), .ZN(n11087) );
  AOI22_X1 U7394 ( .A1(ram[2362]), .A2(n6890), .B1(n11093), .B2(n9103), .ZN(
        n6900) );
  INV_X1 U7395 ( .A(n6901), .ZN(n11088) );
  AOI22_X1 U7396 ( .A1(ram[2363]), .A2(n6890), .B1(n11093), .B2(n9127), .ZN(
        n6901) );
  INV_X1 U7397 ( .A(n6902), .ZN(n11089) );
  AOI22_X1 U7398 ( .A1(ram[2364]), .A2(n6890), .B1(n11093), .B2(n9151), .ZN(
        n6902) );
  INV_X1 U7399 ( .A(n6903), .ZN(n11090) );
  AOI22_X1 U7400 ( .A1(ram[2365]), .A2(n6890), .B1(n11093), .B2(n9175), .ZN(
        n6903) );
  INV_X1 U7401 ( .A(n6904), .ZN(n11091) );
  AOI22_X1 U7402 ( .A1(ram[2366]), .A2(n6890), .B1(n11093), .B2(n9199), .ZN(
        n6904) );
  INV_X1 U7403 ( .A(n6905), .ZN(n11092) );
  AOI22_X1 U7404 ( .A1(ram[2367]), .A2(n6890), .B1(n11093), .B2(n9223), .ZN(
        n6905) );
  INV_X1 U7405 ( .A(n6923), .ZN(n11043) );
  AOI22_X1 U7406 ( .A1(ram[2384]), .A2(n6924), .B1(n11059), .B2(n8862), .ZN(
        n6923) );
  INV_X1 U7407 ( .A(n6925), .ZN(n11044) );
  AOI22_X1 U7408 ( .A1(ram[2385]), .A2(n6924), .B1(n11059), .B2(n8886), .ZN(
        n6925) );
  INV_X1 U7409 ( .A(n6926), .ZN(n11045) );
  AOI22_X1 U7410 ( .A1(ram[2386]), .A2(n6924), .B1(n11059), .B2(n8910), .ZN(
        n6926) );
  INV_X1 U7411 ( .A(n6927), .ZN(n11046) );
  AOI22_X1 U7412 ( .A1(ram[2387]), .A2(n6924), .B1(n11059), .B2(n8934), .ZN(
        n6927) );
  INV_X1 U7413 ( .A(n6928), .ZN(n11047) );
  AOI22_X1 U7414 ( .A1(ram[2388]), .A2(n6924), .B1(n11059), .B2(n8958), .ZN(
        n6928) );
  INV_X1 U7415 ( .A(n6929), .ZN(n11048) );
  AOI22_X1 U7416 ( .A1(ram[2389]), .A2(n6924), .B1(n11059), .B2(n8982), .ZN(
        n6929) );
  INV_X1 U7417 ( .A(n6930), .ZN(n11049) );
  AOI22_X1 U7418 ( .A1(ram[2390]), .A2(n6924), .B1(n11059), .B2(n9006), .ZN(
        n6930) );
  INV_X1 U7419 ( .A(n6931), .ZN(n11050) );
  AOI22_X1 U7420 ( .A1(ram[2391]), .A2(n6924), .B1(n11059), .B2(n9030), .ZN(
        n6931) );
  INV_X1 U7421 ( .A(n6932), .ZN(n11051) );
  AOI22_X1 U7422 ( .A1(ram[2392]), .A2(n6924), .B1(n11059), .B2(n9054), .ZN(
        n6932) );
  INV_X1 U7423 ( .A(n6933), .ZN(n11052) );
  AOI22_X1 U7424 ( .A1(ram[2393]), .A2(n6924), .B1(n11059), .B2(n9078), .ZN(
        n6933) );
  INV_X1 U7425 ( .A(n6934), .ZN(n11053) );
  AOI22_X1 U7426 ( .A1(ram[2394]), .A2(n6924), .B1(n11059), .B2(n9102), .ZN(
        n6934) );
  INV_X1 U7427 ( .A(n6935), .ZN(n11054) );
  AOI22_X1 U7428 ( .A1(ram[2395]), .A2(n6924), .B1(n11059), .B2(n9126), .ZN(
        n6935) );
  INV_X1 U7429 ( .A(n6936), .ZN(n11055) );
  AOI22_X1 U7430 ( .A1(ram[2396]), .A2(n6924), .B1(n11059), .B2(n9150), .ZN(
        n6936) );
  INV_X1 U7431 ( .A(n6937), .ZN(n11056) );
  AOI22_X1 U7432 ( .A1(ram[2397]), .A2(n6924), .B1(n11059), .B2(n9174), .ZN(
        n6937) );
  INV_X1 U7433 ( .A(n6938), .ZN(n11057) );
  AOI22_X1 U7434 ( .A1(ram[2398]), .A2(n6924), .B1(n11059), .B2(n9198), .ZN(
        n6938) );
  INV_X1 U7435 ( .A(n6939), .ZN(n11058) );
  AOI22_X1 U7436 ( .A1(ram[2399]), .A2(n6924), .B1(n11059), .B2(n9222), .ZN(
        n6939) );
  INV_X1 U7437 ( .A(n6957), .ZN(n11009) );
  AOI22_X1 U7438 ( .A1(ram[2416]), .A2(n6958), .B1(n11025), .B2(n8862), .ZN(
        n6957) );
  INV_X1 U7439 ( .A(n6959), .ZN(n11010) );
  AOI22_X1 U7440 ( .A1(ram[2417]), .A2(n6958), .B1(n11025), .B2(n8886), .ZN(
        n6959) );
  INV_X1 U7441 ( .A(n6960), .ZN(n11011) );
  AOI22_X1 U7442 ( .A1(ram[2418]), .A2(n6958), .B1(n11025), .B2(n8910), .ZN(
        n6960) );
  INV_X1 U7443 ( .A(n6961), .ZN(n11012) );
  AOI22_X1 U7444 ( .A1(ram[2419]), .A2(n6958), .B1(n11025), .B2(n8934), .ZN(
        n6961) );
  INV_X1 U7445 ( .A(n6962), .ZN(n11013) );
  AOI22_X1 U7446 ( .A1(ram[2420]), .A2(n6958), .B1(n11025), .B2(n8958), .ZN(
        n6962) );
  INV_X1 U7447 ( .A(n6963), .ZN(n11014) );
  AOI22_X1 U7448 ( .A1(ram[2421]), .A2(n6958), .B1(n11025), .B2(n8982), .ZN(
        n6963) );
  INV_X1 U7449 ( .A(n6964), .ZN(n11015) );
  AOI22_X1 U7450 ( .A1(ram[2422]), .A2(n6958), .B1(n11025), .B2(n9006), .ZN(
        n6964) );
  INV_X1 U7451 ( .A(n6965), .ZN(n11016) );
  AOI22_X1 U7452 ( .A1(ram[2423]), .A2(n6958), .B1(n11025), .B2(n9030), .ZN(
        n6965) );
  INV_X1 U7453 ( .A(n6966), .ZN(n11017) );
  AOI22_X1 U7454 ( .A1(ram[2424]), .A2(n6958), .B1(n11025), .B2(n9054), .ZN(
        n6966) );
  INV_X1 U7455 ( .A(n6967), .ZN(n11018) );
  AOI22_X1 U7456 ( .A1(ram[2425]), .A2(n6958), .B1(n11025), .B2(n9078), .ZN(
        n6967) );
  INV_X1 U7457 ( .A(n6968), .ZN(n11019) );
  AOI22_X1 U7458 ( .A1(ram[2426]), .A2(n6958), .B1(n11025), .B2(n9102), .ZN(
        n6968) );
  INV_X1 U7459 ( .A(n6969), .ZN(n11020) );
  AOI22_X1 U7460 ( .A1(ram[2427]), .A2(n6958), .B1(n11025), .B2(n9126), .ZN(
        n6969) );
  INV_X1 U7461 ( .A(n6970), .ZN(n11021) );
  AOI22_X1 U7462 ( .A1(ram[2428]), .A2(n6958), .B1(n11025), .B2(n9150), .ZN(
        n6970) );
  INV_X1 U7463 ( .A(n6971), .ZN(n11022) );
  AOI22_X1 U7464 ( .A1(ram[2429]), .A2(n6958), .B1(n11025), .B2(n9174), .ZN(
        n6971) );
  INV_X1 U7465 ( .A(n6972), .ZN(n11023) );
  AOI22_X1 U7466 ( .A1(ram[2430]), .A2(n6958), .B1(n11025), .B2(n9198), .ZN(
        n6972) );
  INV_X1 U7467 ( .A(n6973), .ZN(n11024) );
  AOI22_X1 U7468 ( .A1(ram[2431]), .A2(n6958), .B1(n11025), .B2(n9222), .ZN(
        n6973) );
  INV_X1 U7469 ( .A(n6991), .ZN(n10975) );
  AOI22_X1 U7470 ( .A1(ram[2448]), .A2(n6992), .B1(n10991), .B2(n8862), .ZN(
        n6991) );
  INV_X1 U7471 ( .A(n6993), .ZN(n10976) );
  AOI22_X1 U7472 ( .A1(ram[2449]), .A2(n6992), .B1(n10991), .B2(n8886), .ZN(
        n6993) );
  INV_X1 U7473 ( .A(n6994), .ZN(n10977) );
  AOI22_X1 U7474 ( .A1(ram[2450]), .A2(n6992), .B1(n10991), .B2(n8910), .ZN(
        n6994) );
  INV_X1 U7475 ( .A(n6995), .ZN(n10978) );
  AOI22_X1 U7476 ( .A1(ram[2451]), .A2(n6992), .B1(n10991), .B2(n8934), .ZN(
        n6995) );
  INV_X1 U7477 ( .A(n6996), .ZN(n10979) );
  AOI22_X1 U7478 ( .A1(ram[2452]), .A2(n6992), .B1(n10991), .B2(n8958), .ZN(
        n6996) );
  INV_X1 U7479 ( .A(n6997), .ZN(n10980) );
  AOI22_X1 U7480 ( .A1(ram[2453]), .A2(n6992), .B1(n10991), .B2(n8982), .ZN(
        n6997) );
  INV_X1 U7481 ( .A(n6998), .ZN(n10981) );
  AOI22_X1 U7482 ( .A1(ram[2454]), .A2(n6992), .B1(n10991), .B2(n9006), .ZN(
        n6998) );
  INV_X1 U7483 ( .A(n6999), .ZN(n10982) );
  AOI22_X1 U7484 ( .A1(ram[2455]), .A2(n6992), .B1(n10991), .B2(n9030), .ZN(
        n6999) );
  INV_X1 U7485 ( .A(n7000), .ZN(n10983) );
  AOI22_X1 U7486 ( .A1(ram[2456]), .A2(n6992), .B1(n10991), .B2(n9054), .ZN(
        n7000) );
  INV_X1 U7487 ( .A(n7001), .ZN(n10984) );
  AOI22_X1 U7488 ( .A1(ram[2457]), .A2(n6992), .B1(n10991), .B2(n9078), .ZN(
        n7001) );
  INV_X1 U7489 ( .A(n7002), .ZN(n10985) );
  AOI22_X1 U7490 ( .A1(ram[2458]), .A2(n6992), .B1(n10991), .B2(n9102), .ZN(
        n7002) );
  INV_X1 U7491 ( .A(n7003), .ZN(n10986) );
  AOI22_X1 U7492 ( .A1(ram[2459]), .A2(n6992), .B1(n10991), .B2(n9126), .ZN(
        n7003) );
  INV_X1 U7493 ( .A(n7004), .ZN(n10987) );
  AOI22_X1 U7494 ( .A1(ram[2460]), .A2(n6992), .B1(n10991), .B2(n9150), .ZN(
        n7004) );
  INV_X1 U7495 ( .A(n7005), .ZN(n10988) );
  AOI22_X1 U7496 ( .A1(ram[2461]), .A2(n6992), .B1(n10991), .B2(n9174), .ZN(
        n7005) );
  INV_X1 U7497 ( .A(n7006), .ZN(n10989) );
  AOI22_X1 U7498 ( .A1(ram[2462]), .A2(n6992), .B1(n10991), .B2(n9198), .ZN(
        n7006) );
  INV_X1 U7499 ( .A(n7007), .ZN(n10990) );
  AOI22_X1 U7500 ( .A1(ram[2463]), .A2(n6992), .B1(n10991), .B2(n9222), .ZN(
        n7007) );
  INV_X1 U7501 ( .A(n7025), .ZN(n10941) );
  AOI22_X1 U7502 ( .A1(ram[2480]), .A2(n7026), .B1(n10957), .B2(n8862), .ZN(
        n7025) );
  INV_X1 U7503 ( .A(n7027), .ZN(n10942) );
  AOI22_X1 U7504 ( .A1(ram[2481]), .A2(n7026), .B1(n10957), .B2(n8886), .ZN(
        n7027) );
  INV_X1 U7505 ( .A(n7028), .ZN(n10943) );
  AOI22_X1 U7506 ( .A1(ram[2482]), .A2(n7026), .B1(n10957), .B2(n8910), .ZN(
        n7028) );
  INV_X1 U7507 ( .A(n7029), .ZN(n10944) );
  AOI22_X1 U7508 ( .A1(ram[2483]), .A2(n7026), .B1(n10957), .B2(n8934), .ZN(
        n7029) );
  INV_X1 U7509 ( .A(n7030), .ZN(n10945) );
  AOI22_X1 U7510 ( .A1(ram[2484]), .A2(n7026), .B1(n10957), .B2(n8958), .ZN(
        n7030) );
  INV_X1 U7511 ( .A(n7031), .ZN(n10946) );
  AOI22_X1 U7512 ( .A1(ram[2485]), .A2(n7026), .B1(n10957), .B2(n8982), .ZN(
        n7031) );
  INV_X1 U7513 ( .A(n7032), .ZN(n10947) );
  AOI22_X1 U7514 ( .A1(ram[2486]), .A2(n7026), .B1(n10957), .B2(n9006), .ZN(
        n7032) );
  INV_X1 U7515 ( .A(n7033), .ZN(n10948) );
  AOI22_X1 U7516 ( .A1(ram[2487]), .A2(n7026), .B1(n10957), .B2(n9030), .ZN(
        n7033) );
  INV_X1 U7517 ( .A(n7034), .ZN(n10949) );
  AOI22_X1 U7518 ( .A1(ram[2488]), .A2(n7026), .B1(n10957), .B2(n9054), .ZN(
        n7034) );
  INV_X1 U7519 ( .A(n7035), .ZN(n10950) );
  AOI22_X1 U7520 ( .A1(ram[2489]), .A2(n7026), .B1(n10957), .B2(n9078), .ZN(
        n7035) );
  INV_X1 U7521 ( .A(n7036), .ZN(n10951) );
  AOI22_X1 U7522 ( .A1(ram[2490]), .A2(n7026), .B1(n10957), .B2(n9102), .ZN(
        n7036) );
  INV_X1 U7523 ( .A(n7037), .ZN(n10952) );
  AOI22_X1 U7524 ( .A1(ram[2491]), .A2(n7026), .B1(n10957), .B2(n9126), .ZN(
        n7037) );
  INV_X1 U7525 ( .A(n7038), .ZN(n10953) );
  AOI22_X1 U7526 ( .A1(ram[2492]), .A2(n7026), .B1(n10957), .B2(n9150), .ZN(
        n7038) );
  INV_X1 U7527 ( .A(n7039), .ZN(n10954) );
  AOI22_X1 U7528 ( .A1(ram[2493]), .A2(n7026), .B1(n10957), .B2(n9174), .ZN(
        n7039) );
  INV_X1 U7529 ( .A(n7040), .ZN(n10955) );
  AOI22_X1 U7530 ( .A1(ram[2494]), .A2(n7026), .B1(n10957), .B2(n9198), .ZN(
        n7040) );
  INV_X1 U7531 ( .A(n7041), .ZN(n10956) );
  AOI22_X1 U7532 ( .A1(ram[2495]), .A2(n7026), .B1(n10957), .B2(n9222), .ZN(
        n7041) );
  INV_X1 U7533 ( .A(n7059), .ZN(n10907) );
  AOI22_X1 U7534 ( .A1(ram[2512]), .A2(n7060), .B1(n10923), .B2(n8862), .ZN(
        n7059) );
  INV_X1 U7535 ( .A(n7061), .ZN(n10908) );
  AOI22_X1 U7536 ( .A1(ram[2513]), .A2(n7060), .B1(n10923), .B2(n8886), .ZN(
        n7061) );
  INV_X1 U7537 ( .A(n7062), .ZN(n10909) );
  AOI22_X1 U7538 ( .A1(ram[2514]), .A2(n7060), .B1(n10923), .B2(n8910), .ZN(
        n7062) );
  INV_X1 U7539 ( .A(n7063), .ZN(n10910) );
  AOI22_X1 U7540 ( .A1(ram[2515]), .A2(n7060), .B1(n10923), .B2(n8934), .ZN(
        n7063) );
  INV_X1 U7541 ( .A(n7064), .ZN(n10911) );
  AOI22_X1 U7542 ( .A1(ram[2516]), .A2(n7060), .B1(n10923), .B2(n8958), .ZN(
        n7064) );
  INV_X1 U7543 ( .A(n7065), .ZN(n10912) );
  AOI22_X1 U7544 ( .A1(ram[2517]), .A2(n7060), .B1(n10923), .B2(n8982), .ZN(
        n7065) );
  INV_X1 U7545 ( .A(n7066), .ZN(n10913) );
  AOI22_X1 U7546 ( .A1(ram[2518]), .A2(n7060), .B1(n10923), .B2(n9006), .ZN(
        n7066) );
  INV_X1 U7547 ( .A(n7067), .ZN(n10914) );
  AOI22_X1 U7548 ( .A1(ram[2519]), .A2(n7060), .B1(n10923), .B2(n9030), .ZN(
        n7067) );
  INV_X1 U7549 ( .A(n7068), .ZN(n10915) );
  AOI22_X1 U7550 ( .A1(ram[2520]), .A2(n7060), .B1(n10923), .B2(n9054), .ZN(
        n7068) );
  INV_X1 U7551 ( .A(n7069), .ZN(n10916) );
  AOI22_X1 U7552 ( .A1(ram[2521]), .A2(n7060), .B1(n10923), .B2(n9078), .ZN(
        n7069) );
  INV_X1 U7553 ( .A(n7070), .ZN(n10917) );
  AOI22_X1 U7554 ( .A1(ram[2522]), .A2(n7060), .B1(n10923), .B2(n9102), .ZN(
        n7070) );
  INV_X1 U7555 ( .A(n7071), .ZN(n10918) );
  AOI22_X1 U7556 ( .A1(ram[2523]), .A2(n7060), .B1(n10923), .B2(n9126), .ZN(
        n7071) );
  INV_X1 U7557 ( .A(n7072), .ZN(n10919) );
  AOI22_X1 U7558 ( .A1(ram[2524]), .A2(n7060), .B1(n10923), .B2(n9150), .ZN(
        n7072) );
  INV_X1 U7559 ( .A(n7073), .ZN(n10920) );
  AOI22_X1 U7560 ( .A1(ram[2525]), .A2(n7060), .B1(n10923), .B2(n9174), .ZN(
        n7073) );
  INV_X1 U7561 ( .A(n7074), .ZN(n10921) );
  AOI22_X1 U7562 ( .A1(ram[2526]), .A2(n7060), .B1(n10923), .B2(n9198), .ZN(
        n7074) );
  INV_X1 U7563 ( .A(n7075), .ZN(n10922) );
  AOI22_X1 U7564 ( .A1(ram[2527]), .A2(n7060), .B1(n10923), .B2(n9222), .ZN(
        n7075) );
  INV_X1 U7565 ( .A(n7093), .ZN(n10873) );
  AOI22_X1 U7566 ( .A1(ram[2544]), .A2(n7094), .B1(n10889), .B2(n8862), .ZN(
        n7093) );
  INV_X1 U7567 ( .A(n7095), .ZN(n10874) );
  AOI22_X1 U7568 ( .A1(ram[2545]), .A2(n7094), .B1(n10889), .B2(n8886), .ZN(
        n7095) );
  INV_X1 U7569 ( .A(n7096), .ZN(n10875) );
  AOI22_X1 U7570 ( .A1(ram[2546]), .A2(n7094), .B1(n10889), .B2(n8910), .ZN(
        n7096) );
  INV_X1 U7571 ( .A(n7097), .ZN(n10876) );
  AOI22_X1 U7572 ( .A1(ram[2547]), .A2(n7094), .B1(n10889), .B2(n8934), .ZN(
        n7097) );
  INV_X1 U7573 ( .A(n7098), .ZN(n10877) );
  AOI22_X1 U7574 ( .A1(ram[2548]), .A2(n7094), .B1(n10889), .B2(n8958), .ZN(
        n7098) );
  INV_X1 U7575 ( .A(n7099), .ZN(n10878) );
  AOI22_X1 U7576 ( .A1(ram[2549]), .A2(n7094), .B1(n10889), .B2(n8982), .ZN(
        n7099) );
  INV_X1 U7577 ( .A(n7100), .ZN(n10879) );
  AOI22_X1 U7578 ( .A1(ram[2550]), .A2(n7094), .B1(n10889), .B2(n9006), .ZN(
        n7100) );
  INV_X1 U7579 ( .A(n7101), .ZN(n10880) );
  AOI22_X1 U7580 ( .A1(ram[2551]), .A2(n7094), .B1(n10889), .B2(n9030), .ZN(
        n7101) );
  INV_X1 U7581 ( .A(n7102), .ZN(n10881) );
  AOI22_X1 U7582 ( .A1(ram[2552]), .A2(n7094), .B1(n10889), .B2(n9054), .ZN(
        n7102) );
  INV_X1 U7583 ( .A(n7103), .ZN(n10882) );
  AOI22_X1 U7584 ( .A1(ram[2553]), .A2(n7094), .B1(n10889), .B2(n9078), .ZN(
        n7103) );
  INV_X1 U7585 ( .A(n7104), .ZN(n10883) );
  AOI22_X1 U7586 ( .A1(ram[2554]), .A2(n7094), .B1(n10889), .B2(n9102), .ZN(
        n7104) );
  INV_X1 U7587 ( .A(n7105), .ZN(n10884) );
  AOI22_X1 U7588 ( .A1(ram[2555]), .A2(n7094), .B1(n10889), .B2(n9126), .ZN(
        n7105) );
  INV_X1 U7589 ( .A(n7106), .ZN(n10885) );
  AOI22_X1 U7590 ( .A1(ram[2556]), .A2(n7094), .B1(n10889), .B2(n9150), .ZN(
        n7106) );
  INV_X1 U7591 ( .A(n7107), .ZN(n10886) );
  AOI22_X1 U7592 ( .A1(ram[2557]), .A2(n7094), .B1(n10889), .B2(n9174), .ZN(
        n7107) );
  INV_X1 U7593 ( .A(n7108), .ZN(n10887) );
  AOI22_X1 U7594 ( .A1(ram[2558]), .A2(n7094), .B1(n10889), .B2(n9198), .ZN(
        n7108) );
  INV_X1 U7595 ( .A(n7109), .ZN(n10888) );
  AOI22_X1 U7596 ( .A1(ram[2559]), .A2(n7094), .B1(n10889), .B2(n9222), .ZN(
        n7109) );
  INV_X1 U7597 ( .A(n7128), .ZN(n10839) );
  AOI22_X1 U7598 ( .A1(ram[2576]), .A2(n7129), .B1(n10855), .B2(n8861), .ZN(
        n7128) );
  INV_X1 U7599 ( .A(n7130), .ZN(n10840) );
  AOI22_X1 U7600 ( .A1(ram[2577]), .A2(n7129), .B1(n10855), .B2(n8885), .ZN(
        n7130) );
  INV_X1 U7601 ( .A(n7131), .ZN(n10841) );
  AOI22_X1 U7602 ( .A1(ram[2578]), .A2(n7129), .B1(n10855), .B2(n8909), .ZN(
        n7131) );
  INV_X1 U7603 ( .A(n7132), .ZN(n10842) );
  AOI22_X1 U7604 ( .A1(ram[2579]), .A2(n7129), .B1(n10855), .B2(n8933), .ZN(
        n7132) );
  INV_X1 U7605 ( .A(n7133), .ZN(n10843) );
  AOI22_X1 U7606 ( .A1(ram[2580]), .A2(n7129), .B1(n10855), .B2(n8957), .ZN(
        n7133) );
  INV_X1 U7607 ( .A(n7134), .ZN(n10844) );
  AOI22_X1 U7608 ( .A1(ram[2581]), .A2(n7129), .B1(n10855), .B2(n8981), .ZN(
        n7134) );
  INV_X1 U7609 ( .A(n7135), .ZN(n10845) );
  AOI22_X1 U7610 ( .A1(ram[2582]), .A2(n7129), .B1(n10855), .B2(n9005), .ZN(
        n7135) );
  INV_X1 U7611 ( .A(n7136), .ZN(n10846) );
  AOI22_X1 U7612 ( .A1(ram[2583]), .A2(n7129), .B1(n10855), .B2(n9029), .ZN(
        n7136) );
  INV_X1 U7613 ( .A(n7137), .ZN(n10847) );
  AOI22_X1 U7614 ( .A1(ram[2584]), .A2(n7129), .B1(n10855), .B2(n9053), .ZN(
        n7137) );
  INV_X1 U7615 ( .A(n7138), .ZN(n10848) );
  AOI22_X1 U7616 ( .A1(ram[2585]), .A2(n7129), .B1(n10855), .B2(n9077), .ZN(
        n7138) );
  INV_X1 U7617 ( .A(n7139), .ZN(n10849) );
  AOI22_X1 U7618 ( .A1(ram[2586]), .A2(n7129), .B1(n10855), .B2(n9101), .ZN(
        n7139) );
  INV_X1 U7619 ( .A(n7140), .ZN(n10850) );
  AOI22_X1 U7620 ( .A1(ram[2587]), .A2(n7129), .B1(n10855), .B2(n9125), .ZN(
        n7140) );
  INV_X1 U7621 ( .A(n7141), .ZN(n10851) );
  AOI22_X1 U7622 ( .A1(ram[2588]), .A2(n7129), .B1(n10855), .B2(n9149), .ZN(
        n7141) );
  INV_X1 U7623 ( .A(n7142), .ZN(n10852) );
  AOI22_X1 U7624 ( .A1(ram[2589]), .A2(n7129), .B1(n10855), .B2(n9173), .ZN(
        n7142) );
  INV_X1 U7625 ( .A(n7143), .ZN(n10853) );
  AOI22_X1 U7626 ( .A1(ram[2590]), .A2(n7129), .B1(n10855), .B2(n9197), .ZN(
        n7143) );
  INV_X1 U7627 ( .A(n7144), .ZN(n10854) );
  AOI22_X1 U7628 ( .A1(ram[2591]), .A2(n7129), .B1(n10855), .B2(n9221), .ZN(
        n7144) );
  INV_X1 U7629 ( .A(n7162), .ZN(n10805) );
  AOI22_X1 U7630 ( .A1(ram[2608]), .A2(n7163), .B1(n10821), .B2(n8861), .ZN(
        n7162) );
  INV_X1 U7631 ( .A(n7164), .ZN(n10806) );
  AOI22_X1 U7632 ( .A1(ram[2609]), .A2(n7163), .B1(n10821), .B2(n8885), .ZN(
        n7164) );
  INV_X1 U7633 ( .A(n7165), .ZN(n10807) );
  AOI22_X1 U7634 ( .A1(ram[2610]), .A2(n7163), .B1(n10821), .B2(n8909), .ZN(
        n7165) );
  INV_X1 U7635 ( .A(n7166), .ZN(n10808) );
  AOI22_X1 U7636 ( .A1(ram[2611]), .A2(n7163), .B1(n10821), .B2(n8933), .ZN(
        n7166) );
  INV_X1 U7637 ( .A(n7167), .ZN(n10809) );
  AOI22_X1 U7638 ( .A1(ram[2612]), .A2(n7163), .B1(n10821), .B2(n8957), .ZN(
        n7167) );
  INV_X1 U7639 ( .A(n7168), .ZN(n10810) );
  AOI22_X1 U7640 ( .A1(ram[2613]), .A2(n7163), .B1(n10821), .B2(n8981), .ZN(
        n7168) );
  INV_X1 U7641 ( .A(n7169), .ZN(n10811) );
  AOI22_X1 U7642 ( .A1(ram[2614]), .A2(n7163), .B1(n10821), .B2(n9005), .ZN(
        n7169) );
  INV_X1 U7643 ( .A(n7170), .ZN(n10812) );
  AOI22_X1 U7644 ( .A1(ram[2615]), .A2(n7163), .B1(n10821), .B2(n9029), .ZN(
        n7170) );
  INV_X1 U7645 ( .A(n7171), .ZN(n10813) );
  AOI22_X1 U7646 ( .A1(ram[2616]), .A2(n7163), .B1(n10821), .B2(n9053), .ZN(
        n7171) );
  INV_X1 U7647 ( .A(n7172), .ZN(n10814) );
  AOI22_X1 U7648 ( .A1(ram[2617]), .A2(n7163), .B1(n10821), .B2(n9077), .ZN(
        n7172) );
  INV_X1 U7649 ( .A(n7173), .ZN(n10815) );
  AOI22_X1 U7650 ( .A1(ram[2618]), .A2(n7163), .B1(n10821), .B2(n9101), .ZN(
        n7173) );
  INV_X1 U7651 ( .A(n7174), .ZN(n10816) );
  AOI22_X1 U7652 ( .A1(ram[2619]), .A2(n7163), .B1(n10821), .B2(n9125), .ZN(
        n7174) );
  INV_X1 U7653 ( .A(n7175), .ZN(n10817) );
  AOI22_X1 U7654 ( .A1(ram[2620]), .A2(n7163), .B1(n10821), .B2(n9149), .ZN(
        n7175) );
  INV_X1 U7655 ( .A(n7176), .ZN(n10818) );
  AOI22_X1 U7656 ( .A1(ram[2621]), .A2(n7163), .B1(n10821), .B2(n9173), .ZN(
        n7176) );
  INV_X1 U7657 ( .A(n7177), .ZN(n10819) );
  AOI22_X1 U7658 ( .A1(ram[2622]), .A2(n7163), .B1(n10821), .B2(n9197), .ZN(
        n7177) );
  INV_X1 U7659 ( .A(n7178), .ZN(n10820) );
  AOI22_X1 U7660 ( .A1(ram[2623]), .A2(n7163), .B1(n10821), .B2(n9221), .ZN(
        n7178) );
  INV_X1 U7661 ( .A(n7196), .ZN(n10771) );
  AOI22_X1 U7662 ( .A1(ram[2640]), .A2(n7197), .B1(n10787), .B2(n8861), .ZN(
        n7196) );
  INV_X1 U7663 ( .A(n7198), .ZN(n10772) );
  AOI22_X1 U7664 ( .A1(ram[2641]), .A2(n7197), .B1(n10787), .B2(n8885), .ZN(
        n7198) );
  INV_X1 U7665 ( .A(n7199), .ZN(n10773) );
  AOI22_X1 U7666 ( .A1(ram[2642]), .A2(n7197), .B1(n10787), .B2(n8909), .ZN(
        n7199) );
  INV_X1 U7667 ( .A(n7200), .ZN(n10774) );
  AOI22_X1 U7668 ( .A1(ram[2643]), .A2(n7197), .B1(n10787), .B2(n8933), .ZN(
        n7200) );
  INV_X1 U7669 ( .A(n7201), .ZN(n10775) );
  AOI22_X1 U7670 ( .A1(ram[2644]), .A2(n7197), .B1(n10787), .B2(n8957), .ZN(
        n7201) );
  INV_X1 U7671 ( .A(n7202), .ZN(n10776) );
  AOI22_X1 U7672 ( .A1(ram[2645]), .A2(n7197), .B1(n10787), .B2(n8981), .ZN(
        n7202) );
  INV_X1 U7673 ( .A(n7203), .ZN(n10777) );
  AOI22_X1 U7674 ( .A1(ram[2646]), .A2(n7197), .B1(n10787), .B2(n9005), .ZN(
        n7203) );
  INV_X1 U7675 ( .A(n7204), .ZN(n10778) );
  AOI22_X1 U7676 ( .A1(ram[2647]), .A2(n7197), .B1(n10787), .B2(n9029), .ZN(
        n7204) );
  INV_X1 U7677 ( .A(n7205), .ZN(n10779) );
  AOI22_X1 U7678 ( .A1(ram[2648]), .A2(n7197), .B1(n10787), .B2(n9053), .ZN(
        n7205) );
  INV_X1 U7679 ( .A(n7206), .ZN(n10780) );
  AOI22_X1 U7680 ( .A1(ram[2649]), .A2(n7197), .B1(n10787), .B2(n9077), .ZN(
        n7206) );
  INV_X1 U7681 ( .A(n7207), .ZN(n10781) );
  AOI22_X1 U7682 ( .A1(ram[2650]), .A2(n7197), .B1(n10787), .B2(n9101), .ZN(
        n7207) );
  INV_X1 U7683 ( .A(n7208), .ZN(n10782) );
  AOI22_X1 U7684 ( .A1(ram[2651]), .A2(n7197), .B1(n10787), .B2(n9125), .ZN(
        n7208) );
  INV_X1 U7685 ( .A(n7209), .ZN(n10783) );
  AOI22_X1 U7686 ( .A1(ram[2652]), .A2(n7197), .B1(n10787), .B2(n9149), .ZN(
        n7209) );
  INV_X1 U7687 ( .A(n7210), .ZN(n10784) );
  AOI22_X1 U7688 ( .A1(ram[2653]), .A2(n7197), .B1(n10787), .B2(n9173), .ZN(
        n7210) );
  INV_X1 U7689 ( .A(n7211), .ZN(n10785) );
  AOI22_X1 U7690 ( .A1(ram[2654]), .A2(n7197), .B1(n10787), .B2(n9197), .ZN(
        n7211) );
  INV_X1 U7691 ( .A(n7212), .ZN(n10786) );
  AOI22_X1 U7692 ( .A1(ram[2655]), .A2(n7197), .B1(n10787), .B2(n9221), .ZN(
        n7212) );
  INV_X1 U7693 ( .A(n7230), .ZN(n10737) );
  AOI22_X1 U7694 ( .A1(ram[2672]), .A2(n7231), .B1(n10753), .B2(n8861), .ZN(
        n7230) );
  INV_X1 U7695 ( .A(n7232), .ZN(n10738) );
  AOI22_X1 U7696 ( .A1(ram[2673]), .A2(n7231), .B1(n10753), .B2(n8885), .ZN(
        n7232) );
  INV_X1 U7697 ( .A(n7233), .ZN(n10739) );
  AOI22_X1 U7698 ( .A1(ram[2674]), .A2(n7231), .B1(n10753), .B2(n8909), .ZN(
        n7233) );
  INV_X1 U7699 ( .A(n7234), .ZN(n10740) );
  AOI22_X1 U7700 ( .A1(ram[2675]), .A2(n7231), .B1(n10753), .B2(n8933), .ZN(
        n7234) );
  INV_X1 U7701 ( .A(n7235), .ZN(n10741) );
  AOI22_X1 U7702 ( .A1(ram[2676]), .A2(n7231), .B1(n10753), .B2(n8957), .ZN(
        n7235) );
  INV_X1 U7703 ( .A(n7236), .ZN(n10742) );
  AOI22_X1 U7704 ( .A1(ram[2677]), .A2(n7231), .B1(n10753), .B2(n8981), .ZN(
        n7236) );
  INV_X1 U7705 ( .A(n7237), .ZN(n10743) );
  AOI22_X1 U7706 ( .A1(ram[2678]), .A2(n7231), .B1(n10753), .B2(n9005), .ZN(
        n7237) );
  INV_X1 U7707 ( .A(n7238), .ZN(n10744) );
  AOI22_X1 U7708 ( .A1(ram[2679]), .A2(n7231), .B1(n10753), .B2(n9029), .ZN(
        n7238) );
  INV_X1 U7709 ( .A(n7239), .ZN(n10745) );
  AOI22_X1 U7710 ( .A1(ram[2680]), .A2(n7231), .B1(n10753), .B2(n9053), .ZN(
        n7239) );
  INV_X1 U7711 ( .A(n7240), .ZN(n10746) );
  AOI22_X1 U7712 ( .A1(ram[2681]), .A2(n7231), .B1(n10753), .B2(n9077), .ZN(
        n7240) );
  INV_X1 U7713 ( .A(n7241), .ZN(n10747) );
  AOI22_X1 U7714 ( .A1(ram[2682]), .A2(n7231), .B1(n10753), .B2(n9101), .ZN(
        n7241) );
  INV_X1 U7715 ( .A(n7242), .ZN(n10748) );
  AOI22_X1 U7716 ( .A1(ram[2683]), .A2(n7231), .B1(n10753), .B2(n9125), .ZN(
        n7242) );
  INV_X1 U7717 ( .A(n7243), .ZN(n10749) );
  AOI22_X1 U7718 ( .A1(ram[2684]), .A2(n7231), .B1(n10753), .B2(n9149), .ZN(
        n7243) );
  INV_X1 U7719 ( .A(n7244), .ZN(n10750) );
  AOI22_X1 U7720 ( .A1(ram[2685]), .A2(n7231), .B1(n10753), .B2(n9173), .ZN(
        n7244) );
  INV_X1 U7721 ( .A(n7245), .ZN(n10751) );
  AOI22_X1 U7722 ( .A1(ram[2686]), .A2(n7231), .B1(n10753), .B2(n9197), .ZN(
        n7245) );
  INV_X1 U7723 ( .A(n7246), .ZN(n10752) );
  AOI22_X1 U7724 ( .A1(ram[2687]), .A2(n7231), .B1(n10753), .B2(n9221), .ZN(
        n7246) );
  INV_X1 U7725 ( .A(n7264), .ZN(n10703) );
  AOI22_X1 U7726 ( .A1(ram[2704]), .A2(n7265), .B1(n10719), .B2(n8861), .ZN(
        n7264) );
  INV_X1 U7727 ( .A(n7266), .ZN(n10704) );
  AOI22_X1 U7728 ( .A1(ram[2705]), .A2(n7265), .B1(n10719), .B2(n8885), .ZN(
        n7266) );
  INV_X1 U7729 ( .A(n7267), .ZN(n10705) );
  AOI22_X1 U7730 ( .A1(ram[2706]), .A2(n7265), .B1(n10719), .B2(n8909), .ZN(
        n7267) );
  INV_X1 U7731 ( .A(n7268), .ZN(n10706) );
  AOI22_X1 U7732 ( .A1(ram[2707]), .A2(n7265), .B1(n10719), .B2(n8933), .ZN(
        n7268) );
  INV_X1 U7733 ( .A(n7269), .ZN(n10707) );
  AOI22_X1 U7734 ( .A1(ram[2708]), .A2(n7265), .B1(n10719), .B2(n8957), .ZN(
        n7269) );
  INV_X1 U7735 ( .A(n7270), .ZN(n10708) );
  AOI22_X1 U7736 ( .A1(ram[2709]), .A2(n7265), .B1(n10719), .B2(n8981), .ZN(
        n7270) );
  INV_X1 U7737 ( .A(n7271), .ZN(n10709) );
  AOI22_X1 U7738 ( .A1(ram[2710]), .A2(n7265), .B1(n10719), .B2(n9005), .ZN(
        n7271) );
  INV_X1 U7739 ( .A(n7272), .ZN(n10710) );
  AOI22_X1 U7740 ( .A1(ram[2711]), .A2(n7265), .B1(n10719), .B2(n9029), .ZN(
        n7272) );
  INV_X1 U7741 ( .A(n7273), .ZN(n10711) );
  AOI22_X1 U7742 ( .A1(ram[2712]), .A2(n7265), .B1(n10719), .B2(n9053), .ZN(
        n7273) );
  INV_X1 U7743 ( .A(n7274), .ZN(n10712) );
  AOI22_X1 U7744 ( .A1(ram[2713]), .A2(n7265), .B1(n10719), .B2(n9077), .ZN(
        n7274) );
  INV_X1 U7745 ( .A(n7275), .ZN(n10713) );
  AOI22_X1 U7746 ( .A1(ram[2714]), .A2(n7265), .B1(n10719), .B2(n9101), .ZN(
        n7275) );
  INV_X1 U7747 ( .A(n7276), .ZN(n10714) );
  AOI22_X1 U7748 ( .A1(ram[2715]), .A2(n7265), .B1(n10719), .B2(n9125), .ZN(
        n7276) );
  INV_X1 U7749 ( .A(n7277), .ZN(n10715) );
  AOI22_X1 U7750 ( .A1(ram[2716]), .A2(n7265), .B1(n10719), .B2(n9149), .ZN(
        n7277) );
  INV_X1 U7751 ( .A(n7278), .ZN(n10716) );
  AOI22_X1 U7752 ( .A1(ram[2717]), .A2(n7265), .B1(n10719), .B2(n9173), .ZN(
        n7278) );
  INV_X1 U7753 ( .A(n7279), .ZN(n10717) );
  AOI22_X1 U7754 ( .A1(ram[2718]), .A2(n7265), .B1(n10719), .B2(n9197), .ZN(
        n7279) );
  INV_X1 U7755 ( .A(n7280), .ZN(n10718) );
  AOI22_X1 U7756 ( .A1(ram[2719]), .A2(n7265), .B1(n10719), .B2(n9221), .ZN(
        n7280) );
  INV_X1 U7757 ( .A(n7298), .ZN(n10669) );
  AOI22_X1 U7758 ( .A1(ram[2736]), .A2(n7299), .B1(n10685), .B2(n8861), .ZN(
        n7298) );
  INV_X1 U7759 ( .A(n7300), .ZN(n10670) );
  AOI22_X1 U7760 ( .A1(ram[2737]), .A2(n7299), .B1(n10685), .B2(n8885), .ZN(
        n7300) );
  INV_X1 U7761 ( .A(n7301), .ZN(n10671) );
  AOI22_X1 U7762 ( .A1(ram[2738]), .A2(n7299), .B1(n10685), .B2(n8909), .ZN(
        n7301) );
  INV_X1 U7763 ( .A(n7302), .ZN(n10672) );
  AOI22_X1 U7764 ( .A1(ram[2739]), .A2(n7299), .B1(n10685), .B2(n8933), .ZN(
        n7302) );
  INV_X1 U7765 ( .A(n7303), .ZN(n10673) );
  AOI22_X1 U7766 ( .A1(ram[2740]), .A2(n7299), .B1(n10685), .B2(n8957), .ZN(
        n7303) );
  INV_X1 U7767 ( .A(n7304), .ZN(n10674) );
  AOI22_X1 U7768 ( .A1(ram[2741]), .A2(n7299), .B1(n10685), .B2(n8981), .ZN(
        n7304) );
  INV_X1 U7769 ( .A(n7305), .ZN(n10675) );
  AOI22_X1 U7770 ( .A1(ram[2742]), .A2(n7299), .B1(n10685), .B2(n9005), .ZN(
        n7305) );
  INV_X1 U7771 ( .A(n7306), .ZN(n10676) );
  AOI22_X1 U7772 ( .A1(ram[2743]), .A2(n7299), .B1(n10685), .B2(n9029), .ZN(
        n7306) );
  INV_X1 U7773 ( .A(n7307), .ZN(n10677) );
  AOI22_X1 U7774 ( .A1(ram[2744]), .A2(n7299), .B1(n10685), .B2(n9053), .ZN(
        n7307) );
  INV_X1 U7775 ( .A(n7308), .ZN(n10678) );
  AOI22_X1 U7776 ( .A1(ram[2745]), .A2(n7299), .B1(n10685), .B2(n9077), .ZN(
        n7308) );
  INV_X1 U7777 ( .A(n7309), .ZN(n10679) );
  AOI22_X1 U7778 ( .A1(ram[2746]), .A2(n7299), .B1(n10685), .B2(n9101), .ZN(
        n7309) );
  INV_X1 U7779 ( .A(n7310), .ZN(n10680) );
  AOI22_X1 U7780 ( .A1(ram[2747]), .A2(n7299), .B1(n10685), .B2(n9125), .ZN(
        n7310) );
  INV_X1 U7781 ( .A(n7311), .ZN(n10681) );
  AOI22_X1 U7782 ( .A1(ram[2748]), .A2(n7299), .B1(n10685), .B2(n9149), .ZN(
        n7311) );
  INV_X1 U7783 ( .A(n7312), .ZN(n10682) );
  AOI22_X1 U7784 ( .A1(ram[2749]), .A2(n7299), .B1(n10685), .B2(n9173), .ZN(
        n7312) );
  INV_X1 U7785 ( .A(n7313), .ZN(n10683) );
  AOI22_X1 U7786 ( .A1(ram[2750]), .A2(n7299), .B1(n10685), .B2(n9197), .ZN(
        n7313) );
  INV_X1 U7787 ( .A(n7314), .ZN(n10684) );
  AOI22_X1 U7788 ( .A1(ram[2751]), .A2(n7299), .B1(n10685), .B2(n9221), .ZN(
        n7314) );
  INV_X1 U7789 ( .A(n7332), .ZN(n10635) );
  AOI22_X1 U7790 ( .A1(ram[2768]), .A2(n7333), .B1(n10651), .B2(n8860), .ZN(
        n7332) );
  INV_X1 U7791 ( .A(n7334), .ZN(n10636) );
  AOI22_X1 U7792 ( .A1(ram[2769]), .A2(n7333), .B1(n10651), .B2(n8884), .ZN(
        n7334) );
  INV_X1 U7793 ( .A(n7335), .ZN(n10637) );
  AOI22_X1 U7794 ( .A1(ram[2770]), .A2(n7333), .B1(n10651), .B2(n8908), .ZN(
        n7335) );
  INV_X1 U7795 ( .A(n7336), .ZN(n10638) );
  AOI22_X1 U7796 ( .A1(ram[2771]), .A2(n7333), .B1(n10651), .B2(n8932), .ZN(
        n7336) );
  INV_X1 U7797 ( .A(n7337), .ZN(n10639) );
  AOI22_X1 U7798 ( .A1(ram[2772]), .A2(n7333), .B1(n10651), .B2(n8956), .ZN(
        n7337) );
  INV_X1 U7799 ( .A(n7338), .ZN(n10640) );
  AOI22_X1 U7800 ( .A1(ram[2773]), .A2(n7333), .B1(n10651), .B2(n8980), .ZN(
        n7338) );
  INV_X1 U7801 ( .A(n7339), .ZN(n10641) );
  AOI22_X1 U7802 ( .A1(ram[2774]), .A2(n7333), .B1(n10651), .B2(n9004), .ZN(
        n7339) );
  INV_X1 U7803 ( .A(n7340), .ZN(n10642) );
  AOI22_X1 U7804 ( .A1(ram[2775]), .A2(n7333), .B1(n10651), .B2(n9028), .ZN(
        n7340) );
  INV_X1 U7805 ( .A(n7341), .ZN(n10643) );
  AOI22_X1 U7806 ( .A1(ram[2776]), .A2(n7333), .B1(n10651), .B2(n9052), .ZN(
        n7341) );
  INV_X1 U7807 ( .A(n7342), .ZN(n10644) );
  AOI22_X1 U7808 ( .A1(ram[2777]), .A2(n7333), .B1(n10651), .B2(n9076), .ZN(
        n7342) );
  INV_X1 U7809 ( .A(n7343), .ZN(n10645) );
  AOI22_X1 U7810 ( .A1(ram[2778]), .A2(n7333), .B1(n10651), .B2(n9100), .ZN(
        n7343) );
  INV_X1 U7811 ( .A(n7344), .ZN(n10646) );
  AOI22_X1 U7812 ( .A1(ram[2779]), .A2(n7333), .B1(n10651), .B2(n9124), .ZN(
        n7344) );
  INV_X1 U7813 ( .A(n7345), .ZN(n10647) );
  AOI22_X1 U7814 ( .A1(ram[2780]), .A2(n7333), .B1(n10651), .B2(n9148), .ZN(
        n7345) );
  INV_X1 U7815 ( .A(n7346), .ZN(n10648) );
  AOI22_X1 U7816 ( .A1(ram[2781]), .A2(n7333), .B1(n10651), .B2(n9172), .ZN(
        n7346) );
  INV_X1 U7817 ( .A(n7347), .ZN(n10649) );
  AOI22_X1 U7818 ( .A1(ram[2782]), .A2(n7333), .B1(n10651), .B2(n9196), .ZN(
        n7347) );
  INV_X1 U7819 ( .A(n7348), .ZN(n10650) );
  AOI22_X1 U7820 ( .A1(ram[2783]), .A2(n7333), .B1(n10651), .B2(n9220), .ZN(
        n7348) );
  INV_X1 U7821 ( .A(n7366), .ZN(n10601) );
  AOI22_X1 U7822 ( .A1(ram[2800]), .A2(n7367), .B1(n10617), .B2(n8860), .ZN(
        n7366) );
  INV_X1 U7823 ( .A(n7368), .ZN(n10602) );
  AOI22_X1 U7824 ( .A1(ram[2801]), .A2(n7367), .B1(n10617), .B2(n8884), .ZN(
        n7368) );
  INV_X1 U7825 ( .A(n7369), .ZN(n10603) );
  AOI22_X1 U7826 ( .A1(ram[2802]), .A2(n7367), .B1(n10617), .B2(n8908), .ZN(
        n7369) );
  INV_X1 U7827 ( .A(n7370), .ZN(n10604) );
  AOI22_X1 U7828 ( .A1(ram[2803]), .A2(n7367), .B1(n10617), .B2(n8932), .ZN(
        n7370) );
  INV_X1 U7829 ( .A(n7371), .ZN(n10605) );
  AOI22_X1 U7830 ( .A1(ram[2804]), .A2(n7367), .B1(n10617), .B2(n8956), .ZN(
        n7371) );
  INV_X1 U7831 ( .A(n7372), .ZN(n10606) );
  AOI22_X1 U7832 ( .A1(ram[2805]), .A2(n7367), .B1(n10617), .B2(n8980), .ZN(
        n7372) );
  INV_X1 U7833 ( .A(n7373), .ZN(n10607) );
  AOI22_X1 U7834 ( .A1(ram[2806]), .A2(n7367), .B1(n10617), .B2(n9004), .ZN(
        n7373) );
  INV_X1 U7835 ( .A(n7374), .ZN(n10608) );
  AOI22_X1 U7836 ( .A1(ram[2807]), .A2(n7367), .B1(n10617), .B2(n9028), .ZN(
        n7374) );
  INV_X1 U7837 ( .A(n7375), .ZN(n10609) );
  AOI22_X1 U7838 ( .A1(ram[2808]), .A2(n7367), .B1(n10617), .B2(n9052), .ZN(
        n7375) );
  INV_X1 U7839 ( .A(n7376), .ZN(n10610) );
  AOI22_X1 U7840 ( .A1(ram[2809]), .A2(n7367), .B1(n10617), .B2(n9076), .ZN(
        n7376) );
  INV_X1 U7841 ( .A(n7377), .ZN(n10611) );
  AOI22_X1 U7842 ( .A1(ram[2810]), .A2(n7367), .B1(n10617), .B2(n9100), .ZN(
        n7377) );
  INV_X1 U7843 ( .A(n7378), .ZN(n10612) );
  AOI22_X1 U7844 ( .A1(ram[2811]), .A2(n7367), .B1(n10617), .B2(n9124), .ZN(
        n7378) );
  INV_X1 U7845 ( .A(n7379), .ZN(n10613) );
  AOI22_X1 U7846 ( .A1(ram[2812]), .A2(n7367), .B1(n10617), .B2(n9148), .ZN(
        n7379) );
  INV_X1 U7847 ( .A(n7380), .ZN(n10614) );
  AOI22_X1 U7848 ( .A1(ram[2813]), .A2(n7367), .B1(n10617), .B2(n9172), .ZN(
        n7380) );
  INV_X1 U7849 ( .A(n7381), .ZN(n10615) );
  AOI22_X1 U7850 ( .A1(ram[2814]), .A2(n7367), .B1(n10617), .B2(n9196), .ZN(
        n7381) );
  INV_X1 U7851 ( .A(n7382), .ZN(n10616) );
  AOI22_X1 U7852 ( .A1(ram[2815]), .A2(n7367), .B1(n10617), .B2(n9220), .ZN(
        n7382) );
  INV_X1 U7853 ( .A(n7401), .ZN(n10567) );
  AOI22_X1 U7854 ( .A1(ram[2832]), .A2(n7402), .B1(n10583), .B2(n8860), .ZN(
        n7401) );
  INV_X1 U7855 ( .A(n7403), .ZN(n10568) );
  AOI22_X1 U7856 ( .A1(ram[2833]), .A2(n7402), .B1(n10583), .B2(n8884), .ZN(
        n7403) );
  INV_X1 U7857 ( .A(n7404), .ZN(n10569) );
  AOI22_X1 U7858 ( .A1(ram[2834]), .A2(n7402), .B1(n10583), .B2(n8908), .ZN(
        n7404) );
  INV_X1 U7859 ( .A(n7405), .ZN(n10570) );
  AOI22_X1 U7860 ( .A1(ram[2835]), .A2(n7402), .B1(n10583), .B2(n8932), .ZN(
        n7405) );
  INV_X1 U7861 ( .A(n7406), .ZN(n10571) );
  AOI22_X1 U7862 ( .A1(ram[2836]), .A2(n7402), .B1(n10583), .B2(n8956), .ZN(
        n7406) );
  INV_X1 U7863 ( .A(n7407), .ZN(n10572) );
  AOI22_X1 U7864 ( .A1(ram[2837]), .A2(n7402), .B1(n10583), .B2(n8980), .ZN(
        n7407) );
  INV_X1 U7865 ( .A(n7408), .ZN(n10573) );
  AOI22_X1 U7866 ( .A1(ram[2838]), .A2(n7402), .B1(n10583), .B2(n9004), .ZN(
        n7408) );
  INV_X1 U7867 ( .A(n7409), .ZN(n10574) );
  AOI22_X1 U7868 ( .A1(ram[2839]), .A2(n7402), .B1(n10583), .B2(n9028), .ZN(
        n7409) );
  INV_X1 U7869 ( .A(n7410), .ZN(n10575) );
  AOI22_X1 U7870 ( .A1(ram[2840]), .A2(n7402), .B1(n10583), .B2(n9052), .ZN(
        n7410) );
  INV_X1 U7871 ( .A(n7411), .ZN(n10576) );
  AOI22_X1 U7872 ( .A1(ram[2841]), .A2(n7402), .B1(n10583), .B2(n9076), .ZN(
        n7411) );
  INV_X1 U7873 ( .A(n7412), .ZN(n10577) );
  AOI22_X1 U7874 ( .A1(ram[2842]), .A2(n7402), .B1(n10583), .B2(n9100), .ZN(
        n7412) );
  INV_X1 U7875 ( .A(n7413), .ZN(n10578) );
  AOI22_X1 U7876 ( .A1(ram[2843]), .A2(n7402), .B1(n10583), .B2(n9124), .ZN(
        n7413) );
  INV_X1 U7877 ( .A(n7414), .ZN(n10579) );
  AOI22_X1 U7878 ( .A1(ram[2844]), .A2(n7402), .B1(n10583), .B2(n9148), .ZN(
        n7414) );
  INV_X1 U7879 ( .A(n7415), .ZN(n10580) );
  AOI22_X1 U7880 ( .A1(ram[2845]), .A2(n7402), .B1(n10583), .B2(n9172), .ZN(
        n7415) );
  INV_X1 U7881 ( .A(n7416), .ZN(n10581) );
  AOI22_X1 U7882 ( .A1(ram[2846]), .A2(n7402), .B1(n10583), .B2(n9196), .ZN(
        n7416) );
  INV_X1 U7883 ( .A(n7417), .ZN(n10582) );
  AOI22_X1 U7884 ( .A1(ram[2847]), .A2(n7402), .B1(n10583), .B2(n9220), .ZN(
        n7417) );
  INV_X1 U7885 ( .A(n7435), .ZN(n10533) );
  AOI22_X1 U7886 ( .A1(ram[2864]), .A2(n7436), .B1(n10549), .B2(n8860), .ZN(
        n7435) );
  INV_X1 U7887 ( .A(n7437), .ZN(n10534) );
  AOI22_X1 U7888 ( .A1(ram[2865]), .A2(n7436), .B1(n10549), .B2(n8884), .ZN(
        n7437) );
  INV_X1 U7889 ( .A(n7438), .ZN(n10535) );
  AOI22_X1 U7890 ( .A1(ram[2866]), .A2(n7436), .B1(n10549), .B2(n8908), .ZN(
        n7438) );
  INV_X1 U7891 ( .A(n7439), .ZN(n10536) );
  AOI22_X1 U7892 ( .A1(ram[2867]), .A2(n7436), .B1(n10549), .B2(n8932), .ZN(
        n7439) );
  INV_X1 U7893 ( .A(n7440), .ZN(n10537) );
  AOI22_X1 U7894 ( .A1(ram[2868]), .A2(n7436), .B1(n10549), .B2(n8956), .ZN(
        n7440) );
  INV_X1 U7895 ( .A(n7441), .ZN(n10538) );
  AOI22_X1 U7896 ( .A1(ram[2869]), .A2(n7436), .B1(n10549), .B2(n8980), .ZN(
        n7441) );
  INV_X1 U7897 ( .A(n7442), .ZN(n10539) );
  AOI22_X1 U7898 ( .A1(ram[2870]), .A2(n7436), .B1(n10549), .B2(n9004), .ZN(
        n7442) );
  INV_X1 U7899 ( .A(n7443), .ZN(n10540) );
  AOI22_X1 U7900 ( .A1(ram[2871]), .A2(n7436), .B1(n10549), .B2(n9028), .ZN(
        n7443) );
  INV_X1 U7901 ( .A(n7444), .ZN(n10541) );
  AOI22_X1 U7902 ( .A1(ram[2872]), .A2(n7436), .B1(n10549), .B2(n9052), .ZN(
        n7444) );
  INV_X1 U7903 ( .A(n7445), .ZN(n10542) );
  AOI22_X1 U7904 ( .A1(ram[2873]), .A2(n7436), .B1(n10549), .B2(n9076), .ZN(
        n7445) );
  INV_X1 U7905 ( .A(n7446), .ZN(n10543) );
  AOI22_X1 U7906 ( .A1(ram[2874]), .A2(n7436), .B1(n10549), .B2(n9100), .ZN(
        n7446) );
  INV_X1 U7907 ( .A(n7447), .ZN(n10544) );
  AOI22_X1 U7908 ( .A1(ram[2875]), .A2(n7436), .B1(n10549), .B2(n9124), .ZN(
        n7447) );
  INV_X1 U7909 ( .A(n7448), .ZN(n10545) );
  AOI22_X1 U7910 ( .A1(ram[2876]), .A2(n7436), .B1(n10549), .B2(n9148), .ZN(
        n7448) );
  INV_X1 U7911 ( .A(n7449), .ZN(n10546) );
  AOI22_X1 U7912 ( .A1(ram[2877]), .A2(n7436), .B1(n10549), .B2(n9172), .ZN(
        n7449) );
  INV_X1 U7913 ( .A(n7450), .ZN(n10547) );
  AOI22_X1 U7914 ( .A1(ram[2878]), .A2(n7436), .B1(n10549), .B2(n9196), .ZN(
        n7450) );
  INV_X1 U7915 ( .A(n7451), .ZN(n10548) );
  AOI22_X1 U7916 ( .A1(ram[2879]), .A2(n7436), .B1(n10549), .B2(n9220), .ZN(
        n7451) );
  INV_X1 U7917 ( .A(n7469), .ZN(n10499) );
  AOI22_X1 U7918 ( .A1(ram[2896]), .A2(n7470), .B1(n10515), .B2(n8860), .ZN(
        n7469) );
  INV_X1 U7919 ( .A(n7471), .ZN(n10500) );
  AOI22_X1 U7920 ( .A1(ram[2897]), .A2(n7470), .B1(n10515), .B2(n8884), .ZN(
        n7471) );
  INV_X1 U7921 ( .A(n7472), .ZN(n10501) );
  AOI22_X1 U7922 ( .A1(ram[2898]), .A2(n7470), .B1(n10515), .B2(n8908), .ZN(
        n7472) );
  INV_X1 U7923 ( .A(n7473), .ZN(n10502) );
  AOI22_X1 U7924 ( .A1(ram[2899]), .A2(n7470), .B1(n10515), .B2(n8932), .ZN(
        n7473) );
  INV_X1 U7925 ( .A(n7474), .ZN(n10503) );
  AOI22_X1 U7926 ( .A1(ram[2900]), .A2(n7470), .B1(n10515), .B2(n8956), .ZN(
        n7474) );
  INV_X1 U7927 ( .A(n7475), .ZN(n10504) );
  AOI22_X1 U7928 ( .A1(ram[2901]), .A2(n7470), .B1(n10515), .B2(n8980), .ZN(
        n7475) );
  INV_X1 U7929 ( .A(n7476), .ZN(n10505) );
  AOI22_X1 U7930 ( .A1(ram[2902]), .A2(n7470), .B1(n10515), .B2(n9004), .ZN(
        n7476) );
  INV_X1 U7931 ( .A(n7477), .ZN(n10506) );
  AOI22_X1 U7932 ( .A1(ram[2903]), .A2(n7470), .B1(n10515), .B2(n9028), .ZN(
        n7477) );
  INV_X1 U7933 ( .A(n7478), .ZN(n10507) );
  AOI22_X1 U7934 ( .A1(ram[2904]), .A2(n7470), .B1(n10515), .B2(n9052), .ZN(
        n7478) );
  INV_X1 U7935 ( .A(n7479), .ZN(n10508) );
  AOI22_X1 U7936 ( .A1(ram[2905]), .A2(n7470), .B1(n10515), .B2(n9076), .ZN(
        n7479) );
  INV_X1 U7937 ( .A(n7480), .ZN(n10509) );
  AOI22_X1 U7938 ( .A1(ram[2906]), .A2(n7470), .B1(n10515), .B2(n9100), .ZN(
        n7480) );
  INV_X1 U7939 ( .A(n7481), .ZN(n10510) );
  AOI22_X1 U7940 ( .A1(ram[2907]), .A2(n7470), .B1(n10515), .B2(n9124), .ZN(
        n7481) );
  INV_X1 U7941 ( .A(n7482), .ZN(n10511) );
  AOI22_X1 U7942 ( .A1(ram[2908]), .A2(n7470), .B1(n10515), .B2(n9148), .ZN(
        n7482) );
  INV_X1 U7943 ( .A(n7483), .ZN(n10512) );
  AOI22_X1 U7944 ( .A1(ram[2909]), .A2(n7470), .B1(n10515), .B2(n9172), .ZN(
        n7483) );
  INV_X1 U7945 ( .A(n7484), .ZN(n10513) );
  AOI22_X1 U7946 ( .A1(ram[2910]), .A2(n7470), .B1(n10515), .B2(n9196), .ZN(
        n7484) );
  INV_X1 U7947 ( .A(n7485), .ZN(n10514) );
  AOI22_X1 U7948 ( .A1(ram[2911]), .A2(n7470), .B1(n10515), .B2(n9220), .ZN(
        n7485) );
  INV_X1 U7949 ( .A(n7503), .ZN(n10465) );
  AOI22_X1 U7950 ( .A1(ram[2928]), .A2(n7504), .B1(n10481), .B2(n8860), .ZN(
        n7503) );
  INV_X1 U7951 ( .A(n7505), .ZN(n10466) );
  AOI22_X1 U7952 ( .A1(ram[2929]), .A2(n7504), .B1(n10481), .B2(n8884), .ZN(
        n7505) );
  INV_X1 U7953 ( .A(n7506), .ZN(n10467) );
  AOI22_X1 U7954 ( .A1(ram[2930]), .A2(n7504), .B1(n10481), .B2(n8908), .ZN(
        n7506) );
  INV_X1 U7955 ( .A(n7507), .ZN(n10468) );
  AOI22_X1 U7956 ( .A1(ram[2931]), .A2(n7504), .B1(n10481), .B2(n8932), .ZN(
        n7507) );
  INV_X1 U7957 ( .A(n7508), .ZN(n10469) );
  AOI22_X1 U7958 ( .A1(ram[2932]), .A2(n7504), .B1(n10481), .B2(n8956), .ZN(
        n7508) );
  INV_X1 U7959 ( .A(n7509), .ZN(n10470) );
  AOI22_X1 U7960 ( .A1(ram[2933]), .A2(n7504), .B1(n10481), .B2(n8980), .ZN(
        n7509) );
  INV_X1 U7961 ( .A(n7510), .ZN(n10471) );
  AOI22_X1 U7962 ( .A1(ram[2934]), .A2(n7504), .B1(n10481), .B2(n9004), .ZN(
        n7510) );
  INV_X1 U7963 ( .A(n7511), .ZN(n10472) );
  AOI22_X1 U7964 ( .A1(ram[2935]), .A2(n7504), .B1(n10481), .B2(n9028), .ZN(
        n7511) );
  INV_X1 U7965 ( .A(n7512), .ZN(n10473) );
  AOI22_X1 U7966 ( .A1(ram[2936]), .A2(n7504), .B1(n10481), .B2(n9052), .ZN(
        n7512) );
  INV_X1 U7967 ( .A(n7513), .ZN(n10474) );
  AOI22_X1 U7968 ( .A1(ram[2937]), .A2(n7504), .B1(n10481), .B2(n9076), .ZN(
        n7513) );
  INV_X1 U7969 ( .A(n7514), .ZN(n10475) );
  AOI22_X1 U7970 ( .A1(ram[2938]), .A2(n7504), .B1(n10481), .B2(n9100), .ZN(
        n7514) );
  INV_X1 U7971 ( .A(n7515), .ZN(n10476) );
  AOI22_X1 U7972 ( .A1(ram[2939]), .A2(n7504), .B1(n10481), .B2(n9124), .ZN(
        n7515) );
  INV_X1 U7973 ( .A(n7516), .ZN(n10477) );
  AOI22_X1 U7974 ( .A1(ram[2940]), .A2(n7504), .B1(n10481), .B2(n9148), .ZN(
        n7516) );
  INV_X1 U7975 ( .A(n7517), .ZN(n10478) );
  AOI22_X1 U7976 ( .A1(ram[2941]), .A2(n7504), .B1(n10481), .B2(n9172), .ZN(
        n7517) );
  INV_X1 U7977 ( .A(n7518), .ZN(n10479) );
  AOI22_X1 U7978 ( .A1(ram[2942]), .A2(n7504), .B1(n10481), .B2(n9196), .ZN(
        n7518) );
  INV_X1 U7979 ( .A(n7519), .ZN(n10480) );
  AOI22_X1 U7980 ( .A1(ram[2943]), .A2(n7504), .B1(n10481), .B2(n9220), .ZN(
        n7519) );
  INV_X1 U7981 ( .A(n7537), .ZN(n10431) );
  AOI22_X1 U7982 ( .A1(ram[2960]), .A2(n7538), .B1(n10447), .B2(n8859), .ZN(
        n7537) );
  INV_X1 U7983 ( .A(n7539), .ZN(n10432) );
  AOI22_X1 U7984 ( .A1(ram[2961]), .A2(n7538), .B1(n10447), .B2(n8883), .ZN(
        n7539) );
  INV_X1 U7985 ( .A(n7540), .ZN(n10433) );
  AOI22_X1 U7986 ( .A1(ram[2962]), .A2(n7538), .B1(n10447), .B2(n8907), .ZN(
        n7540) );
  INV_X1 U7987 ( .A(n7541), .ZN(n10434) );
  AOI22_X1 U7988 ( .A1(ram[2963]), .A2(n7538), .B1(n10447), .B2(n8931), .ZN(
        n7541) );
  INV_X1 U7989 ( .A(n7542), .ZN(n10435) );
  AOI22_X1 U7990 ( .A1(ram[2964]), .A2(n7538), .B1(n10447), .B2(n8955), .ZN(
        n7542) );
  INV_X1 U7991 ( .A(n7543), .ZN(n10436) );
  AOI22_X1 U7992 ( .A1(ram[2965]), .A2(n7538), .B1(n10447), .B2(n8979), .ZN(
        n7543) );
  INV_X1 U7993 ( .A(n7544), .ZN(n10437) );
  AOI22_X1 U7994 ( .A1(ram[2966]), .A2(n7538), .B1(n10447), .B2(n9003), .ZN(
        n7544) );
  INV_X1 U7995 ( .A(n7545), .ZN(n10438) );
  AOI22_X1 U7996 ( .A1(ram[2967]), .A2(n7538), .B1(n10447), .B2(n9027), .ZN(
        n7545) );
  INV_X1 U7997 ( .A(n7546), .ZN(n10439) );
  AOI22_X1 U7998 ( .A1(ram[2968]), .A2(n7538), .B1(n10447), .B2(n9051), .ZN(
        n7546) );
  INV_X1 U7999 ( .A(n7547), .ZN(n10440) );
  AOI22_X1 U8000 ( .A1(ram[2969]), .A2(n7538), .B1(n10447), .B2(n9075), .ZN(
        n7547) );
  INV_X1 U8001 ( .A(n7548), .ZN(n10441) );
  AOI22_X1 U8002 ( .A1(ram[2970]), .A2(n7538), .B1(n10447), .B2(n9099), .ZN(
        n7548) );
  INV_X1 U8003 ( .A(n7549), .ZN(n10442) );
  AOI22_X1 U8004 ( .A1(ram[2971]), .A2(n7538), .B1(n10447), .B2(n9123), .ZN(
        n7549) );
  INV_X1 U8005 ( .A(n7550), .ZN(n10443) );
  AOI22_X1 U8006 ( .A1(ram[2972]), .A2(n7538), .B1(n10447), .B2(n9147), .ZN(
        n7550) );
  INV_X1 U8007 ( .A(n7551), .ZN(n10444) );
  AOI22_X1 U8008 ( .A1(ram[2973]), .A2(n7538), .B1(n10447), .B2(n9171), .ZN(
        n7551) );
  INV_X1 U8009 ( .A(n7552), .ZN(n10445) );
  AOI22_X1 U8010 ( .A1(ram[2974]), .A2(n7538), .B1(n10447), .B2(n9195), .ZN(
        n7552) );
  INV_X1 U8011 ( .A(n7553), .ZN(n10446) );
  AOI22_X1 U8012 ( .A1(ram[2975]), .A2(n7538), .B1(n10447), .B2(n9219), .ZN(
        n7553) );
  INV_X1 U8013 ( .A(n7571), .ZN(n10397) );
  AOI22_X1 U8014 ( .A1(ram[2992]), .A2(n7572), .B1(n10413), .B2(n8859), .ZN(
        n7571) );
  INV_X1 U8015 ( .A(n7573), .ZN(n10398) );
  AOI22_X1 U8016 ( .A1(ram[2993]), .A2(n7572), .B1(n10413), .B2(n8883), .ZN(
        n7573) );
  INV_X1 U8017 ( .A(n7574), .ZN(n10399) );
  AOI22_X1 U8018 ( .A1(ram[2994]), .A2(n7572), .B1(n10413), .B2(n8907), .ZN(
        n7574) );
  INV_X1 U8019 ( .A(n7575), .ZN(n10400) );
  AOI22_X1 U8020 ( .A1(ram[2995]), .A2(n7572), .B1(n10413), .B2(n8931), .ZN(
        n7575) );
  INV_X1 U8021 ( .A(n7576), .ZN(n10401) );
  AOI22_X1 U8022 ( .A1(ram[2996]), .A2(n7572), .B1(n10413), .B2(n8955), .ZN(
        n7576) );
  INV_X1 U8023 ( .A(n7577), .ZN(n10402) );
  AOI22_X1 U8024 ( .A1(ram[2997]), .A2(n7572), .B1(n10413), .B2(n8979), .ZN(
        n7577) );
  INV_X1 U8025 ( .A(n7578), .ZN(n10403) );
  AOI22_X1 U8026 ( .A1(ram[2998]), .A2(n7572), .B1(n10413), .B2(n9003), .ZN(
        n7578) );
  INV_X1 U8027 ( .A(n7579), .ZN(n10404) );
  AOI22_X1 U8028 ( .A1(ram[2999]), .A2(n7572), .B1(n10413), .B2(n9027), .ZN(
        n7579) );
  INV_X1 U8029 ( .A(n7580), .ZN(n10405) );
  AOI22_X1 U8030 ( .A1(ram[3000]), .A2(n7572), .B1(n10413), .B2(n9051), .ZN(
        n7580) );
  INV_X1 U8031 ( .A(n7581), .ZN(n10406) );
  AOI22_X1 U8032 ( .A1(ram[3001]), .A2(n7572), .B1(n10413), .B2(n9075), .ZN(
        n7581) );
  INV_X1 U8033 ( .A(n7582), .ZN(n10407) );
  AOI22_X1 U8034 ( .A1(ram[3002]), .A2(n7572), .B1(n10413), .B2(n9099), .ZN(
        n7582) );
  INV_X1 U8035 ( .A(n7583), .ZN(n10408) );
  AOI22_X1 U8036 ( .A1(ram[3003]), .A2(n7572), .B1(n10413), .B2(n9123), .ZN(
        n7583) );
  INV_X1 U8037 ( .A(n7584), .ZN(n10409) );
  AOI22_X1 U8038 ( .A1(ram[3004]), .A2(n7572), .B1(n10413), .B2(n9147), .ZN(
        n7584) );
  INV_X1 U8039 ( .A(n7585), .ZN(n10410) );
  AOI22_X1 U8040 ( .A1(ram[3005]), .A2(n7572), .B1(n10413), .B2(n9171), .ZN(
        n7585) );
  INV_X1 U8041 ( .A(n7586), .ZN(n10411) );
  AOI22_X1 U8042 ( .A1(ram[3006]), .A2(n7572), .B1(n10413), .B2(n9195), .ZN(
        n7586) );
  INV_X1 U8043 ( .A(n7587), .ZN(n10412) );
  AOI22_X1 U8044 ( .A1(ram[3007]), .A2(n7572), .B1(n10413), .B2(n9219), .ZN(
        n7587) );
  INV_X1 U8045 ( .A(n7605), .ZN(n10363) );
  AOI22_X1 U8046 ( .A1(ram[3024]), .A2(n7606), .B1(n10379), .B2(n8859), .ZN(
        n7605) );
  INV_X1 U8047 ( .A(n7607), .ZN(n10364) );
  AOI22_X1 U8048 ( .A1(ram[3025]), .A2(n7606), .B1(n10379), .B2(n8883), .ZN(
        n7607) );
  INV_X1 U8049 ( .A(n7608), .ZN(n10365) );
  AOI22_X1 U8050 ( .A1(ram[3026]), .A2(n7606), .B1(n10379), .B2(n8907), .ZN(
        n7608) );
  INV_X1 U8051 ( .A(n7609), .ZN(n10366) );
  AOI22_X1 U8052 ( .A1(ram[3027]), .A2(n7606), .B1(n10379), .B2(n8931), .ZN(
        n7609) );
  INV_X1 U8053 ( .A(n7610), .ZN(n10367) );
  AOI22_X1 U8054 ( .A1(ram[3028]), .A2(n7606), .B1(n10379), .B2(n8955), .ZN(
        n7610) );
  INV_X1 U8055 ( .A(n7611), .ZN(n10368) );
  AOI22_X1 U8056 ( .A1(ram[3029]), .A2(n7606), .B1(n10379), .B2(n8979), .ZN(
        n7611) );
  INV_X1 U8057 ( .A(n7612), .ZN(n10369) );
  AOI22_X1 U8058 ( .A1(ram[3030]), .A2(n7606), .B1(n10379), .B2(n9003), .ZN(
        n7612) );
  INV_X1 U8059 ( .A(n7613), .ZN(n10370) );
  AOI22_X1 U8060 ( .A1(ram[3031]), .A2(n7606), .B1(n10379), .B2(n9027), .ZN(
        n7613) );
  INV_X1 U8061 ( .A(n7614), .ZN(n10371) );
  AOI22_X1 U8062 ( .A1(ram[3032]), .A2(n7606), .B1(n10379), .B2(n9051), .ZN(
        n7614) );
  INV_X1 U8063 ( .A(n7615), .ZN(n10372) );
  AOI22_X1 U8064 ( .A1(ram[3033]), .A2(n7606), .B1(n10379), .B2(n9075), .ZN(
        n7615) );
  INV_X1 U8065 ( .A(n7616), .ZN(n10373) );
  AOI22_X1 U8066 ( .A1(ram[3034]), .A2(n7606), .B1(n10379), .B2(n9099), .ZN(
        n7616) );
  INV_X1 U8067 ( .A(n7617), .ZN(n10374) );
  AOI22_X1 U8068 ( .A1(ram[3035]), .A2(n7606), .B1(n10379), .B2(n9123), .ZN(
        n7617) );
  INV_X1 U8069 ( .A(n7618), .ZN(n10375) );
  AOI22_X1 U8070 ( .A1(ram[3036]), .A2(n7606), .B1(n10379), .B2(n9147), .ZN(
        n7618) );
  INV_X1 U8071 ( .A(n7619), .ZN(n10376) );
  AOI22_X1 U8072 ( .A1(ram[3037]), .A2(n7606), .B1(n10379), .B2(n9171), .ZN(
        n7619) );
  INV_X1 U8073 ( .A(n7620), .ZN(n10377) );
  AOI22_X1 U8074 ( .A1(ram[3038]), .A2(n7606), .B1(n10379), .B2(n9195), .ZN(
        n7620) );
  INV_X1 U8075 ( .A(n7621), .ZN(n10378) );
  AOI22_X1 U8076 ( .A1(ram[3039]), .A2(n7606), .B1(n10379), .B2(n9219), .ZN(
        n7621) );
  INV_X1 U8077 ( .A(n7639), .ZN(n10329) );
  AOI22_X1 U8078 ( .A1(ram[3056]), .A2(n7640), .B1(n10345), .B2(n8859), .ZN(
        n7639) );
  INV_X1 U8079 ( .A(n7641), .ZN(n10330) );
  AOI22_X1 U8080 ( .A1(ram[3057]), .A2(n7640), .B1(n10345), .B2(n8883), .ZN(
        n7641) );
  INV_X1 U8081 ( .A(n7642), .ZN(n10331) );
  AOI22_X1 U8082 ( .A1(ram[3058]), .A2(n7640), .B1(n10345), .B2(n8907), .ZN(
        n7642) );
  INV_X1 U8083 ( .A(n7643), .ZN(n10332) );
  AOI22_X1 U8084 ( .A1(ram[3059]), .A2(n7640), .B1(n10345), .B2(n8931), .ZN(
        n7643) );
  INV_X1 U8085 ( .A(n7644), .ZN(n10333) );
  AOI22_X1 U8086 ( .A1(ram[3060]), .A2(n7640), .B1(n10345), .B2(n8955), .ZN(
        n7644) );
  INV_X1 U8087 ( .A(n7645), .ZN(n10334) );
  AOI22_X1 U8088 ( .A1(ram[3061]), .A2(n7640), .B1(n10345), .B2(n8979), .ZN(
        n7645) );
  INV_X1 U8089 ( .A(n7646), .ZN(n10335) );
  AOI22_X1 U8090 ( .A1(ram[3062]), .A2(n7640), .B1(n10345), .B2(n9003), .ZN(
        n7646) );
  INV_X1 U8091 ( .A(n7647), .ZN(n10336) );
  AOI22_X1 U8092 ( .A1(ram[3063]), .A2(n7640), .B1(n10345), .B2(n9027), .ZN(
        n7647) );
  INV_X1 U8093 ( .A(n7648), .ZN(n10337) );
  AOI22_X1 U8094 ( .A1(ram[3064]), .A2(n7640), .B1(n10345), .B2(n9051), .ZN(
        n7648) );
  INV_X1 U8095 ( .A(n7649), .ZN(n10338) );
  AOI22_X1 U8096 ( .A1(ram[3065]), .A2(n7640), .B1(n10345), .B2(n9075), .ZN(
        n7649) );
  INV_X1 U8097 ( .A(n7650), .ZN(n10339) );
  AOI22_X1 U8098 ( .A1(ram[3066]), .A2(n7640), .B1(n10345), .B2(n9099), .ZN(
        n7650) );
  INV_X1 U8099 ( .A(n7651), .ZN(n10340) );
  AOI22_X1 U8100 ( .A1(ram[3067]), .A2(n7640), .B1(n10345), .B2(n9123), .ZN(
        n7651) );
  INV_X1 U8101 ( .A(n7652), .ZN(n10341) );
  AOI22_X1 U8102 ( .A1(ram[3068]), .A2(n7640), .B1(n10345), .B2(n9147), .ZN(
        n7652) );
  INV_X1 U8103 ( .A(n7653), .ZN(n10342) );
  AOI22_X1 U8104 ( .A1(ram[3069]), .A2(n7640), .B1(n10345), .B2(n9171), .ZN(
        n7653) );
  INV_X1 U8105 ( .A(n7654), .ZN(n10343) );
  AOI22_X1 U8106 ( .A1(ram[3070]), .A2(n7640), .B1(n10345), .B2(n9195), .ZN(
        n7654) );
  INV_X1 U8107 ( .A(n7655), .ZN(n10344) );
  AOI22_X1 U8108 ( .A1(ram[3071]), .A2(n7640), .B1(n10345), .B2(n9219), .ZN(
        n7655) );
  INV_X1 U8109 ( .A(n7674), .ZN(n10295) );
  AOI22_X1 U8110 ( .A1(ram[3088]), .A2(n7675), .B1(n10311), .B2(n8859), .ZN(
        n7674) );
  INV_X1 U8111 ( .A(n7676), .ZN(n10296) );
  AOI22_X1 U8112 ( .A1(ram[3089]), .A2(n7675), .B1(n10311), .B2(n8883), .ZN(
        n7676) );
  INV_X1 U8113 ( .A(n7677), .ZN(n10297) );
  AOI22_X1 U8114 ( .A1(ram[3090]), .A2(n7675), .B1(n10311), .B2(n8907), .ZN(
        n7677) );
  INV_X1 U8115 ( .A(n7678), .ZN(n10298) );
  AOI22_X1 U8116 ( .A1(ram[3091]), .A2(n7675), .B1(n10311), .B2(n8931), .ZN(
        n7678) );
  INV_X1 U8117 ( .A(n7679), .ZN(n10299) );
  AOI22_X1 U8118 ( .A1(ram[3092]), .A2(n7675), .B1(n10311), .B2(n8955), .ZN(
        n7679) );
  INV_X1 U8119 ( .A(n7680), .ZN(n10300) );
  AOI22_X1 U8120 ( .A1(ram[3093]), .A2(n7675), .B1(n10311), .B2(n8979), .ZN(
        n7680) );
  INV_X1 U8121 ( .A(n7681), .ZN(n10301) );
  AOI22_X1 U8122 ( .A1(ram[3094]), .A2(n7675), .B1(n10311), .B2(n9003), .ZN(
        n7681) );
  INV_X1 U8123 ( .A(n7682), .ZN(n10302) );
  AOI22_X1 U8124 ( .A1(ram[3095]), .A2(n7675), .B1(n10311), .B2(n9027), .ZN(
        n7682) );
  INV_X1 U8125 ( .A(n7683), .ZN(n10303) );
  AOI22_X1 U8126 ( .A1(ram[3096]), .A2(n7675), .B1(n10311), .B2(n9051), .ZN(
        n7683) );
  INV_X1 U8127 ( .A(n7684), .ZN(n10304) );
  AOI22_X1 U8128 ( .A1(ram[3097]), .A2(n7675), .B1(n10311), .B2(n9075), .ZN(
        n7684) );
  INV_X1 U8129 ( .A(n7685), .ZN(n10305) );
  AOI22_X1 U8130 ( .A1(ram[3098]), .A2(n7675), .B1(n10311), .B2(n9099), .ZN(
        n7685) );
  INV_X1 U8131 ( .A(n7686), .ZN(n10306) );
  AOI22_X1 U8132 ( .A1(ram[3099]), .A2(n7675), .B1(n10311), .B2(n9123), .ZN(
        n7686) );
  INV_X1 U8133 ( .A(n7687), .ZN(n10307) );
  AOI22_X1 U8134 ( .A1(ram[3100]), .A2(n7675), .B1(n10311), .B2(n9147), .ZN(
        n7687) );
  INV_X1 U8135 ( .A(n7688), .ZN(n10308) );
  AOI22_X1 U8136 ( .A1(ram[3101]), .A2(n7675), .B1(n10311), .B2(n9171), .ZN(
        n7688) );
  INV_X1 U8137 ( .A(n7689), .ZN(n10309) );
  AOI22_X1 U8138 ( .A1(ram[3102]), .A2(n7675), .B1(n10311), .B2(n9195), .ZN(
        n7689) );
  INV_X1 U8139 ( .A(n7690), .ZN(n10310) );
  AOI22_X1 U8140 ( .A1(ram[3103]), .A2(n7675), .B1(n10311), .B2(n9219), .ZN(
        n7690) );
  INV_X1 U8141 ( .A(n7708), .ZN(n10261) );
  AOI22_X1 U8142 ( .A1(ram[3120]), .A2(n7709), .B1(n10277), .B2(n8859), .ZN(
        n7708) );
  INV_X1 U8143 ( .A(n7710), .ZN(n10262) );
  AOI22_X1 U8144 ( .A1(ram[3121]), .A2(n7709), .B1(n10277), .B2(n8883), .ZN(
        n7710) );
  INV_X1 U8145 ( .A(n7711), .ZN(n10263) );
  AOI22_X1 U8146 ( .A1(ram[3122]), .A2(n7709), .B1(n10277), .B2(n8907), .ZN(
        n7711) );
  INV_X1 U8147 ( .A(n7712), .ZN(n10264) );
  AOI22_X1 U8148 ( .A1(ram[3123]), .A2(n7709), .B1(n10277), .B2(n8931), .ZN(
        n7712) );
  INV_X1 U8149 ( .A(n7713), .ZN(n10265) );
  AOI22_X1 U8150 ( .A1(ram[3124]), .A2(n7709), .B1(n10277), .B2(n8955), .ZN(
        n7713) );
  INV_X1 U8151 ( .A(n7714), .ZN(n10266) );
  AOI22_X1 U8152 ( .A1(ram[3125]), .A2(n7709), .B1(n10277), .B2(n8979), .ZN(
        n7714) );
  INV_X1 U8153 ( .A(n7715), .ZN(n10267) );
  AOI22_X1 U8154 ( .A1(ram[3126]), .A2(n7709), .B1(n10277), .B2(n9003), .ZN(
        n7715) );
  INV_X1 U8155 ( .A(n7716), .ZN(n10268) );
  AOI22_X1 U8156 ( .A1(ram[3127]), .A2(n7709), .B1(n10277), .B2(n9027), .ZN(
        n7716) );
  INV_X1 U8157 ( .A(n7717), .ZN(n10269) );
  AOI22_X1 U8158 ( .A1(ram[3128]), .A2(n7709), .B1(n10277), .B2(n9051), .ZN(
        n7717) );
  INV_X1 U8159 ( .A(n7718), .ZN(n10270) );
  AOI22_X1 U8160 ( .A1(ram[3129]), .A2(n7709), .B1(n10277), .B2(n9075), .ZN(
        n7718) );
  INV_X1 U8161 ( .A(n7719), .ZN(n10271) );
  AOI22_X1 U8162 ( .A1(ram[3130]), .A2(n7709), .B1(n10277), .B2(n9099), .ZN(
        n7719) );
  INV_X1 U8163 ( .A(n7720), .ZN(n10272) );
  AOI22_X1 U8164 ( .A1(ram[3131]), .A2(n7709), .B1(n10277), .B2(n9123), .ZN(
        n7720) );
  INV_X1 U8165 ( .A(n7721), .ZN(n10273) );
  AOI22_X1 U8166 ( .A1(ram[3132]), .A2(n7709), .B1(n10277), .B2(n9147), .ZN(
        n7721) );
  INV_X1 U8167 ( .A(n7722), .ZN(n10274) );
  AOI22_X1 U8168 ( .A1(ram[3133]), .A2(n7709), .B1(n10277), .B2(n9171), .ZN(
        n7722) );
  INV_X1 U8169 ( .A(n7723), .ZN(n10275) );
  AOI22_X1 U8170 ( .A1(ram[3134]), .A2(n7709), .B1(n10277), .B2(n9195), .ZN(
        n7723) );
  INV_X1 U8171 ( .A(n7724), .ZN(n10276) );
  AOI22_X1 U8172 ( .A1(ram[3135]), .A2(n7709), .B1(n10277), .B2(n9219), .ZN(
        n7724) );
  INV_X1 U8173 ( .A(n7742), .ZN(n10227) );
  AOI22_X1 U8174 ( .A1(ram[3152]), .A2(n7743), .B1(n10243), .B2(n8858), .ZN(
        n7742) );
  INV_X1 U8175 ( .A(n7744), .ZN(n10228) );
  AOI22_X1 U8176 ( .A1(ram[3153]), .A2(n7743), .B1(n10243), .B2(n8882), .ZN(
        n7744) );
  INV_X1 U8177 ( .A(n7745), .ZN(n10229) );
  AOI22_X1 U8178 ( .A1(ram[3154]), .A2(n7743), .B1(n10243), .B2(n8906), .ZN(
        n7745) );
  INV_X1 U8179 ( .A(n7746), .ZN(n10230) );
  AOI22_X1 U8180 ( .A1(ram[3155]), .A2(n7743), .B1(n10243), .B2(n8930), .ZN(
        n7746) );
  INV_X1 U8181 ( .A(n7747), .ZN(n10231) );
  AOI22_X1 U8182 ( .A1(ram[3156]), .A2(n7743), .B1(n10243), .B2(n8954), .ZN(
        n7747) );
  INV_X1 U8183 ( .A(n7748), .ZN(n10232) );
  AOI22_X1 U8184 ( .A1(ram[3157]), .A2(n7743), .B1(n10243), .B2(n8978), .ZN(
        n7748) );
  INV_X1 U8185 ( .A(n7749), .ZN(n10233) );
  AOI22_X1 U8186 ( .A1(ram[3158]), .A2(n7743), .B1(n10243), .B2(n9002), .ZN(
        n7749) );
  INV_X1 U8187 ( .A(n7750), .ZN(n10234) );
  AOI22_X1 U8188 ( .A1(ram[3159]), .A2(n7743), .B1(n10243), .B2(n9026), .ZN(
        n7750) );
  INV_X1 U8189 ( .A(n7751), .ZN(n10235) );
  AOI22_X1 U8190 ( .A1(ram[3160]), .A2(n7743), .B1(n10243), .B2(n9050), .ZN(
        n7751) );
  INV_X1 U8191 ( .A(n7752), .ZN(n10236) );
  AOI22_X1 U8192 ( .A1(ram[3161]), .A2(n7743), .B1(n10243), .B2(n9074), .ZN(
        n7752) );
  INV_X1 U8193 ( .A(n7753), .ZN(n10237) );
  AOI22_X1 U8194 ( .A1(ram[3162]), .A2(n7743), .B1(n10243), .B2(n9098), .ZN(
        n7753) );
  INV_X1 U8195 ( .A(n7754), .ZN(n10238) );
  AOI22_X1 U8196 ( .A1(ram[3163]), .A2(n7743), .B1(n10243), .B2(n9122), .ZN(
        n7754) );
  INV_X1 U8197 ( .A(n7755), .ZN(n10239) );
  AOI22_X1 U8198 ( .A1(ram[3164]), .A2(n7743), .B1(n10243), .B2(n9146), .ZN(
        n7755) );
  INV_X1 U8199 ( .A(n7756), .ZN(n10240) );
  AOI22_X1 U8200 ( .A1(ram[3165]), .A2(n7743), .B1(n10243), .B2(n9170), .ZN(
        n7756) );
  INV_X1 U8201 ( .A(n7757), .ZN(n10241) );
  AOI22_X1 U8202 ( .A1(ram[3166]), .A2(n7743), .B1(n10243), .B2(n9194), .ZN(
        n7757) );
  INV_X1 U8203 ( .A(n7758), .ZN(n10242) );
  AOI22_X1 U8204 ( .A1(ram[3167]), .A2(n7743), .B1(n10243), .B2(n9218), .ZN(
        n7758) );
  INV_X1 U8205 ( .A(n7776), .ZN(n10193) );
  AOI22_X1 U8206 ( .A1(ram[3184]), .A2(n7777), .B1(n10209), .B2(n8858), .ZN(
        n7776) );
  INV_X1 U8207 ( .A(n7778), .ZN(n10194) );
  AOI22_X1 U8208 ( .A1(ram[3185]), .A2(n7777), .B1(n10209), .B2(n8882), .ZN(
        n7778) );
  INV_X1 U8209 ( .A(n7779), .ZN(n10195) );
  AOI22_X1 U8210 ( .A1(ram[3186]), .A2(n7777), .B1(n10209), .B2(n8906), .ZN(
        n7779) );
  INV_X1 U8211 ( .A(n7780), .ZN(n10196) );
  AOI22_X1 U8212 ( .A1(ram[3187]), .A2(n7777), .B1(n10209), .B2(n8930), .ZN(
        n7780) );
  INV_X1 U8213 ( .A(n7781), .ZN(n10197) );
  AOI22_X1 U8214 ( .A1(ram[3188]), .A2(n7777), .B1(n10209), .B2(n8954), .ZN(
        n7781) );
  INV_X1 U8215 ( .A(n7782), .ZN(n10198) );
  AOI22_X1 U8216 ( .A1(ram[3189]), .A2(n7777), .B1(n10209), .B2(n8978), .ZN(
        n7782) );
  INV_X1 U8217 ( .A(n7783), .ZN(n10199) );
  AOI22_X1 U8218 ( .A1(ram[3190]), .A2(n7777), .B1(n10209), .B2(n9002), .ZN(
        n7783) );
  INV_X1 U8219 ( .A(n7784), .ZN(n10200) );
  AOI22_X1 U8220 ( .A1(ram[3191]), .A2(n7777), .B1(n10209), .B2(n9026), .ZN(
        n7784) );
  INV_X1 U8221 ( .A(n7785), .ZN(n10201) );
  AOI22_X1 U8222 ( .A1(ram[3192]), .A2(n7777), .B1(n10209), .B2(n9050), .ZN(
        n7785) );
  INV_X1 U8223 ( .A(n7786), .ZN(n10202) );
  AOI22_X1 U8224 ( .A1(ram[3193]), .A2(n7777), .B1(n10209), .B2(n9074), .ZN(
        n7786) );
  INV_X1 U8225 ( .A(n7787), .ZN(n10203) );
  AOI22_X1 U8226 ( .A1(ram[3194]), .A2(n7777), .B1(n10209), .B2(n9098), .ZN(
        n7787) );
  INV_X1 U8227 ( .A(n7788), .ZN(n10204) );
  AOI22_X1 U8228 ( .A1(ram[3195]), .A2(n7777), .B1(n10209), .B2(n9122), .ZN(
        n7788) );
  INV_X1 U8229 ( .A(n7789), .ZN(n10205) );
  AOI22_X1 U8230 ( .A1(ram[3196]), .A2(n7777), .B1(n10209), .B2(n9146), .ZN(
        n7789) );
  INV_X1 U8231 ( .A(n7790), .ZN(n10206) );
  AOI22_X1 U8232 ( .A1(ram[3197]), .A2(n7777), .B1(n10209), .B2(n9170), .ZN(
        n7790) );
  INV_X1 U8233 ( .A(n7791), .ZN(n10207) );
  AOI22_X1 U8234 ( .A1(ram[3198]), .A2(n7777), .B1(n10209), .B2(n9194), .ZN(
        n7791) );
  INV_X1 U8235 ( .A(n7792), .ZN(n10208) );
  AOI22_X1 U8236 ( .A1(ram[3199]), .A2(n7777), .B1(n10209), .B2(n9218), .ZN(
        n7792) );
  INV_X1 U8237 ( .A(n7810), .ZN(n10159) );
  AOI22_X1 U8238 ( .A1(ram[3216]), .A2(n7811), .B1(n10175), .B2(n8858), .ZN(
        n7810) );
  INV_X1 U8239 ( .A(n7812), .ZN(n10160) );
  AOI22_X1 U8240 ( .A1(ram[3217]), .A2(n7811), .B1(n10175), .B2(n8882), .ZN(
        n7812) );
  INV_X1 U8241 ( .A(n7813), .ZN(n10161) );
  AOI22_X1 U8242 ( .A1(ram[3218]), .A2(n7811), .B1(n10175), .B2(n8906), .ZN(
        n7813) );
  INV_X1 U8243 ( .A(n7814), .ZN(n10162) );
  AOI22_X1 U8244 ( .A1(ram[3219]), .A2(n7811), .B1(n10175), .B2(n8930), .ZN(
        n7814) );
  INV_X1 U8245 ( .A(n7815), .ZN(n10163) );
  AOI22_X1 U8246 ( .A1(ram[3220]), .A2(n7811), .B1(n10175), .B2(n8954), .ZN(
        n7815) );
  INV_X1 U8247 ( .A(n7816), .ZN(n10164) );
  AOI22_X1 U8248 ( .A1(ram[3221]), .A2(n7811), .B1(n10175), .B2(n8978), .ZN(
        n7816) );
  INV_X1 U8249 ( .A(n7817), .ZN(n10165) );
  AOI22_X1 U8250 ( .A1(ram[3222]), .A2(n7811), .B1(n10175), .B2(n9002), .ZN(
        n7817) );
  INV_X1 U8251 ( .A(n7818), .ZN(n10166) );
  AOI22_X1 U8252 ( .A1(ram[3223]), .A2(n7811), .B1(n10175), .B2(n9026), .ZN(
        n7818) );
  INV_X1 U8253 ( .A(n7819), .ZN(n10167) );
  AOI22_X1 U8254 ( .A1(ram[3224]), .A2(n7811), .B1(n10175), .B2(n9050), .ZN(
        n7819) );
  INV_X1 U8255 ( .A(n7820), .ZN(n10168) );
  AOI22_X1 U8256 ( .A1(ram[3225]), .A2(n7811), .B1(n10175), .B2(n9074), .ZN(
        n7820) );
  INV_X1 U8257 ( .A(n7821), .ZN(n10169) );
  AOI22_X1 U8258 ( .A1(ram[3226]), .A2(n7811), .B1(n10175), .B2(n9098), .ZN(
        n7821) );
  INV_X1 U8259 ( .A(n7822), .ZN(n10170) );
  AOI22_X1 U8260 ( .A1(ram[3227]), .A2(n7811), .B1(n10175), .B2(n9122), .ZN(
        n7822) );
  INV_X1 U8261 ( .A(n7823), .ZN(n10171) );
  AOI22_X1 U8262 ( .A1(ram[3228]), .A2(n7811), .B1(n10175), .B2(n9146), .ZN(
        n7823) );
  INV_X1 U8263 ( .A(n7824), .ZN(n10172) );
  AOI22_X1 U8264 ( .A1(ram[3229]), .A2(n7811), .B1(n10175), .B2(n9170), .ZN(
        n7824) );
  INV_X1 U8265 ( .A(n7825), .ZN(n10173) );
  AOI22_X1 U8266 ( .A1(ram[3230]), .A2(n7811), .B1(n10175), .B2(n9194), .ZN(
        n7825) );
  INV_X1 U8267 ( .A(n7826), .ZN(n10174) );
  AOI22_X1 U8268 ( .A1(ram[3231]), .A2(n7811), .B1(n10175), .B2(n9218), .ZN(
        n7826) );
  INV_X1 U8269 ( .A(n7844), .ZN(n10125) );
  AOI22_X1 U8270 ( .A1(ram[3248]), .A2(n7845), .B1(n10141), .B2(n8858), .ZN(
        n7844) );
  INV_X1 U8271 ( .A(n7846), .ZN(n10126) );
  AOI22_X1 U8272 ( .A1(ram[3249]), .A2(n7845), .B1(n10141), .B2(n8882), .ZN(
        n7846) );
  INV_X1 U8273 ( .A(n7847), .ZN(n10127) );
  AOI22_X1 U8274 ( .A1(ram[3250]), .A2(n7845), .B1(n10141), .B2(n8906), .ZN(
        n7847) );
  INV_X1 U8275 ( .A(n7848), .ZN(n10128) );
  AOI22_X1 U8276 ( .A1(ram[3251]), .A2(n7845), .B1(n10141), .B2(n8930), .ZN(
        n7848) );
  INV_X1 U8277 ( .A(n7849), .ZN(n10129) );
  AOI22_X1 U8278 ( .A1(ram[3252]), .A2(n7845), .B1(n10141), .B2(n8954), .ZN(
        n7849) );
  INV_X1 U8279 ( .A(n7850), .ZN(n10130) );
  AOI22_X1 U8280 ( .A1(ram[3253]), .A2(n7845), .B1(n10141), .B2(n8978), .ZN(
        n7850) );
  INV_X1 U8281 ( .A(n7851), .ZN(n10131) );
  AOI22_X1 U8282 ( .A1(ram[3254]), .A2(n7845), .B1(n10141), .B2(n9002), .ZN(
        n7851) );
  INV_X1 U8283 ( .A(n7852), .ZN(n10132) );
  AOI22_X1 U8284 ( .A1(ram[3255]), .A2(n7845), .B1(n10141), .B2(n9026), .ZN(
        n7852) );
  INV_X1 U8285 ( .A(n7853), .ZN(n10133) );
  AOI22_X1 U8286 ( .A1(ram[3256]), .A2(n7845), .B1(n10141), .B2(n9050), .ZN(
        n7853) );
  INV_X1 U8287 ( .A(n7854), .ZN(n10134) );
  AOI22_X1 U8288 ( .A1(ram[3257]), .A2(n7845), .B1(n10141), .B2(n9074), .ZN(
        n7854) );
  INV_X1 U8289 ( .A(n7855), .ZN(n10135) );
  AOI22_X1 U8290 ( .A1(ram[3258]), .A2(n7845), .B1(n10141), .B2(n9098), .ZN(
        n7855) );
  INV_X1 U8291 ( .A(n7856), .ZN(n10136) );
  AOI22_X1 U8292 ( .A1(ram[3259]), .A2(n7845), .B1(n10141), .B2(n9122), .ZN(
        n7856) );
  INV_X1 U8293 ( .A(n7857), .ZN(n10137) );
  AOI22_X1 U8294 ( .A1(ram[3260]), .A2(n7845), .B1(n10141), .B2(n9146), .ZN(
        n7857) );
  INV_X1 U8295 ( .A(n7858), .ZN(n10138) );
  AOI22_X1 U8296 ( .A1(ram[3261]), .A2(n7845), .B1(n10141), .B2(n9170), .ZN(
        n7858) );
  INV_X1 U8297 ( .A(n7859), .ZN(n10139) );
  AOI22_X1 U8298 ( .A1(ram[3262]), .A2(n7845), .B1(n10141), .B2(n9194), .ZN(
        n7859) );
  INV_X1 U8299 ( .A(n7860), .ZN(n10140) );
  AOI22_X1 U8300 ( .A1(ram[3263]), .A2(n7845), .B1(n10141), .B2(n9218), .ZN(
        n7860) );
  INV_X1 U8301 ( .A(n7878), .ZN(n10091) );
  AOI22_X1 U8302 ( .A1(ram[3280]), .A2(n7879), .B1(n10107), .B2(n8858), .ZN(
        n7878) );
  INV_X1 U8303 ( .A(n7880), .ZN(n10092) );
  AOI22_X1 U8304 ( .A1(ram[3281]), .A2(n7879), .B1(n10107), .B2(n8882), .ZN(
        n7880) );
  INV_X1 U8305 ( .A(n7881), .ZN(n10093) );
  AOI22_X1 U8306 ( .A1(ram[3282]), .A2(n7879), .B1(n10107), .B2(n8906), .ZN(
        n7881) );
  INV_X1 U8307 ( .A(n7882), .ZN(n10094) );
  AOI22_X1 U8308 ( .A1(ram[3283]), .A2(n7879), .B1(n10107), .B2(n8930), .ZN(
        n7882) );
  INV_X1 U8309 ( .A(n7883), .ZN(n10095) );
  AOI22_X1 U8310 ( .A1(ram[3284]), .A2(n7879), .B1(n10107), .B2(n8954), .ZN(
        n7883) );
  INV_X1 U8311 ( .A(n7884), .ZN(n10096) );
  AOI22_X1 U8312 ( .A1(ram[3285]), .A2(n7879), .B1(n10107), .B2(n8978), .ZN(
        n7884) );
  INV_X1 U8313 ( .A(n7885), .ZN(n10097) );
  AOI22_X1 U8314 ( .A1(ram[3286]), .A2(n7879), .B1(n10107), .B2(n9002), .ZN(
        n7885) );
  INV_X1 U8315 ( .A(n7886), .ZN(n10098) );
  AOI22_X1 U8316 ( .A1(ram[3287]), .A2(n7879), .B1(n10107), .B2(n9026), .ZN(
        n7886) );
  INV_X1 U8317 ( .A(n7887), .ZN(n10099) );
  AOI22_X1 U8318 ( .A1(ram[3288]), .A2(n7879), .B1(n10107), .B2(n9050), .ZN(
        n7887) );
  INV_X1 U8319 ( .A(n7888), .ZN(n10100) );
  AOI22_X1 U8320 ( .A1(ram[3289]), .A2(n7879), .B1(n10107), .B2(n9074), .ZN(
        n7888) );
  INV_X1 U8321 ( .A(n7889), .ZN(n10101) );
  AOI22_X1 U8322 ( .A1(ram[3290]), .A2(n7879), .B1(n10107), .B2(n9098), .ZN(
        n7889) );
  INV_X1 U8323 ( .A(n7890), .ZN(n10102) );
  AOI22_X1 U8324 ( .A1(ram[3291]), .A2(n7879), .B1(n10107), .B2(n9122), .ZN(
        n7890) );
  INV_X1 U8325 ( .A(n7891), .ZN(n10103) );
  AOI22_X1 U8326 ( .A1(ram[3292]), .A2(n7879), .B1(n10107), .B2(n9146), .ZN(
        n7891) );
  INV_X1 U8327 ( .A(n7892), .ZN(n10104) );
  AOI22_X1 U8328 ( .A1(ram[3293]), .A2(n7879), .B1(n10107), .B2(n9170), .ZN(
        n7892) );
  INV_X1 U8329 ( .A(n7893), .ZN(n10105) );
  AOI22_X1 U8330 ( .A1(ram[3294]), .A2(n7879), .B1(n10107), .B2(n9194), .ZN(
        n7893) );
  INV_X1 U8331 ( .A(n7894), .ZN(n10106) );
  AOI22_X1 U8332 ( .A1(ram[3295]), .A2(n7879), .B1(n10107), .B2(n9218), .ZN(
        n7894) );
  INV_X1 U8333 ( .A(n7912), .ZN(n10057) );
  AOI22_X1 U8334 ( .A1(ram[3312]), .A2(n7913), .B1(n10073), .B2(n8858), .ZN(
        n7912) );
  INV_X1 U8335 ( .A(n7914), .ZN(n10058) );
  AOI22_X1 U8336 ( .A1(ram[3313]), .A2(n7913), .B1(n10073), .B2(n8882), .ZN(
        n7914) );
  INV_X1 U8337 ( .A(n7915), .ZN(n10059) );
  AOI22_X1 U8338 ( .A1(ram[3314]), .A2(n7913), .B1(n10073), .B2(n8906), .ZN(
        n7915) );
  INV_X1 U8339 ( .A(n7916), .ZN(n10060) );
  AOI22_X1 U8340 ( .A1(ram[3315]), .A2(n7913), .B1(n10073), .B2(n8930), .ZN(
        n7916) );
  INV_X1 U8341 ( .A(n7917), .ZN(n10061) );
  AOI22_X1 U8342 ( .A1(ram[3316]), .A2(n7913), .B1(n10073), .B2(n8954), .ZN(
        n7917) );
  INV_X1 U8343 ( .A(n7918), .ZN(n10062) );
  AOI22_X1 U8344 ( .A1(ram[3317]), .A2(n7913), .B1(n10073), .B2(n8978), .ZN(
        n7918) );
  INV_X1 U8345 ( .A(n7919), .ZN(n10063) );
  AOI22_X1 U8346 ( .A1(ram[3318]), .A2(n7913), .B1(n10073), .B2(n9002), .ZN(
        n7919) );
  INV_X1 U8347 ( .A(n7920), .ZN(n10064) );
  AOI22_X1 U8348 ( .A1(ram[3319]), .A2(n7913), .B1(n10073), .B2(n9026), .ZN(
        n7920) );
  INV_X1 U8349 ( .A(n7921), .ZN(n10065) );
  AOI22_X1 U8350 ( .A1(ram[3320]), .A2(n7913), .B1(n10073), .B2(n9050), .ZN(
        n7921) );
  INV_X1 U8351 ( .A(n7922), .ZN(n10066) );
  AOI22_X1 U8352 ( .A1(ram[3321]), .A2(n7913), .B1(n10073), .B2(n9074), .ZN(
        n7922) );
  INV_X1 U8353 ( .A(n7923), .ZN(n10067) );
  AOI22_X1 U8354 ( .A1(ram[3322]), .A2(n7913), .B1(n10073), .B2(n9098), .ZN(
        n7923) );
  INV_X1 U8355 ( .A(n7924), .ZN(n10068) );
  AOI22_X1 U8356 ( .A1(ram[3323]), .A2(n7913), .B1(n10073), .B2(n9122), .ZN(
        n7924) );
  INV_X1 U8357 ( .A(n7925), .ZN(n10069) );
  AOI22_X1 U8358 ( .A1(ram[3324]), .A2(n7913), .B1(n10073), .B2(n9146), .ZN(
        n7925) );
  INV_X1 U8359 ( .A(n7926), .ZN(n10070) );
  AOI22_X1 U8360 ( .A1(ram[3325]), .A2(n7913), .B1(n10073), .B2(n9170), .ZN(
        n7926) );
  INV_X1 U8361 ( .A(n7927), .ZN(n10071) );
  AOI22_X1 U8362 ( .A1(ram[3326]), .A2(n7913), .B1(n10073), .B2(n9194), .ZN(
        n7927) );
  INV_X1 U8363 ( .A(n7928), .ZN(n10072) );
  AOI22_X1 U8364 ( .A1(ram[3327]), .A2(n7913), .B1(n10073), .B2(n9218), .ZN(
        n7928) );
  INV_X1 U8365 ( .A(n7948), .ZN(n10023) );
  AOI22_X1 U8366 ( .A1(ram[3344]), .A2(n7949), .B1(n10039), .B2(n8857), .ZN(
        n7948) );
  INV_X1 U8367 ( .A(n7950), .ZN(n10024) );
  AOI22_X1 U8368 ( .A1(ram[3345]), .A2(n7949), .B1(n10039), .B2(n8881), .ZN(
        n7950) );
  INV_X1 U8369 ( .A(n7951), .ZN(n10025) );
  AOI22_X1 U8370 ( .A1(ram[3346]), .A2(n7949), .B1(n10039), .B2(n8905), .ZN(
        n7951) );
  INV_X1 U8371 ( .A(n7952), .ZN(n10026) );
  AOI22_X1 U8372 ( .A1(ram[3347]), .A2(n7949), .B1(n10039), .B2(n8929), .ZN(
        n7952) );
  INV_X1 U8373 ( .A(n7953), .ZN(n10027) );
  AOI22_X1 U8374 ( .A1(ram[3348]), .A2(n7949), .B1(n10039), .B2(n8953), .ZN(
        n7953) );
  INV_X1 U8375 ( .A(n7954), .ZN(n10028) );
  AOI22_X1 U8376 ( .A1(ram[3349]), .A2(n7949), .B1(n10039), .B2(n8977), .ZN(
        n7954) );
  INV_X1 U8377 ( .A(n7955), .ZN(n10029) );
  AOI22_X1 U8378 ( .A1(ram[3350]), .A2(n7949), .B1(n10039), .B2(n9001), .ZN(
        n7955) );
  INV_X1 U8379 ( .A(n7956), .ZN(n10030) );
  AOI22_X1 U8380 ( .A1(ram[3351]), .A2(n7949), .B1(n10039), .B2(n9025), .ZN(
        n7956) );
  INV_X1 U8381 ( .A(n7957), .ZN(n10031) );
  AOI22_X1 U8382 ( .A1(ram[3352]), .A2(n7949), .B1(n10039), .B2(n9049), .ZN(
        n7957) );
  INV_X1 U8383 ( .A(n7958), .ZN(n10032) );
  AOI22_X1 U8384 ( .A1(ram[3353]), .A2(n7949), .B1(n10039), .B2(n9073), .ZN(
        n7958) );
  INV_X1 U8385 ( .A(n7959), .ZN(n10033) );
  AOI22_X1 U8386 ( .A1(ram[3354]), .A2(n7949), .B1(n10039), .B2(n9097), .ZN(
        n7959) );
  INV_X1 U8387 ( .A(n7960), .ZN(n10034) );
  AOI22_X1 U8388 ( .A1(ram[3355]), .A2(n7949), .B1(n10039), .B2(n9121), .ZN(
        n7960) );
  INV_X1 U8389 ( .A(n7961), .ZN(n10035) );
  AOI22_X1 U8390 ( .A1(ram[3356]), .A2(n7949), .B1(n10039), .B2(n9145), .ZN(
        n7961) );
  INV_X1 U8391 ( .A(n7962), .ZN(n10036) );
  AOI22_X1 U8392 ( .A1(ram[3357]), .A2(n7949), .B1(n10039), .B2(n9169), .ZN(
        n7962) );
  INV_X1 U8393 ( .A(n7963), .ZN(n10037) );
  AOI22_X1 U8394 ( .A1(ram[3358]), .A2(n7949), .B1(n10039), .B2(n9193), .ZN(
        n7963) );
  INV_X1 U8395 ( .A(n7964), .ZN(n10038) );
  AOI22_X1 U8396 ( .A1(ram[3359]), .A2(n7949), .B1(n10039), .B2(n9217), .ZN(
        n7964) );
  INV_X1 U8397 ( .A(n7982), .ZN(n9989) );
  AOI22_X1 U8398 ( .A1(ram[3376]), .A2(n7983), .B1(n10005), .B2(n8857), .ZN(
        n7982) );
  INV_X1 U8399 ( .A(n7984), .ZN(n9990) );
  AOI22_X1 U8400 ( .A1(ram[3377]), .A2(n7983), .B1(n10005), .B2(n8881), .ZN(
        n7984) );
  INV_X1 U8401 ( .A(n7985), .ZN(n9991) );
  AOI22_X1 U8402 ( .A1(ram[3378]), .A2(n7983), .B1(n10005), .B2(n8905), .ZN(
        n7985) );
  INV_X1 U8403 ( .A(n7986), .ZN(n9992) );
  AOI22_X1 U8404 ( .A1(ram[3379]), .A2(n7983), .B1(n10005), .B2(n8929), .ZN(
        n7986) );
  INV_X1 U8405 ( .A(n7987), .ZN(n9993) );
  AOI22_X1 U8406 ( .A1(ram[3380]), .A2(n7983), .B1(n10005), .B2(n8953), .ZN(
        n7987) );
  INV_X1 U8407 ( .A(n7988), .ZN(n9994) );
  AOI22_X1 U8408 ( .A1(ram[3381]), .A2(n7983), .B1(n10005), .B2(n8977), .ZN(
        n7988) );
  INV_X1 U8409 ( .A(n7989), .ZN(n9995) );
  AOI22_X1 U8410 ( .A1(ram[3382]), .A2(n7983), .B1(n10005), .B2(n9001), .ZN(
        n7989) );
  INV_X1 U8411 ( .A(n7990), .ZN(n9996) );
  AOI22_X1 U8412 ( .A1(ram[3383]), .A2(n7983), .B1(n10005), .B2(n9025), .ZN(
        n7990) );
  INV_X1 U8413 ( .A(n7991), .ZN(n9997) );
  AOI22_X1 U8414 ( .A1(ram[3384]), .A2(n7983), .B1(n10005), .B2(n9049), .ZN(
        n7991) );
  INV_X1 U8415 ( .A(n7992), .ZN(n9998) );
  AOI22_X1 U8416 ( .A1(ram[3385]), .A2(n7983), .B1(n10005), .B2(n9073), .ZN(
        n7992) );
  INV_X1 U8417 ( .A(n7993), .ZN(n9999) );
  AOI22_X1 U8418 ( .A1(ram[3386]), .A2(n7983), .B1(n10005), .B2(n9097), .ZN(
        n7993) );
  INV_X1 U8419 ( .A(n7994), .ZN(n10000) );
  AOI22_X1 U8420 ( .A1(ram[3387]), .A2(n7983), .B1(n10005), .B2(n9121), .ZN(
        n7994) );
  INV_X1 U8421 ( .A(n7995), .ZN(n10001) );
  AOI22_X1 U8422 ( .A1(ram[3388]), .A2(n7983), .B1(n10005), .B2(n9145), .ZN(
        n7995) );
  INV_X1 U8423 ( .A(n7996), .ZN(n10002) );
  AOI22_X1 U8424 ( .A1(ram[3389]), .A2(n7983), .B1(n10005), .B2(n9169), .ZN(
        n7996) );
  INV_X1 U8425 ( .A(n7997), .ZN(n10003) );
  AOI22_X1 U8426 ( .A1(ram[3390]), .A2(n7983), .B1(n10005), .B2(n9193), .ZN(
        n7997) );
  INV_X1 U8427 ( .A(n7998), .ZN(n10004) );
  AOI22_X1 U8428 ( .A1(ram[3391]), .A2(n7983), .B1(n10005), .B2(n9217), .ZN(
        n7998) );
  INV_X1 U8429 ( .A(n8016), .ZN(n9955) );
  AOI22_X1 U8430 ( .A1(ram[3408]), .A2(n8017), .B1(n9971), .B2(n8857), .ZN(
        n8016) );
  INV_X1 U8431 ( .A(n8018), .ZN(n9956) );
  AOI22_X1 U8432 ( .A1(ram[3409]), .A2(n8017), .B1(n9971), .B2(n8881), .ZN(
        n8018) );
  INV_X1 U8433 ( .A(n8019), .ZN(n9957) );
  AOI22_X1 U8434 ( .A1(ram[3410]), .A2(n8017), .B1(n9971), .B2(n8905), .ZN(
        n8019) );
  INV_X1 U8435 ( .A(n8020), .ZN(n9958) );
  AOI22_X1 U8436 ( .A1(ram[3411]), .A2(n8017), .B1(n9971), .B2(n8929), .ZN(
        n8020) );
  INV_X1 U8437 ( .A(n8021), .ZN(n9959) );
  AOI22_X1 U8438 ( .A1(ram[3412]), .A2(n8017), .B1(n9971), .B2(n8953), .ZN(
        n8021) );
  INV_X1 U8439 ( .A(n8022), .ZN(n9960) );
  AOI22_X1 U8440 ( .A1(ram[3413]), .A2(n8017), .B1(n9971), .B2(n8977), .ZN(
        n8022) );
  INV_X1 U8441 ( .A(n8023), .ZN(n9961) );
  AOI22_X1 U8442 ( .A1(ram[3414]), .A2(n8017), .B1(n9971), .B2(n9001), .ZN(
        n8023) );
  INV_X1 U8443 ( .A(n8024), .ZN(n9962) );
  AOI22_X1 U8444 ( .A1(ram[3415]), .A2(n8017), .B1(n9971), .B2(n9025), .ZN(
        n8024) );
  INV_X1 U8445 ( .A(n8025), .ZN(n9963) );
  AOI22_X1 U8446 ( .A1(ram[3416]), .A2(n8017), .B1(n9971), .B2(n9049), .ZN(
        n8025) );
  INV_X1 U8447 ( .A(n8026), .ZN(n9964) );
  AOI22_X1 U8448 ( .A1(ram[3417]), .A2(n8017), .B1(n9971), .B2(n9073), .ZN(
        n8026) );
  INV_X1 U8449 ( .A(n8027), .ZN(n9965) );
  AOI22_X1 U8450 ( .A1(ram[3418]), .A2(n8017), .B1(n9971), .B2(n9097), .ZN(
        n8027) );
  INV_X1 U8451 ( .A(n8028), .ZN(n9966) );
  AOI22_X1 U8452 ( .A1(ram[3419]), .A2(n8017), .B1(n9971), .B2(n9121), .ZN(
        n8028) );
  INV_X1 U8453 ( .A(n8029), .ZN(n9967) );
  AOI22_X1 U8454 ( .A1(ram[3420]), .A2(n8017), .B1(n9971), .B2(n9145), .ZN(
        n8029) );
  INV_X1 U8455 ( .A(n8030), .ZN(n9968) );
  AOI22_X1 U8456 ( .A1(ram[3421]), .A2(n8017), .B1(n9971), .B2(n9169), .ZN(
        n8030) );
  INV_X1 U8457 ( .A(n8031), .ZN(n9969) );
  AOI22_X1 U8458 ( .A1(ram[3422]), .A2(n8017), .B1(n9971), .B2(n9193), .ZN(
        n8031) );
  INV_X1 U8459 ( .A(n8032), .ZN(n9970) );
  AOI22_X1 U8460 ( .A1(ram[3423]), .A2(n8017), .B1(n9971), .B2(n9217), .ZN(
        n8032) );
  INV_X1 U8461 ( .A(n8050), .ZN(n9921) );
  AOI22_X1 U8462 ( .A1(ram[3440]), .A2(n8051), .B1(n9937), .B2(n8857), .ZN(
        n8050) );
  INV_X1 U8463 ( .A(n8052), .ZN(n9922) );
  AOI22_X1 U8464 ( .A1(ram[3441]), .A2(n8051), .B1(n9937), .B2(n8881), .ZN(
        n8052) );
  INV_X1 U8465 ( .A(n8053), .ZN(n9923) );
  AOI22_X1 U8466 ( .A1(ram[3442]), .A2(n8051), .B1(n9937), .B2(n8905), .ZN(
        n8053) );
  INV_X1 U8467 ( .A(n8054), .ZN(n9924) );
  AOI22_X1 U8468 ( .A1(ram[3443]), .A2(n8051), .B1(n9937), .B2(n8929), .ZN(
        n8054) );
  INV_X1 U8469 ( .A(n8055), .ZN(n9925) );
  AOI22_X1 U8470 ( .A1(ram[3444]), .A2(n8051), .B1(n9937), .B2(n8953), .ZN(
        n8055) );
  INV_X1 U8471 ( .A(n8056), .ZN(n9926) );
  AOI22_X1 U8472 ( .A1(ram[3445]), .A2(n8051), .B1(n9937), .B2(n8977), .ZN(
        n8056) );
  INV_X1 U8473 ( .A(n8057), .ZN(n9927) );
  AOI22_X1 U8474 ( .A1(ram[3446]), .A2(n8051), .B1(n9937), .B2(n9001), .ZN(
        n8057) );
  INV_X1 U8475 ( .A(n8058), .ZN(n9928) );
  AOI22_X1 U8476 ( .A1(ram[3447]), .A2(n8051), .B1(n9937), .B2(n9025), .ZN(
        n8058) );
  INV_X1 U8477 ( .A(n8059), .ZN(n9929) );
  AOI22_X1 U8478 ( .A1(ram[3448]), .A2(n8051), .B1(n9937), .B2(n9049), .ZN(
        n8059) );
  INV_X1 U8479 ( .A(n8060), .ZN(n9930) );
  AOI22_X1 U8480 ( .A1(ram[3449]), .A2(n8051), .B1(n9937), .B2(n9073), .ZN(
        n8060) );
  INV_X1 U8481 ( .A(n8061), .ZN(n9931) );
  AOI22_X1 U8482 ( .A1(ram[3450]), .A2(n8051), .B1(n9937), .B2(n9097), .ZN(
        n8061) );
  INV_X1 U8483 ( .A(n8062), .ZN(n9932) );
  AOI22_X1 U8484 ( .A1(ram[3451]), .A2(n8051), .B1(n9937), .B2(n9121), .ZN(
        n8062) );
  INV_X1 U8485 ( .A(n8063), .ZN(n9933) );
  AOI22_X1 U8486 ( .A1(ram[3452]), .A2(n8051), .B1(n9937), .B2(n9145), .ZN(
        n8063) );
  INV_X1 U8487 ( .A(n8064), .ZN(n9934) );
  AOI22_X1 U8488 ( .A1(ram[3453]), .A2(n8051), .B1(n9937), .B2(n9169), .ZN(
        n8064) );
  INV_X1 U8489 ( .A(n8065), .ZN(n9935) );
  AOI22_X1 U8490 ( .A1(ram[3454]), .A2(n8051), .B1(n9937), .B2(n9193), .ZN(
        n8065) );
  INV_X1 U8491 ( .A(n8066), .ZN(n9936) );
  AOI22_X1 U8492 ( .A1(ram[3455]), .A2(n8051), .B1(n9937), .B2(n9217), .ZN(
        n8066) );
  INV_X1 U8493 ( .A(n8084), .ZN(n9887) );
  AOI22_X1 U8494 ( .A1(ram[3472]), .A2(n8085), .B1(n9903), .B2(n8857), .ZN(
        n8084) );
  INV_X1 U8495 ( .A(n8086), .ZN(n9888) );
  AOI22_X1 U8496 ( .A1(ram[3473]), .A2(n8085), .B1(n9903), .B2(n8881), .ZN(
        n8086) );
  INV_X1 U8497 ( .A(n8087), .ZN(n9889) );
  AOI22_X1 U8498 ( .A1(ram[3474]), .A2(n8085), .B1(n9903), .B2(n8905), .ZN(
        n8087) );
  INV_X1 U8499 ( .A(n8088), .ZN(n9890) );
  AOI22_X1 U8500 ( .A1(ram[3475]), .A2(n8085), .B1(n9903), .B2(n8929), .ZN(
        n8088) );
  INV_X1 U8501 ( .A(n8089), .ZN(n9891) );
  AOI22_X1 U8502 ( .A1(ram[3476]), .A2(n8085), .B1(n9903), .B2(n8953), .ZN(
        n8089) );
  INV_X1 U8503 ( .A(n8090), .ZN(n9892) );
  AOI22_X1 U8504 ( .A1(ram[3477]), .A2(n8085), .B1(n9903), .B2(n8977), .ZN(
        n8090) );
  INV_X1 U8505 ( .A(n8091), .ZN(n9893) );
  AOI22_X1 U8506 ( .A1(ram[3478]), .A2(n8085), .B1(n9903), .B2(n9001), .ZN(
        n8091) );
  INV_X1 U8507 ( .A(n8092), .ZN(n9894) );
  AOI22_X1 U8508 ( .A1(ram[3479]), .A2(n8085), .B1(n9903), .B2(n9025), .ZN(
        n8092) );
  INV_X1 U8509 ( .A(n8093), .ZN(n9895) );
  AOI22_X1 U8510 ( .A1(ram[3480]), .A2(n8085), .B1(n9903), .B2(n9049), .ZN(
        n8093) );
  INV_X1 U8511 ( .A(n8094), .ZN(n9896) );
  AOI22_X1 U8512 ( .A1(ram[3481]), .A2(n8085), .B1(n9903), .B2(n9073), .ZN(
        n8094) );
  INV_X1 U8513 ( .A(n8095), .ZN(n9897) );
  AOI22_X1 U8514 ( .A1(ram[3482]), .A2(n8085), .B1(n9903), .B2(n9097), .ZN(
        n8095) );
  INV_X1 U8515 ( .A(n8096), .ZN(n9898) );
  AOI22_X1 U8516 ( .A1(ram[3483]), .A2(n8085), .B1(n9903), .B2(n9121), .ZN(
        n8096) );
  INV_X1 U8517 ( .A(n8097), .ZN(n9899) );
  AOI22_X1 U8518 ( .A1(ram[3484]), .A2(n8085), .B1(n9903), .B2(n9145), .ZN(
        n8097) );
  INV_X1 U8519 ( .A(n8098), .ZN(n9900) );
  AOI22_X1 U8520 ( .A1(ram[3485]), .A2(n8085), .B1(n9903), .B2(n9169), .ZN(
        n8098) );
  INV_X1 U8521 ( .A(n8099), .ZN(n9901) );
  AOI22_X1 U8522 ( .A1(ram[3486]), .A2(n8085), .B1(n9903), .B2(n9193), .ZN(
        n8099) );
  INV_X1 U8523 ( .A(n8100), .ZN(n9902) );
  AOI22_X1 U8524 ( .A1(ram[3487]), .A2(n8085), .B1(n9903), .B2(n9217), .ZN(
        n8100) );
  INV_X1 U8525 ( .A(n8118), .ZN(n9853) );
  AOI22_X1 U8526 ( .A1(ram[3504]), .A2(n8119), .B1(n9869), .B2(n8857), .ZN(
        n8118) );
  INV_X1 U8527 ( .A(n8120), .ZN(n9854) );
  AOI22_X1 U8528 ( .A1(ram[3505]), .A2(n8119), .B1(n9869), .B2(n8881), .ZN(
        n8120) );
  INV_X1 U8529 ( .A(n8121), .ZN(n9855) );
  AOI22_X1 U8530 ( .A1(ram[3506]), .A2(n8119), .B1(n9869), .B2(n8905), .ZN(
        n8121) );
  INV_X1 U8531 ( .A(n8122), .ZN(n9856) );
  AOI22_X1 U8532 ( .A1(ram[3507]), .A2(n8119), .B1(n9869), .B2(n8929), .ZN(
        n8122) );
  INV_X1 U8533 ( .A(n8123), .ZN(n9857) );
  AOI22_X1 U8534 ( .A1(ram[3508]), .A2(n8119), .B1(n9869), .B2(n8953), .ZN(
        n8123) );
  INV_X1 U8535 ( .A(n8124), .ZN(n9858) );
  AOI22_X1 U8536 ( .A1(ram[3509]), .A2(n8119), .B1(n9869), .B2(n8977), .ZN(
        n8124) );
  INV_X1 U8537 ( .A(n8125), .ZN(n9859) );
  AOI22_X1 U8538 ( .A1(ram[3510]), .A2(n8119), .B1(n9869), .B2(n9001), .ZN(
        n8125) );
  INV_X1 U8539 ( .A(n8126), .ZN(n9860) );
  AOI22_X1 U8540 ( .A1(ram[3511]), .A2(n8119), .B1(n9869), .B2(n9025), .ZN(
        n8126) );
  INV_X1 U8541 ( .A(n8127), .ZN(n9861) );
  AOI22_X1 U8542 ( .A1(ram[3512]), .A2(n8119), .B1(n9869), .B2(n9049), .ZN(
        n8127) );
  INV_X1 U8543 ( .A(n8128), .ZN(n9862) );
  AOI22_X1 U8544 ( .A1(ram[3513]), .A2(n8119), .B1(n9869), .B2(n9073), .ZN(
        n8128) );
  INV_X1 U8545 ( .A(n8129), .ZN(n9863) );
  AOI22_X1 U8546 ( .A1(ram[3514]), .A2(n8119), .B1(n9869), .B2(n9097), .ZN(
        n8129) );
  INV_X1 U8547 ( .A(n8130), .ZN(n9864) );
  AOI22_X1 U8548 ( .A1(ram[3515]), .A2(n8119), .B1(n9869), .B2(n9121), .ZN(
        n8130) );
  INV_X1 U8549 ( .A(n8131), .ZN(n9865) );
  AOI22_X1 U8550 ( .A1(ram[3516]), .A2(n8119), .B1(n9869), .B2(n9145), .ZN(
        n8131) );
  INV_X1 U8551 ( .A(n8132), .ZN(n9866) );
  AOI22_X1 U8552 ( .A1(ram[3517]), .A2(n8119), .B1(n9869), .B2(n9169), .ZN(
        n8132) );
  INV_X1 U8553 ( .A(n8133), .ZN(n9867) );
  AOI22_X1 U8554 ( .A1(ram[3518]), .A2(n8119), .B1(n9869), .B2(n9193), .ZN(
        n8133) );
  INV_X1 U8555 ( .A(n8134), .ZN(n9868) );
  AOI22_X1 U8556 ( .A1(ram[3519]), .A2(n8119), .B1(n9869), .B2(n9217), .ZN(
        n8134) );
  INV_X1 U8557 ( .A(n8152), .ZN(n9819) );
  AOI22_X1 U8558 ( .A1(ram[3536]), .A2(n8153), .B1(n9835), .B2(n8856), .ZN(
        n8152) );
  INV_X1 U8559 ( .A(n8154), .ZN(n9820) );
  AOI22_X1 U8560 ( .A1(ram[3537]), .A2(n8153), .B1(n9835), .B2(n8880), .ZN(
        n8154) );
  INV_X1 U8561 ( .A(n8155), .ZN(n9821) );
  AOI22_X1 U8562 ( .A1(ram[3538]), .A2(n8153), .B1(n9835), .B2(n8904), .ZN(
        n8155) );
  INV_X1 U8563 ( .A(n8156), .ZN(n9822) );
  AOI22_X1 U8564 ( .A1(ram[3539]), .A2(n8153), .B1(n9835), .B2(n8928), .ZN(
        n8156) );
  INV_X1 U8565 ( .A(n8157), .ZN(n9823) );
  AOI22_X1 U8566 ( .A1(ram[3540]), .A2(n8153), .B1(n9835), .B2(n8952), .ZN(
        n8157) );
  INV_X1 U8567 ( .A(n8158), .ZN(n9824) );
  AOI22_X1 U8568 ( .A1(ram[3541]), .A2(n8153), .B1(n9835), .B2(n8976), .ZN(
        n8158) );
  INV_X1 U8569 ( .A(n8159), .ZN(n9825) );
  AOI22_X1 U8570 ( .A1(ram[3542]), .A2(n8153), .B1(n9835), .B2(n9000), .ZN(
        n8159) );
  INV_X1 U8571 ( .A(n8160), .ZN(n9826) );
  AOI22_X1 U8572 ( .A1(ram[3543]), .A2(n8153), .B1(n9835), .B2(n9024), .ZN(
        n8160) );
  INV_X1 U8573 ( .A(n8161), .ZN(n9827) );
  AOI22_X1 U8574 ( .A1(ram[3544]), .A2(n8153), .B1(n9835), .B2(n9048), .ZN(
        n8161) );
  INV_X1 U8575 ( .A(n8162), .ZN(n9828) );
  AOI22_X1 U8576 ( .A1(ram[3545]), .A2(n8153), .B1(n9835), .B2(n9072), .ZN(
        n8162) );
  INV_X1 U8577 ( .A(n8163), .ZN(n9829) );
  AOI22_X1 U8578 ( .A1(ram[3546]), .A2(n8153), .B1(n9835), .B2(n9096), .ZN(
        n8163) );
  INV_X1 U8579 ( .A(n8164), .ZN(n9830) );
  AOI22_X1 U8580 ( .A1(ram[3547]), .A2(n8153), .B1(n9835), .B2(n9120), .ZN(
        n8164) );
  INV_X1 U8581 ( .A(n8165), .ZN(n9831) );
  AOI22_X1 U8582 ( .A1(ram[3548]), .A2(n8153), .B1(n9835), .B2(n9144), .ZN(
        n8165) );
  INV_X1 U8583 ( .A(n8166), .ZN(n9832) );
  AOI22_X1 U8584 ( .A1(ram[3549]), .A2(n8153), .B1(n9835), .B2(n9168), .ZN(
        n8166) );
  INV_X1 U8585 ( .A(n8167), .ZN(n9833) );
  AOI22_X1 U8586 ( .A1(ram[3550]), .A2(n8153), .B1(n9835), .B2(n9192), .ZN(
        n8167) );
  INV_X1 U8587 ( .A(n8168), .ZN(n9834) );
  AOI22_X1 U8588 ( .A1(ram[3551]), .A2(n8153), .B1(n9835), .B2(n9216), .ZN(
        n8168) );
  INV_X1 U8589 ( .A(n8186), .ZN(n9785) );
  AOI22_X1 U8590 ( .A1(ram[3568]), .A2(n8187), .B1(n9801), .B2(n8856), .ZN(
        n8186) );
  INV_X1 U8591 ( .A(n8188), .ZN(n9786) );
  AOI22_X1 U8592 ( .A1(ram[3569]), .A2(n8187), .B1(n9801), .B2(n8880), .ZN(
        n8188) );
  INV_X1 U8593 ( .A(n8189), .ZN(n9787) );
  AOI22_X1 U8594 ( .A1(ram[3570]), .A2(n8187), .B1(n9801), .B2(n8904), .ZN(
        n8189) );
  INV_X1 U8595 ( .A(n8190), .ZN(n9788) );
  AOI22_X1 U8596 ( .A1(ram[3571]), .A2(n8187), .B1(n9801), .B2(n8928), .ZN(
        n8190) );
  INV_X1 U8597 ( .A(n8191), .ZN(n9789) );
  AOI22_X1 U8598 ( .A1(ram[3572]), .A2(n8187), .B1(n9801), .B2(n8952), .ZN(
        n8191) );
  INV_X1 U8599 ( .A(n8192), .ZN(n9790) );
  AOI22_X1 U8600 ( .A1(ram[3573]), .A2(n8187), .B1(n9801), .B2(n8976), .ZN(
        n8192) );
  INV_X1 U8601 ( .A(n8193), .ZN(n9791) );
  AOI22_X1 U8602 ( .A1(ram[3574]), .A2(n8187), .B1(n9801), .B2(n9000), .ZN(
        n8193) );
  INV_X1 U8603 ( .A(n8194), .ZN(n9792) );
  AOI22_X1 U8604 ( .A1(ram[3575]), .A2(n8187), .B1(n9801), .B2(n9024), .ZN(
        n8194) );
  INV_X1 U8605 ( .A(n8195), .ZN(n9793) );
  AOI22_X1 U8606 ( .A1(ram[3576]), .A2(n8187), .B1(n9801), .B2(n9048), .ZN(
        n8195) );
  INV_X1 U8607 ( .A(n8196), .ZN(n9794) );
  AOI22_X1 U8608 ( .A1(ram[3577]), .A2(n8187), .B1(n9801), .B2(n9072), .ZN(
        n8196) );
  INV_X1 U8609 ( .A(n8197), .ZN(n9795) );
  AOI22_X1 U8610 ( .A1(ram[3578]), .A2(n8187), .B1(n9801), .B2(n9096), .ZN(
        n8197) );
  INV_X1 U8611 ( .A(n8198), .ZN(n9796) );
  AOI22_X1 U8612 ( .A1(ram[3579]), .A2(n8187), .B1(n9801), .B2(n9120), .ZN(
        n8198) );
  INV_X1 U8613 ( .A(n8199), .ZN(n9797) );
  AOI22_X1 U8614 ( .A1(ram[3580]), .A2(n8187), .B1(n9801), .B2(n9144), .ZN(
        n8199) );
  INV_X1 U8615 ( .A(n8200), .ZN(n9798) );
  AOI22_X1 U8616 ( .A1(ram[3581]), .A2(n8187), .B1(n9801), .B2(n9168), .ZN(
        n8200) );
  INV_X1 U8617 ( .A(n8201), .ZN(n9799) );
  AOI22_X1 U8618 ( .A1(ram[3582]), .A2(n8187), .B1(n9801), .B2(n9192), .ZN(
        n8201) );
  INV_X1 U8619 ( .A(n8202), .ZN(n9800) );
  AOI22_X1 U8620 ( .A1(ram[3583]), .A2(n8187), .B1(n9801), .B2(n9216), .ZN(
        n8202) );
  INV_X1 U8621 ( .A(n8221), .ZN(n9751) );
  AOI22_X1 U8622 ( .A1(ram[3600]), .A2(n8222), .B1(n9767), .B2(n8856), .ZN(
        n8221) );
  INV_X1 U8623 ( .A(n8223), .ZN(n9752) );
  AOI22_X1 U8624 ( .A1(ram[3601]), .A2(n8222), .B1(n9767), .B2(n8880), .ZN(
        n8223) );
  INV_X1 U8625 ( .A(n8224), .ZN(n9753) );
  AOI22_X1 U8626 ( .A1(ram[3602]), .A2(n8222), .B1(n9767), .B2(n8904), .ZN(
        n8224) );
  INV_X1 U8627 ( .A(n8225), .ZN(n9754) );
  AOI22_X1 U8628 ( .A1(ram[3603]), .A2(n8222), .B1(n9767), .B2(n8928), .ZN(
        n8225) );
  INV_X1 U8629 ( .A(n8226), .ZN(n9755) );
  AOI22_X1 U8630 ( .A1(ram[3604]), .A2(n8222), .B1(n9767), .B2(n8952), .ZN(
        n8226) );
  INV_X1 U8631 ( .A(n8227), .ZN(n9756) );
  AOI22_X1 U8632 ( .A1(ram[3605]), .A2(n8222), .B1(n9767), .B2(n8976), .ZN(
        n8227) );
  INV_X1 U8633 ( .A(n8228), .ZN(n9757) );
  AOI22_X1 U8634 ( .A1(ram[3606]), .A2(n8222), .B1(n9767), .B2(n9000), .ZN(
        n8228) );
  INV_X1 U8635 ( .A(n8229), .ZN(n9758) );
  AOI22_X1 U8636 ( .A1(ram[3607]), .A2(n8222), .B1(n9767), .B2(n9024), .ZN(
        n8229) );
  INV_X1 U8637 ( .A(n8230), .ZN(n9759) );
  AOI22_X1 U8638 ( .A1(ram[3608]), .A2(n8222), .B1(n9767), .B2(n9048), .ZN(
        n8230) );
  INV_X1 U8639 ( .A(n8231), .ZN(n9760) );
  AOI22_X1 U8640 ( .A1(ram[3609]), .A2(n8222), .B1(n9767), .B2(n9072), .ZN(
        n8231) );
  INV_X1 U8641 ( .A(n8232), .ZN(n9761) );
  AOI22_X1 U8642 ( .A1(ram[3610]), .A2(n8222), .B1(n9767), .B2(n9096), .ZN(
        n8232) );
  INV_X1 U8643 ( .A(n8233), .ZN(n9762) );
  AOI22_X1 U8644 ( .A1(ram[3611]), .A2(n8222), .B1(n9767), .B2(n9120), .ZN(
        n8233) );
  INV_X1 U8645 ( .A(n8234), .ZN(n9763) );
  AOI22_X1 U8646 ( .A1(ram[3612]), .A2(n8222), .B1(n9767), .B2(n9144), .ZN(
        n8234) );
  INV_X1 U8647 ( .A(n8235), .ZN(n9764) );
  AOI22_X1 U8648 ( .A1(ram[3613]), .A2(n8222), .B1(n9767), .B2(n9168), .ZN(
        n8235) );
  INV_X1 U8649 ( .A(n8236), .ZN(n9765) );
  AOI22_X1 U8650 ( .A1(ram[3614]), .A2(n8222), .B1(n9767), .B2(n9192), .ZN(
        n8236) );
  INV_X1 U8651 ( .A(n8237), .ZN(n9766) );
  AOI22_X1 U8652 ( .A1(ram[3615]), .A2(n8222), .B1(n9767), .B2(n9216), .ZN(
        n8237) );
  INV_X1 U8653 ( .A(n8255), .ZN(n9717) );
  AOI22_X1 U8654 ( .A1(ram[3632]), .A2(n8256), .B1(n9733), .B2(n8856), .ZN(
        n8255) );
  INV_X1 U8655 ( .A(n8257), .ZN(n9718) );
  AOI22_X1 U8656 ( .A1(ram[3633]), .A2(n8256), .B1(n9733), .B2(n8880), .ZN(
        n8257) );
  INV_X1 U8657 ( .A(n8258), .ZN(n9719) );
  AOI22_X1 U8658 ( .A1(ram[3634]), .A2(n8256), .B1(n9733), .B2(n8904), .ZN(
        n8258) );
  INV_X1 U8659 ( .A(n8259), .ZN(n9720) );
  AOI22_X1 U8660 ( .A1(ram[3635]), .A2(n8256), .B1(n9733), .B2(n8928), .ZN(
        n8259) );
  INV_X1 U8661 ( .A(n8260), .ZN(n9721) );
  AOI22_X1 U8662 ( .A1(ram[3636]), .A2(n8256), .B1(n9733), .B2(n8952), .ZN(
        n8260) );
  INV_X1 U8663 ( .A(n8261), .ZN(n9722) );
  AOI22_X1 U8664 ( .A1(ram[3637]), .A2(n8256), .B1(n9733), .B2(n8976), .ZN(
        n8261) );
  INV_X1 U8665 ( .A(n8262), .ZN(n9723) );
  AOI22_X1 U8666 ( .A1(ram[3638]), .A2(n8256), .B1(n9733), .B2(n9000), .ZN(
        n8262) );
  INV_X1 U8667 ( .A(n8263), .ZN(n9724) );
  AOI22_X1 U8668 ( .A1(ram[3639]), .A2(n8256), .B1(n9733), .B2(n9024), .ZN(
        n8263) );
  INV_X1 U8669 ( .A(n8264), .ZN(n9725) );
  AOI22_X1 U8670 ( .A1(ram[3640]), .A2(n8256), .B1(n9733), .B2(n9048), .ZN(
        n8264) );
  INV_X1 U8671 ( .A(n8265), .ZN(n9726) );
  AOI22_X1 U8672 ( .A1(ram[3641]), .A2(n8256), .B1(n9733), .B2(n9072), .ZN(
        n8265) );
  INV_X1 U8673 ( .A(n8266), .ZN(n9727) );
  AOI22_X1 U8674 ( .A1(ram[3642]), .A2(n8256), .B1(n9733), .B2(n9096), .ZN(
        n8266) );
  INV_X1 U8675 ( .A(n8267), .ZN(n9728) );
  AOI22_X1 U8676 ( .A1(ram[3643]), .A2(n8256), .B1(n9733), .B2(n9120), .ZN(
        n8267) );
  INV_X1 U8677 ( .A(n8268), .ZN(n9729) );
  AOI22_X1 U8678 ( .A1(ram[3644]), .A2(n8256), .B1(n9733), .B2(n9144), .ZN(
        n8268) );
  INV_X1 U8679 ( .A(n8269), .ZN(n9730) );
  AOI22_X1 U8680 ( .A1(ram[3645]), .A2(n8256), .B1(n9733), .B2(n9168), .ZN(
        n8269) );
  INV_X1 U8681 ( .A(n8270), .ZN(n9731) );
  AOI22_X1 U8682 ( .A1(ram[3646]), .A2(n8256), .B1(n9733), .B2(n9192), .ZN(
        n8270) );
  INV_X1 U8683 ( .A(n8271), .ZN(n9732) );
  AOI22_X1 U8684 ( .A1(ram[3647]), .A2(n8256), .B1(n9733), .B2(n9216), .ZN(
        n8271) );
  INV_X1 U8685 ( .A(n8289), .ZN(n9683) );
  AOI22_X1 U8686 ( .A1(ram[3664]), .A2(n8290), .B1(n9699), .B2(n8856), .ZN(
        n8289) );
  INV_X1 U8687 ( .A(n8291), .ZN(n9684) );
  AOI22_X1 U8688 ( .A1(ram[3665]), .A2(n8290), .B1(n9699), .B2(n8880), .ZN(
        n8291) );
  INV_X1 U8689 ( .A(n8292), .ZN(n9685) );
  AOI22_X1 U8690 ( .A1(ram[3666]), .A2(n8290), .B1(n9699), .B2(n8904), .ZN(
        n8292) );
  INV_X1 U8691 ( .A(n8293), .ZN(n9686) );
  AOI22_X1 U8692 ( .A1(ram[3667]), .A2(n8290), .B1(n9699), .B2(n8928), .ZN(
        n8293) );
  INV_X1 U8693 ( .A(n8294), .ZN(n9687) );
  AOI22_X1 U8694 ( .A1(ram[3668]), .A2(n8290), .B1(n9699), .B2(n8952), .ZN(
        n8294) );
  INV_X1 U8695 ( .A(n8295), .ZN(n9688) );
  AOI22_X1 U8696 ( .A1(ram[3669]), .A2(n8290), .B1(n9699), .B2(n8976), .ZN(
        n8295) );
  INV_X1 U8697 ( .A(n8296), .ZN(n9689) );
  AOI22_X1 U8698 ( .A1(ram[3670]), .A2(n8290), .B1(n9699), .B2(n9000), .ZN(
        n8296) );
  INV_X1 U8699 ( .A(n8297), .ZN(n9690) );
  AOI22_X1 U8700 ( .A1(ram[3671]), .A2(n8290), .B1(n9699), .B2(n9024), .ZN(
        n8297) );
  INV_X1 U8701 ( .A(n8298), .ZN(n9691) );
  AOI22_X1 U8702 ( .A1(ram[3672]), .A2(n8290), .B1(n9699), .B2(n9048), .ZN(
        n8298) );
  INV_X1 U8703 ( .A(n8299), .ZN(n9692) );
  AOI22_X1 U8704 ( .A1(ram[3673]), .A2(n8290), .B1(n9699), .B2(n9072), .ZN(
        n8299) );
  INV_X1 U8705 ( .A(n8300), .ZN(n9693) );
  AOI22_X1 U8706 ( .A1(ram[3674]), .A2(n8290), .B1(n9699), .B2(n9096), .ZN(
        n8300) );
  INV_X1 U8707 ( .A(n8301), .ZN(n9694) );
  AOI22_X1 U8708 ( .A1(ram[3675]), .A2(n8290), .B1(n9699), .B2(n9120), .ZN(
        n8301) );
  INV_X1 U8709 ( .A(n8302), .ZN(n9695) );
  AOI22_X1 U8710 ( .A1(ram[3676]), .A2(n8290), .B1(n9699), .B2(n9144), .ZN(
        n8302) );
  INV_X1 U8711 ( .A(n8303), .ZN(n9696) );
  AOI22_X1 U8712 ( .A1(ram[3677]), .A2(n8290), .B1(n9699), .B2(n9168), .ZN(
        n8303) );
  INV_X1 U8713 ( .A(n8304), .ZN(n9697) );
  AOI22_X1 U8714 ( .A1(ram[3678]), .A2(n8290), .B1(n9699), .B2(n9192), .ZN(
        n8304) );
  INV_X1 U8715 ( .A(n8305), .ZN(n9698) );
  AOI22_X1 U8716 ( .A1(ram[3679]), .A2(n8290), .B1(n9699), .B2(n9216), .ZN(
        n8305) );
  INV_X1 U8717 ( .A(n8323), .ZN(n9649) );
  AOI22_X1 U8718 ( .A1(ram[3696]), .A2(n8324), .B1(n9665), .B2(n8856), .ZN(
        n8323) );
  INV_X1 U8719 ( .A(n8325), .ZN(n9650) );
  AOI22_X1 U8720 ( .A1(ram[3697]), .A2(n8324), .B1(n9665), .B2(n8880), .ZN(
        n8325) );
  INV_X1 U8721 ( .A(n8326), .ZN(n9651) );
  AOI22_X1 U8722 ( .A1(ram[3698]), .A2(n8324), .B1(n9665), .B2(n8904), .ZN(
        n8326) );
  INV_X1 U8723 ( .A(n8327), .ZN(n9652) );
  AOI22_X1 U8724 ( .A1(ram[3699]), .A2(n8324), .B1(n9665), .B2(n8928), .ZN(
        n8327) );
  INV_X1 U8725 ( .A(n8328), .ZN(n9653) );
  AOI22_X1 U8726 ( .A1(ram[3700]), .A2(n8324), .B1(n9665), .B2(n8952), .ZN(
        n8328) );
  INV_X1 U8727 ( .A(n8329), .ZN(n9654) );
  AOI22_X1 U8728 ( .A1(ram[3701]), .A2(n8324), .B1(n9665), .B2(n8976), .ZN(
        n8329) );
  INV_X1 U8729 ( .A(n8330), .ZN(n9655) );
  AOI22_X1 U8730 ( .A1(ram[3702]), .A2(n8324), .B1(n9665), .B2(n9000), .ZN(
        n8330) );
  INV_X1 U8731 ( .A(n8331), .ZN(n9656) );
  AOI22_X1 U8732 ( .A1(ram[3703]), .A2(n8324), .B1(n9665), .B2(n9024), .ZN(
        n8331) );
  INV_X1 U8733 ( .A(n8332), .ZN(n9657) );
  AOI22_X1 U8734 ( .A1(ram[3704]), .A2(n8324), .B1(n9665), .B2(n9048), .ZN(
        n8332) );
  INV_X1 U8735 ( .A(n8333), .ZN(n9658) );
  AOI22_X1 U8736 ( .A1(ram[3705]), .A2(n8324), .B1(n9665), .B2(n9072), .ZN(
        n8333) );
  INV_X1 U8737 ( .A(n8334), .ZN(n9659) );
  AOI22_X1 U8738 ( .A1(ram[3706]), .A2(n8324), .B1(n9665), .B2(n9096), .ZN(
        n8334) );
  INV_X1 U8739 ( .A(n8335), .ZN(n9660) );
  AOI22_X1 U8740 ( .A1(ram[3707]), .A2(n8324), .B1(n9665), .B2(n9120), .ZN(
        n8335) );
  INV_X1 U8741 ( .A(n8336), .ZN(n9661) );
  AOI22_X1 U8742 ( .A1(ram[3708]), .A2(n8324), .B1(n9665), .B2(n9144), .ZN(
        n8336) );
  INV_X1 U8743 ( .A(n8337), .ZN(n9662) );
  AOI22_X1 U8744 ( .A1(ram[3709]), .A2(n8324), .B1(n9665), .B2(n9168), .ZN(
        n8337) );
  INV_X1 U8745 ( .A(n8338), .ZN(n9663) );
  AOI22_X1 U8746 ( .A1(ram[3710]), .A2(n8324), .B1(n9665), .B2(n9192), .ZN(
        n8338) );
  INV_X1 U8747 ( .A(n8339), .ZN(n9664) );
  AOI22_X1 U8748 ( .A1(ram[3711]), .A2(n8324), .B1(n9665), .B2(n9216), .ZN(
        n8339) );
  INV_X1 U8749 ( .A(n8357), .ZN(n9615) );
  AOI22_X1 U8750 ( .A1(ram[3728]), .A2(n8358), .B1(n9631), .B2(n8855), .ZN(
        n8357) );
  INV_X1 U8751 ( .A(n8359), .ZN(n9616) );
  AOI22_X1 U8752 ( .A1(ram[3729]), .A2(n8358), .B1(n9631), .B2(n8879), .ZN(
        n8359) );
  INV_X1 U8753 ( .A(n8360), .ZN(n9617) );
  AOI22_X1 U8754 ( .A1(ram[3730]), .A2(n8358), .B1(n9631), .B2(n8903), .ZN(
        n8360) );
  INV_X1 U8755 ( .A(n8361), .ZN(n9618) );
  AOI22_X1 U8756 ( .A1(ram[3731]), .A2(n8358), .B1(n9631), .B2(n8927), .ZN(
        n8361) );
  INV_X1 U8757 ( .A(n8362), .ZN(n9619) );
  AOI22_X1 U8758 ( .A1(ram[3732]), .A2(n8358), .B1(n9631), .B2(n8951), .ZN(
        n8362) );
  INV_X1 U8759 ( .A(n8363), .ZN(n9620) );
  AOI22_X1 U8760 ( .A1(ram[3733]), .A2(n8358), .B1(n9631), .B2(n8975), .ZN(
        n8363) );
  INV_X1 U8761 ( .A(n8364), .ZN(n9621) );
  AOI22_X1 U8762 ( .A1(ram[3734]), .A2(n8358), .B1(n9631), .B2(n8999), .ZN(
        n8364) );
  INV_X1 U8763 ( .A(n8365), .ZN(n9622) );
  AOI22_X1 U8764 ( .A1(ram[3735]), .A2(n8358), .B1(n9631), .B2(n9023), .ZN(
        n8365) );
  INV_X1 U8765 ( .A(n8366), .ZN(n9623) );
  AOI22_X1 U8766 ( .A1(ram[3736]), .A2(n8358), .B1(n9631), .B2(n9047), .ZN(
        n8366) );
  INV_X1 U8767 ( .A(n8367), .ZN(n9624) );
  AOI22_X1 U8768 ( .A1(ram[3737]), .A2(n8358), .B1(n9631), .B2(n9071), .ZN(
        n8367) );
  INV_X1 U8769 ( .A(n8368), .ZN(n9625) );
  AOI22_X1 U8770 ( .A1(ram[3738]), .A2(n8358), .B1(n9631), .B2(n9095), .ZN(
        n8368) );
  INV_X1 U8771 ( .A(n8369), .ZN(n9626) );
  AOI22_X1 U8772 ( .A1(ram[3739]), .A2(n8358), .B1(n9631), .B2(n9119), .ZN(
        n8369) );
  INV_X1 U8773 ( .A(n8370), .ZN(n9627) );
  AOI22_X1 U8774 ( .A1(ram[3740]), .A2(n8358), .B1(n9631), .B2(n9143), .ZN(
        n8370) );
  INV_X1 U8775 ( .A(n8371), .ZN(n9628) );
  AOI22_X1 U8776 ( .A1(ram[3741]), .A2(n8358), .B1(n9631), .B2(n9167), .ZN(
        n8371) );
  INV_X1 U8777 ( .A(n8372), .ZN(n9629) );
  AOI22_X1 U8778 ( .A1(ram[3742]), .A2(n8358), .B1(n9631), .B2(n9191), .ZN(
        n8372) );
  INV_X1 U8779 ( .A(n8373), .ZN(n9630) );
  AOI22_X1 U8780 ( .A1(ram[3743]), .A2(n8358), .B1(n9631), .B2(n9215), .ZN(
        n8373) );
  INV_X1 U8781 ( .A(n8391), .ZN(n9581) );
  AOI22_X1 U8782 ( .A1(ram[3760]), .A2(n8392), .B1(n9597), .B2(n8855), .ZN(
        n8391) );
  INV_X1 U8783 ( .A(n8393), .ZN(n9582) );
  AOI22_X1 U8784 ( .A1(ram[3761]), .A2(n8392), .B1(n9597), .B2(n8879), .ZN(
        n8393) );
  INV_X1 U8785 ( .A(n8394), .ZN(n9583) );
  AOI22_X1 U8786 ( .A1(ram[3762]), .A2(n8392), .B1(n9597), .B2(n8903), .ZN(
        n8394) );
  INV_X1 U8787 ( .A(n8395), .ZN(n9584) );
  AOI22_X1 U8788 ( .A1(ram[3763]), .A2(n8392), .B1(n9597), .B2(n8927), .ZN(
        n8395) );
  INV_X1 U8789 ( .A(n8396), .ZN(n9585) );
  AOI22_X1 U8790 ( .A1(ram[3764]), .A2(n8392), .B1(n9597), .B2(n8951), .ZN(
        n8396) );
  INV_X1 U8791 ( .A(n8397), .ZN(n9586) );
  AOI22_X1 U8792 ( .A1(ram[3765]), .A2(n8392), .B1(n9597), .B2(n8975), .ZN(
        n8397) );
  INV_X1 U8793 ( .A(n8398), .ZN(n9587) );
  AOI22_X1 U8794 ( .A1(ram[3766]), .A2(n8392), .B1(n9597), .B2(n8999), .ZN(
        n8398) );
  INV_X1 U8795 ( .A(n8399), .ZN(n9588) );
  AOI22_X1 U8796 ( .A1(ram[3767]), .A2(n8392), .B1(n9597), .B2(n9023), .ZN(
        n8399) );
  INV_X1 U8797 ( .A(n8400), .ZN(n9589) );
  AOI22_X1 U8798 ( .A1(ram[3768]), .A2(n8392), .B1(n9597), .B2(n9047), .ZN(
        n8400) );
  INV_X1 U8799 ( .A(n8401), .ZN(n9590) );
  AOI22_X1 U8800 ( .A1(ram[3769]), .A2(n8392), .B1(n9597), .B2(n9071), .ZN(
        n8401) );
  INV_X1 U8801 ( .A(n8402), .ZN(n9591) );
  AOI22_X1 U8802 ( .A1(ram[3770]), .A2(n8392), .B1(n9597), .B2(n9095), .ZN(
        n8402) );
  INV_X1 U8803 ( .A(n8403), .ZN(n9592) );
  AOI22_X1 U8804 ( .A1(ram[3771]), .A2(n8392), .B1(n9597), .B2(n9119), .ZN(
        n8403) );
  INV_X1 U8805 ( .A(n8404), .ZN(n9593) );
  AOI22_X1 U8806 ( .A1(ram[3772]), .A2(n8392), .B1(n9597), .B2(n9143), .ZN(
        n8404) );
  INV_X1 U8807 ( .A(n8405), .ZN(n9594) );
  AOI22_X1 U8808 ( .A1(ram[3773]), .A2(n8392), .B1(n9597), .B2(n9167), .ZN(
        n8405) );
  INV_X1 U8809 ( .A(n8406), .ZN(n9595) );
  AOI22_X1 U8810 ( .A1(ram[3774]), .A2(n8392), .B1(n9597), .B2(n9191), .ZN(
        n8406) );
  INV_X1 U8811 ( .A(n8407), .ZN(n9596) );
  AOI22_X1 U8812 ( .A1(ram[3775]), .A2(n8392), .B1(n9597), .B2(n9215), .ZN(
        n8407) );
  INV_X1 U8813 ( .A(n8425), .ZN(n9547) );
  AOI22_X1 U8814 ( .A1(ram[3792]), .A2(n8426), .B1(n9563), .B2(n8855), .ZN(
        n8425) );
  INV_X1 U8815 ( .A(n8427), .ZN(n9548) );
  AOI22_X1 U8816 ( .A1(ram[3793]), .A2(n8426), .B1(n9563), .B2(n8879), .ZN(
        n8427) );
  INV_X1 U8817 ( .A(n8428), .ZN(n9549) );
  AOI22_X1 U8818 ( .A1(ram[3794]), .A2(n8426), .B1(n9563), .B2(n8903), .ZN(
        n8428) );
  INV_X1 U8819 ( .A(n8429), .ZN(n9550) );
  AOI22_X1 U8820 ( .A1(ram[3795]), .A2(n8426), .B1(n9563), .B2(n8927), .ZN(
        n8429) );
  INV_X1 U8821 ( .A(n8430), .ZN(n9551) );
  AOI22_X1 U8822 ( .A1(ram[3796]), .A2(n8426), .B1(n9563), .B2(n8951), .ZN(
        n8430) );
  INV_X1 U8823 ( .A(n8431), .ZN(n9552) );
  AOI22_X1 U8824 ( .A1(ram[3797]), .A2(n8426), .B1(n9563), .B2(n8975), .ZN(
        n8431) );
  INV_X1 U8825 ( .A(n8432), .ZN(n9553) );
  AOI22_X1 U8826 ( .A1(ram[3798]), .A2(n8426), .B1(n9563), .B2(n8999), .ZN(
        n8432) );
  INV_X1 U8827 ( .A(n8433), .ZN(n9554) );
  AOI22_X1 U8828 ( .A1(ram[3799]), .A2(n8426), .B1(n9563), .B2(n9023), .ZN(
        n8433) );
  INV_X1 U8829 ( .A(n8434), .ZN(n9555) );
  AOI22_X1 U8830 ( .A1(ram[3800]), .A2(n8426), .B1(n9563), .B2(n9047), .ZN(
        n8434) );
  INV_X1 U8831 ( .A(n8435), .ZN(n9556) );
  AOI22_X1 U8832 ( .A1(ram[3801]), .A2(n8426), .B1(n9563), .B2(n9071), .ZN(
        n8435) );
  INV_X1 U8833 ( .A(n8436), .ZN(n9557) );
  AOI22_X1 U8834 ( .A1(ram[3802]), .A2(n8426), .B1(n9563), .B2(n9095), .ZN(
        n8436) );
  INV_X1 U8835 ( .A(n8437), .ZN(n9558) );
  AOI22_X1 U8836 ( .A1(ram[3803]), .A2(n8426), .B1(n9563), .B2(n9119), .ZN(
        n8437) );
  INV_X1 U8837 ( .A(n8438), .ZN(n9559) );
  AOI22_X1 U8838 ( .A1(ram[3804]), .A2(n8426), .B1(n9563), .B2(n9143), .ZN(
        n8438) );
  INV_X1 U8839 ( .A(n8439), .ZN(n9560) );
  AOI22_X1 U8840 ( .A1(ram[3805]), .A2(n8426), .B1(n9563), .B2(n9167), .ZN(
        n8439) );
  INV_X1 U8841 ( .A(n8440), .ZN(n9561) );
  AOI22_X1 U8842 ( .A1(ram[3806]), .A2(n8426), .B1(n9563), .B2(n9191), .ZN(
        n8440) );
  INV_X1 U8843 ( .A(n8441), .ZN(n9562) );
  AOI22_X1 U8844 ( .A1(ram[3807]), .A2(n8426), .B1(n9563), .B2(n9215), .ZN(
        n8441) );
  INV_X1 U8845 ( .A(n8459), .ZN(n9513) );
  AOI22_X1 U8846 ( .A1(ram[3824]), .A2(n8460), .B1(n9529), .B2(n8855), .ZN(
        n8459) );
  INV_X1 U8847 ( .A(n8461), .ZN(n9514) );
  AOI22_X1 U8848 ( .A1(ram[3825]), .A2(n8460), .B1(n9529), .B2(n8879), .ZN(
        n8461) );
  INV_X1 U8849 ( .A(n8462), .ZN(n9515) );
  AOI22_X1 U8850 ( .A1(ram[3826]), .A2(n8460), .B1(n9529), .B2(n8903), .ZN(
        n8462) );
  INV_X1 U8851 ( .A(n8463), .ZN(n9516) );
  AOI22_X1 U8852 ( .A1(ram[3827]), .A2(n8460), .B1(n9529), .B2(n8927), .ZN(
        n8463) );
  INV_X1 U8853 ( .A(n8464), .ZN(n9517) );
  AOI22_X1 U8854 ( .A1(ram[3828]), .A2(n8460), .B1(n9529), .B2(n8951), .ZN(
        n8464) );
  INV_X1 U8855 ( .A(n8465), .ZN(n9518) );
  AOI22_X1 U8856 ( .A1(ram[3829]), .A2(n8460), .B1(n9529), .B2(n8975), .ZN(
        n8465) );
  INV_X1 U8857 ( .A(n8466), .ZN(n9519) );
  AOI22_X1 U8858 ( .A1(ram[3830]), .A2(n8460), .B1(n9529), .B2(n8999), .ZN(
        n8466) );
  INV_X1 U8859 ( .A(n8467), .ZN(n9520) );
  AOI22_X1 U8860 ( .A1(ram[3831]), .A2(n8460), .B1(n9529), .B2(n9023), .ZN(
        n8467) );
  INV_X1 U8861 ( .A(n8468), .ZN(n9521) );
  AOI22_X1 U8862 ( .A1(ram[3832]), .A2(n8460), .B1(n9529), .B2(n9047), .ZN(
        n8468) );
  INV_X1 U8863 ( .A(n8469), .ZN(n9522) );
  AOI22_X1 U8864 ( .A1(ram[3833]), .A2(n8460), .B1(n9529), .B2(n9071), .ZN(
        n8469) );
  INV_X1 U8865 ( .A(n8470), .ZN(n9523) );
  AOI22_X1 U8866 ( .A1(ram[3834]), .A2(n8460), .B1(n9529), .B2(n9095), .ZN(
        n8470) );
  INV_X1 U8867 ( .A(n8471), .ZN(n9524) );
  AOI22_X1 U8868 ( .A1(ram[3835]), .A2(n8460), .B1(n9529), .B2(n9119), .ZN(
        n8471) );
  INV_X1 U8869 ( .A(n8472), .ZN(n9525) );
  AOI22_X1 U8870 ( .A1(ram[3836]), .A2(n8460), .B1(n9529), .B2(n9143), .ZN(
        n8472) );
  INV_X1 U8871 ( .A(n8473), .ZN(n9526) );
  AOI22_X1 U8872 ( .A1(ram[3837]), .A2(n8460), .B1(n9529), .B2(n9167), .ZN(
        n8473) );
  INV_X1 U8873 ( .A(n8474), .ZN(n9527) );
  AOI22_X1 U8874 ( .A1(ram[3838]), .A2(n8460), .B1(n9529), .B2(n9191), .ZN(
        n8474) );
  INV_X1 U8875 ( .A(n8475), .ZN(n9528) );
  AOI22_X1 U8876 ( .A1(ram[3839]), .A2(n8460), .B1(n9529), .B2(n9215), .ZN(
        n8475) );
  INV_X1 U8877 ( .A(n8496), .ZN(n9479) );
  AOI22_X1 U8878 ( .A1(ram[3856]), .A2(n8497), .B1(n9495), .B2(n8855), .ZN(
        n8496) );
  INV_X1 U8879 ( .A(n8498), .ZN(n9480) );
  AOI22_X1 U8880 ( .A1(ram[3857]), .A2(n8497), .B1(n9495), .B2(n8879), .ZN(
        n8498) );
  INV_X1 U8881 ( .A(n8499), .ZN(n9481) );
  AOI22_X1 U8882 ( .A1(ram[3858]), .A2(n8497), .B1(n9495), .B2(n8903), .ZN(
        n8499) );
  INV_X1 U8883 ( .A(n8500), .ZN(n9482) );
  AOI22_X1 U8884 ( .A1(ram[3859]), .A2(n8497), .B1(n9495), .B2(n8927), .ZN(
        n8500) );
  INV_X1 U8885 ( .A(n8501), .ZN(n9483) );
  AOI22_X1 U8886 ( .A1(ram[3860]), .A2(n8497), .B1(n9495), .B2(n8951), .ZN(
        n8501) );
  INV_X1 U8887 ( .A(n8502), .ZN(n9484) );
  AOI22_X1 U8888 ( .A1(ram[3861]), .A2(n8497), .B1(n9495), .B2(n8975), .ZN(
        n8502) );
  INV_X1 U8889 ( .A(n8503), .ZN(n9485) );
  AOI22_X1 U8890 ( .A1(ram[3862]), .A2(n8497), .B1(n9495), .B2(n8999), .ZN(
        n8503) );
  INV_X1 U8891 ( .A(n8504), .ZN(n9486) );
  AOI22_X1 U8892 ( .A1(ram[3863]), .A2(n8497), .B1(n9495), .B2(n9023), .ZN(
        n8504) );
  INV_X1 U8893 ( .A(n8505), .ZN(n9487) );
  AOI22_X1 U8894 ( .A1(ram[3864]), .A2(n8497), .B1(n9495), .B2(n9047), .ZN(
        n8505) );
  INV_X1 U8895 ( .A(n8506), .ZN(n9488) );
  AOI22_X1 U8896 ( .A1(ram[3865]), .A2(n8497), .B1(n9495), .B2(n9071), .ZN(
        n8506) );
  INV_X1 U8897 ( .A(n8507), .ZN(n9489) );
  AOI22_X1 U8898 ( .A1(ram[3866]), .A2(n8497), .B1(n9495), .B2(n9095), .ZN(
        n8507) );
  INV_X1 U8899 ( .A(n8508), .ZN(n9490) );
  AOI22_X1 U8900 ( .A1(ram[3867]), .A2(n8497), .B1(n9495), .B2(n9119), .ZN(
        n8508) );
  INV_X1 U8901 ( .A(n8509), .ZN(n9491) );
  AOI22_X1 U8902 ( .A1(ram[3868]), .A2(n8497), .B1(n9495), .B2(n9143), .ZN(
        n8509) );
  INV_X1 U8903 ( .A(n8510), .ZN(n9492) );
  AOI22_X1 U8904 ( .A1(ram[3869]), .A2(n8497), .B1(n9495), .B2(n9167), .ZN(
        n8510) );
  INV_X1 U8905 ( .A(n8511), .ZN(n9493) );
  AOI22_X1 U8906 ( .A1(ram[3870]), .A2(n8497), .B1(n9495), .B2(n9191), .ZN(
        n8511) );
  INV_X1 U8907 ( .A(n8512), .ZN(n9494) );
  AOI22_X1 U8908 ( .A1(ram[3871]), .A2(n8497), .B1(n9495), .B2(n9215), .ZN(
        n8512) );
  INV_X1 U8909 ( .A(n8532), .ZN(n9445) );
  AOI22_X1 U8910 ( .A1(ram[3888]), .A2(n8533), .B1(n9461), .B2(n8855), .ZN(
        n8532) );
  INV_X1 U8911 ( .A(n8534), .ZN(n9446) );
  AOI22_X1 U8912 ( .A1(ram[3889]), .A2(n8533), .B1(n9461), .B2(n8879), .ZN(
        n8534) );
  INV_X1 U8913 ( .A(n8535), .ZN(n9447) );
  AOI22_X1 U8914 ( .A1(ram[3890]), .A2(n8533), .B1(n9461), .B2(n8903), .ZN(
        n8535) );
  INV_X1 U8915 ( .A(n8536), .ZN(n9448) );
  AOI22_X1 U8916 ( .A1(ram[3891]), .A2(n8533), .B1(n9461), .B2(n8927), .ZN(
        n8536) );
  INV_X1 U8917 ( .A(n8537), .ZN(n9449) );
  AOI22_X1 U8918 ( .A1(ram[3892]), .A2(n8533), .B1(n9461), .B2(n8951), .ZN(
        n8537) );
  INV_X1 U8919 ( .A(n8538), .ZN(n9450) );
  AOI22_X1 U8920 ( .A1(ram[3893]), .A2(n8533), .B1(n9461), .B2(n8975), .ZN(
        n8538) );
  INV_X1 U8921 ( .A(n8539), .ZN(n9451) );
  AOI22_X1 U8922 ( .A1(ram[3894]), .A2(n8533), .B1(n9461), .B2(n8999), .ZN(
        n8539) );
  INV_X1 U8923 ( .A(n8540), .ZN(n9452) );
  AOI22_X1 U8924 ( .A1(ram[3895]), .A2(n8533), .B1(n9461), .B2(n9023), .ZN(
        n8540) );
  INV_X1 U8925 ( .A(n8541), .ZN(n9453) );
  AOI22_X1 U8926 ( .A1(ram[3896]), .A2(n8533), .B1(n9461), .B2(n9047), .ZN(
        n8541) );
  INV_X1 U8927 ( .A(n8542), .ZN(n9454) );
  AOI22_X1 U8928 ( .A1(ram[3897]), .A2(n8533), .B1(n9461), .B2(n9071), .ZN(
        n8542) );
  INV_X1 U8929 ( .A(n8543), .ZN(n9455) );
  AOI22_X1 U8930 ( .A1(ram[3898]), .A2(n8533), .B1(n9461), .B2(n9095), .ZN(
        n8543) );
  INV_X1 U8931 ( .A(n8544), .ZN(n9456) );
  AOI22_X1 U8932 ( .A1(ram[3899]), .A2(n8533), .B1(n9461), .B2(n9119), .ZN(
        n8544) );
  INV_X1 U8933 ( .A(n8545), .ZN(n9457) );
  AOI22_X1 U8934 ( .A1(ram[3900]), .A2(n8533), .B1(n9461), .B2(n9143), .ZN(
        n8545) );
  INV_X1 U8935 ( .A(n8546), .ZN(n9458) );
  AOI22_X1 U8936 ( .A1(ram[3901]), .A2(n8533), .B1(n9461), .B2(n9167), .ZN(
        n8546) );
  INV_X1 U8937 ( .A(n8547), .ZN(n9459) );
  AOI22_X1 U8938 ( .A1(ram[3902]), .A2(n8533), .B1(n9461), .B2(n9191), .ZN(
        n8547) );
  INV_X1 U8939 ( .A(n8548), .ZN(n9460) );
  AOI22_X1 U8940 ( .A1(ram[3903]), .A2(n8533), .B1(n9461), .B2(n9215), .ZN(
        n8548) );
  INV_X1 U8941 ( .A(n8568), .ZN(n9411) );
  AOI22_X1 U8942 ( .A1(ram[3920]), .A2(n8569), .B1(n9427), .B2(n8854), .ZN(
        n8568) );
  INV_X1 U8943 ( .A(n8570), .ZN(n9412) );
  AOI22_X1 U8944 ( .A1(ram[3921]), .A2(n8569), .B1(n9427), .B2(n8878), .ZN(
        n8570) );
  INV_X1 U8945 ( .A(n8571), .ZN(n9413) );
  AOI22_X1 U8946 ( .A1(ram[3922]), .A2(n8569), .B1(n9427), .B2(n8902), .ZN(
        n8571) );
  INV_X1 U8947 ( .A(n8572), .ZN(n9414) );
  AOI22_X1 U8948 ( .A1(ram[3923]), .A2(n8569), .B1(n9427), .B2(n8926), .ZN(
        n8572) );
  INV_X1 U8949 ( .A(n8573), .ZN(n9415) );
  AOI22_X1 U8950 ( .A1(ram[3924]), .A2(n8569), .B1(n9427), .B2(n8950), .ZN(
        n8573) );
  INV_X1 U8951 ( .A(n8574), .ZN(n9416) );
  AOI22_X1 U8952 ( .A1(ram[3925]), .A2(n8569), .B1(n9427), .B2(n8974), .ZN(
        n8574) );
  INV_X1 U8953 ( .A(n8575), .ZN(n9417) );
  AOI22_X1 U8954 ( .A1(ram[3926]), .A2(n8569), .B1(n9427), .B2(n8998), .ZN(
        n8575) );
  INV_X1 U8955 ( .A(n8576), .ZN(n9418) );
  AOI22_X1 U8956 ( .A1(ram[3927]), .A2(n8569), .B1(n9427), .B2(n9022), .ZN(
        n8576) );
  INV_X1 U8957 ( .A(n8577), .ZN(n9419) );
  AOI22_X1 U8958 ( .A1(ram[3928]), .A2(n8569), .B1(n9427), .B2(n9046), .ZN(
        n8577) );
  INV_X1 U8959 ( .A(n8578), .ZN(n9420) );
  AOI22_X1 U8960 ( .A1(ram[3929]), .A2(n8569), .B1(n9427), .B2(n9070), .ZN(
        n8578) );
  INV_X1 U8961 ( .A(n8579), .ZN(n9421) );
  AOI22_X1 U8962 ( .A1(ram[3930]), .A2(n8569), .B1(n9427), .B2(n9094), .ZN(
        n8579) );
  INV_X1 U8963 ( .A(n8580), .ZN(n9422) );
  AOI22_X1 U8964 ( .A1(ram[3931]), .A2(n8569), .B1(n9427), .B2(n9118), .ZN(
        n8580) );
  INV_X1 U8965 ( .A(n8581), .ZN(n9423) );
  AOI22_X1 U8966 ( .A1(ram[3932]), .A2(n8569), .B1(n9427), .B2(n9142), .ZN(
        n8581) );
  INV_X1 U8967 ( .A(n8582), .ZN(n9424) );
  AOI22_X1 U8968 ( .A1(ram[3933]), .A2(n8569), .B1(n9427), .B2(n9166), .ZN(
        n8582) );
  INV_X1 U8969 ( .A(n8583), .ZN(n9425) );
  AOI22_X1 U8970 ( .A1(ram[3934]), .A2(n8569), .B1(n9427), .B2(n9190), .ZN(
        n8583) );
  INV_X1 U8971 ( .A(n8584), .ZN(n9426) );
  AOI22_X1 U8972 ( .A1(ram[3935]), .A2(n8569), .B1(n9427), .B2(n9214), .ZN(
        n8584) );
  INV_X1 U8973 ( .A(n8602), .ZN(n9377) );
  AOI22_X1 U8974 ( .A1(ram[3952]), .A2(n8603), .B1(n9393), .B2(n8854), .ZN(
        n8602) );
  INV_X1 U8975 ( .A(n8604), .ZN(n9378) );
  AOI22_X1 U8976 ( .A1(ram[3953]), .A2(n8603), .B1(n9393), .B2(n8878), .ZN(
        n8604) );
  INV_X1 U8977 ( .A(n8605), .ZN(n9379) );
  AOI22_X1 U8978 ( .A1(ram[3954]), .A2(n8603), .B1(n9393), .B2(n8902), .ZN(
        n8605) );
  INV_X1 U8979 ( .A(n8606), .ZN(n9380) );
  AOI22_X1 U8980 ( .A1(ram[3955]), .A2(n8603), .B1(n9393), .B2(n8926), .ZN(
        n8606) );
  INV_X1 U8981 ( .A(n8607), .ZN(n9381) );
  AOI22_X1 U8982 ( .A1(ram[3956]), .A2(n8603), .B1(n9393), .B2(n8950), .ZN(
        n8607) );
  INV_X1 U8983 ( .A(n8608), .ZN(n9382) );
  AOI22_X1 U8984 ( .A1(ram[3957]), .A2(n8603), .B1(n9393), .B2(n8974), .ZN(
        n8608) );
  INV_X1 U8985 ( .A(n8609), .ZN(n9383) );
  AOI22_X1 U8986 ( .A1(ram[3958]), .A2(n8603), .B1(n9393), .B2(n8998), .ZN(
        n8609) );
  INV_X1 U8987 ( .A(n8610), .ZN(n9384) );
  AOI22_X1 U8988 ( .A1(ram[3959]), .A2(n8603), .B1(n9393), .B2(n9022), .ZN(
        n8610) );
  INV_X1 U8989 ( .A(n8611), .ZN(n9385) );
  AOI22_X1 U8990 ( .A1(ram[3960]), .A2(n8603), .B1(n9393), .B2(n9046), .ZN(
        n8611) );
  INV_X1 U8991 ( .A(n8612), .ZN(n9386) );
  AOI22_X1 U8992 ( .A1(ram[3961]), .A2(n8603), .B1(n9393), .B2(n9070), .ZN(
        n8612) );
  INV_X1 U8993 ( .A(n8613), .ZN(n9387) );
  AOI22_X1 U8994 ( .A1(ram[3962]), .A2(n8603), .B1(n9393), .B2(n9094), .ZN(
        n8613) );
  INV_X1 U8995 ( .A(n8614), .ZN(n9388) );
  AOI22_X1 U8996 ( .A1(ram[3963]), .A2(n8603), .B1(n9393), .B2(n9118), .ZN(
        n8614) );
  INV_X1 U8997 ( .A(n8615), .ZN(n9389) );
  AOI22_X1 U8998 ( .A1(ram[3964]), .A2(n8603), .B1(n9393), .B2(n9142), .ZN(
        n8615) );
  INV_X1 U8999 ( .A(n8616), .ZN(n9390) );
  AOI22_X1 U9000 ( .A1(ram[3965]), .A2(n8603), .B1(n9393), .B2(n9166), .ZN(
        n8616) );
  INV_X1 U9001 ( .A(n8617), .ZN(n9391) );
  AOI22_X1 U9002 ( .A1(ram[3966]), .A2(n8603), .B1(n9393), .B2(n9190), .ZN(
        n8617) );
  INV_X1 U9003 ( .A(n8618), .ZN(n9392) );
  AOI22_X1 U9004 ( .A1(ram[3967]), .A2(n8603), .B1(n9393), .B2(n9214), .ZN(
        n8618) );
  INV_X1 U9005 ( .A(n8637), .ZN(n9343) );
  AOI22_X1 U9006 ( .A1(ram[3984]), .A2(n8638), .B1(n9359), .B2(n8854), .ZN(
        n8637) );
  INV_X1 U9007 ( .A(n8639), .ZN(n9344) );
  AOI22_X1 U9008 ( .A1(ram[3985]), .A2(n8638), .B1(n9359), .B2(n8878), .ZN(
        n8639) );
  INV_X1 U9009 ( .A(n8640), .ZN(n9345) );
  AOI22_X1 U9010 ( .A1(ram[3986]), .A2(n8638), .B1(n9359), .B2(n8902), .ZN(
        n8640) );
  INV_X1 U9011 ( .A(n8641), .ZN(n9346) );
  AOI22_X1 U9012 ( .A1(ram[3987]), .A2(n8638), .B1(n9359), .B2(n8926), .ZN(
        n8641) );
  INV_X1 U9013 ( .A(n8642), .ZN(n9347) );
  AOI22_X1 U9014 ( .A1(ram[3988]), .A2(n8638), .B1(n9359), .B2(n8950), .ZN(
        n8642) );
  INV_X1 U9015 ( .A(n8643), .ZN(n9348) );
  AOI22_X1 U9016 ( .A1(ram[3989]), .A2(n8638), .B1(n9359), .B2(n8974), .ZN(
        n8643) );
  INV_X1 U9017 ( .A(n8644), .ZN(n9349) );
  AOI22_X1 U9018 ( .A1(ram[3990]), .A2(n8638), .B1(n9359), .B2(n8998), .ZN(
        n8644) );
  INV_X1 U9019 ( .A(n8645), .ZN(n9350) );
  AOI22_X1 U9020 ( .A1(ram[3991]), .A2(n8638), .B1(n9359), .B2(n9022), .ZN(
        n8645) );
  INV_X1 U9021 ( .A(n8646), .ZN(n9351) );
  AOI22_X1 U9022 ( .A1(ram[3992]), .A2(n8638), .B1(n9359), .B2(n9046), .ZN(
        n8646) );
  INV_X1 U9023 ( .A(n8647), .ZN(n9352) );
  AOI22_X1 U9024 ( .A1(ram[3993]), .A2(n8638), .B1(n9359), .B2(n9070), .ZN(
        n8647) );
  INV_X1 U9025 ( .A(n8648), .ZN(n9353) );
  AOI22_X1 U9026 ( .A1(ram[3994]), .A2(n8638), .B1(n9359), .B2(n9094), .ZN(
        n8648) );
  INV_X1 U9027 ( .A(n8649), .ZN(n9354) );
  AOI22_X1 U9028 ( .A1(ram[3995]), .A2(n8638), .B1(n9359), .B2(n9118), .ZN(
        n8649) );
  INV_X1 U9029 ( .A(n8650), .ZN(n9355) );
  AOI22_X1 U9030 ( .A1(ram[3996]), .A2(n8638), .B1(n9359), .B2(n9142), .ZN(
        n8650) );
  INV_X1 U9031 ( .A(n8651), .ZN(n9356) );
  AOI22_X1 U9032 ( .A1(ram[3997]), .A2(n8638), .B1(n9359), .B2(n9166), .ZN(
        n8651) );
  INV_X1 U9033 ( .A(n8652), .ZN(n9357) );
  AOI22_X1 U9034 ( .A1(ram[3998]), .A2(n8638), .B1(n9359), .B2(n9190), .ZN(
        n8652) );
  INV_X1 U9035 ( .A(n8653), .ZN(n9358) );
  AOI22_X1 U9036 ( .A1(ram[3999]), .A2(n8638), .B1(n9359), .B2(n9214), .ZN(
        n8653) );
  INV_X1 U9037 ( .A(n8671), .ZN(n9309) );
  AOI22_X1 U9038 ( .A1(ram[4016]), .A2(n8672), .B1(n9325), .B2(n8854), .ZN(
        n8671) );
  INV_X1 U9039 ( .A(n8673), .ZN(n9310) );
  AOI22_X1 U9040 ( .A1(ram[4017]), .A2(n8672), .B1(n9325), .B2(n8878), .ZN(
        n8673) );
  INV_X1 U9041 ( .A(n8674), .ZN(n9311) );
  AOI22_X1 U9042 ( .A1(ram[4018]), .A2(n8672), .B1(n9325), .B2(n8902), .ZN(
        n8674) );
  INV_X1 U9043 ( .A(n8675), .ZN(n9312) );
  AOI22_X1 U9044 ( .A1(ram[4019]), .A2(n8672), .B1(n9325), .B2(n8926), .ZN(
        n8675) );
  INV_X1 U9045 ( .A(n8676), .ZN(n9313) );
  AOI22_X1 U9046 ( .A1(ram[4020]), .A2(n8672), .B1(n9325), .B2(n8950), .ZN(
        n8676) );
  INV_X1 U9047 ( .A(n8677), .ZN(n9314) );
  AOI22_X1 U9048 ( .A1(ram[4021]), .A2(n8672), .B1(n9325), .B2(n8974), .ZN(
        n8677) );
  INV_X1 U9049 ( .A(n8678), .ZN(n9315) );
  AOI22_X1 U9050 ( .A1(ram[4022]), .A2(n8672), .B1(n9325), .B2(n8998), .ZN(
        n8678) );
  INV_X1 U9051 ( .A(n8679), .ZN(n9316) );
  AOI22_X1 U9052 ( .A1(ram[4023]), .A2(n8672), .B1(n9325), .B2(n9022), .ZN(
        n8679) );
  INV_X1 U9053 ( .A(n8680), .ZN(n9317) );
  AOI22_X1 U9054 ( .A1(ram[4024]), .A2(n8672), .B1(n9325), .B2(n9046), .ZN(
        n8680) );
  INV_X1 U9055 ( .A(n8681), .ZN(n9318) );
  AOI22_X1 U9056 ( .A1(ram[4025]), .A2(n8672), .B1(n9325), .B2(n9070), .ZN(
        n8681) );
  INV_X1 U9057 ( .A(n8682), .ZN(n9319) );
  AOI22_X1 U9058 ( .A1(ram[4026]), .A2(n8672), .B1(n9325), .B2(n9094), .ZN(
        n8682) );
  INV_X1 U9059 ( .A(n8683), .ZN(n9320) );
  AOI22_X1 U9060 ( .A1(ram[4027]), .A2(n8672), .B1(n9325), .B2(n9118), .ZN(
        n8683) );
  INV_X1 U9061 ( .A(n8684), .ZN(n9321) );
  AOI22_X1 U9062 ( .A1(ram[4028]), .A2(n8672), .B1(n9325), .B2(n9142), .ZN(
        n8684) );
  INV_X1 U9063 ( .A(n8685), .ZN(n9322) );
  AOI22_X1 U9064 ( .A1(ram[4029]), .A2(n8672), .B1(n9325), .B2(n9166), .ZN(
        n8685) );
  INV_X1 U9065 ( .A(n8686), .ZN(n9323) );
  AOI22_X1 U9066 ( .A1(ram[4030]), .A2(n8672), .B1(n9325), .B2(n9190), .ZN(
        n8686) );
  INV_X1 U9067 ( .A(n8687), .ZN(n9324) );
  AOI22_X1 U9068 ( .A1(ram[4031]), .A2(n8672), .B1(n9325), .B2(n9214), .ZN(
        n8687) );
  INV_X1 U9069 ( .A(n8706), .ZN(n9275) );
  AOI22_X1 U9070 ( .A1(ram[4048]), .A2(n8707), .B1(n9291), .B2(n8854), .ZN(
        n8706) );
  INV_X1 U9071 ( .A(n8708), .ZN(n9276) );
  AOI22_X1 U9072 ( .A1(ram[4049]), .A2(n8707), .B1(n9291), .B2(n8878), .ZN(
        n8708) );
  INV_X1 U9073 ( .A(n8709), .ZN(n9277) );
  AOI22_X1 U9074 ( .A1(ram[4050]), .A2(n8707), .B1(n9291), .B2(n8902), .ZN(
        n8709) );
  INV_X1 U9075 ( .A(n8710), .ZN(n9278) );
  AOI22_X1 U9076 ( .A1(ram[4051]), .A2(n8707), .B1(n9291), .B2(n8926), .ZN(
        n8710) );
  INV_X1 U9077 ( .A(n8711), .ZN(n9279) );
  AOI22_X1 U9078 ( .A1(ram[4052]), .A2(n8707), .B1(n9291), .B2(n8950), .ZN(
        n8711) );
  INV_X1 U9079 ( .A(n8712), .ZN(n9280) );
  AOI22_X1 U9080 ( .A1(ram[4053]), .A2(n8707), .B1(n9291), .B2(n8974), .ZN(
        n8712) );
  INV_X1 U9081 ( .A(n8713), .ZN(n9281) );
  AOI22_X1 U9082 ( .A1(ram[4054]), .A2(n8707), .B1(n9291), .B2(n8998), .ZN(
        n8713) );
  INV_X1 U9083 ( .A(n8714), .ZN(n9282) );
  AOI22_X1 U9084 ( .A1(ram[4055]), .A2(n8707), .B1(n9291), .B2(n9022), .ZN(
        n8714) );
  INV_X1 U9085 ( .A(n8715), .ZN(n9283) );
  AOI22_X1 U9086 ( .A1(ram[4056]), .A2(n8707), .B1(n9291), .B2(n9046), .ZN(
        n8715) );
  INV_X1 U9087 ( .A(n8716), .ZN(n9284) );
  AOI22_X1 U9088 ( .A1(ram[4057]), .A2(n8707), .B1(n9291), .B2(n9070), .ZN(
        n8716) );
  INV_X1 U9089 ( .A(n8717), .ZN(n9285) );
  AOI22_X1 U9090 ( .A1(ram[4058]), .A2(n8707), .B1(n9291), .B2(n9094), .ZN(
        n8717) );
  INV_X1 U9091 ( .A(n8718), .ZN(n9286) );
  AOI22_X1 U9092 ( .A1(ram[4059]), .A2(n8707), .B1(n9291), .B2(n9118), .ZN(
        n8718) );
  INV_X1 U9093 ( .A(n8719), .ZN(n9287) );
  AOI22_X1 U9094 ( .A1(ram[4060]), .A2(n8707), .B1(n9291), .B2(n9142), .ZN(
        n8719) );
  INV_X1 U9095 ( .A(n8720), .ZN(n9288) );
  AOI22_X1 U9096 ( .A1(ram[4061]), .A2(n8707), .B1(n9291), .B2(n9166), .ZN(
        n8720) );
  INV_X1 U9097 ( .A(n8721), .ZN(n9289) );
  AOI22_X1 U9098 ( .A1(ram[4062]), .A2(n8707), .B1(n9291), .B2(n9190), .ZN(
        n8721) );
  INV_X1 U9099 ( .A(n8722), .ZN(n9290) );
  AOI22_X1 U9100 ( .A1(ram[4063]), .A2(n8707), .B1(n9291), .B2(n9214), .ZN(
        n8722) );
  INV_X1 U9101 ( .A(n8740), .ZN(n9241) );
  AOI22_X1 U9102 ( .A1(ram[4080]), .A2(n8741), .B1(n9257), .B2(n8854), .ZN(
        n8740) );
  INV_X1 U9103 ( .A(n8742), .ZN(n9242) );
  AOI22_X1 U9104 ( .A1(ram[4081]), .A2(n8741), .B1(n9257), .B2(n8878), .ZN(
        n8742) );
  INV_X1 U9105 ( .A(n8743), .ZN(n9243) );
  AOI22_X1 U9106 ( .A1(ram[4082]), .A2(n8741), .B1(n9257), .B2(n8902), .ZN(
        n8743) );
  INV_X1 U9107 ( .A(n8744), .ZN(n9244) );
  AOI22_X1 U9108 ( .A1(ram[4083]), .A2(n8741), .B1(n9257), .B2(n8926), .ZN(
        n8744) );
  INV_X1 U9109 ( .A(n8745), .ZN(n9245) );
  AOI22_X1 U9110 ( .A1(ram[4084]), .A2(n8741), .B1(n9257), .B2(n8950), .ZN(
        n8745) );
  INV_X1 U9111 ( .A(n8746), .ZN(n9246) );
  AOI22_X1 U9112 ( .A1(ram[4085]), .A2(n8741), .B1(n9257), .B2(n8974), .ZN(
        n8746) );
  INV_X1 U9113 ( .A(n8747), .ZN(n9247) );
  AOI22_X1 U9114 ( .A1(ram[4086]), .A2(n8741), .B1(n9257), .B2(n8998), .ZN(
        n8747) );
  INV_X1 U9115 ( .A(n8748), .ZN(n9248) );
  AOI22_X1 U9116 ( .A1(ram[4087]), .A2(n8741), .B1(n9257), .B2(n9022), .ZN(
        n8748) );
  INV_X1 U9117 ( .A(n8749), .ZN(n9249) );
  AOI22_X1 U9118 ( .A1(ram[4088]), .A2(n8741), .B1(n9257), .B2(n9046), .ZN(
        n8749) );
  INV_X1 U9119 ( .A(n8750), .ZN(n9250) );
  AOI22_X1 U9120 ( .A1(ram[4089]), .A2(n8741), .B1(n9257), .B2(n9070), .ZN(
        n8750) );
  INV_X1 U9121 ( .A(n8751), .ZN(n9251) );
  AOI22_X1 U9122 ( .A1(ram[4090]), .A2(n8741), .B1(n9257), .B2(n9094), .ZN(
        n8751) );
  INV_X1 U9123 ( .A(n8752), .ZN(n9252) );
  AOI22_X1 U9124 ( .A1(ram[4091]), .A2(n8741), .B1(n9257), .B2(n9118), .ZN(
        n8752) );
  INV_X1 U9125 ( .A(n8753), .ZN(n9253) );
  AOI22_X1 U9126 ( .A1(ram[4092]), .A2(n8741), .B1(n9257), .B2(n9142), .ZN(
        n8753) );
  INV_X1 U9127 ( .A(n8754), .ZN(n9254) );
  AOI22_X1 U9128 ( .A1(ram[4093]), .A2(n8741), .B1(n9257), .B2(n9166), .ZN(
        n8754) );
  INV_X1 U9129 ( .A(n8755), .ZN(n9255) );
  AOI22_X1 U9130 ( .A1(ram[4094]), .A2(n8741), .B1(n9257), .B2(n9190), .ZN(
        n8755) );
  INV_X1 U9131 ( .A(n8756), .ZN(n9256) );
  AOI22_X1 U9132 ( .A1(ram[4095]), .A2(n8741), .B1(n9257), .B2(n9214), .ZN(
        n8756) );
  AND2_X1 U9133 ( .A1(N300), .A2(mem_read), .ZN(mem_read_data[1]) );
  MUX2_X1 U9134 ( .A(ram[4064]), .B(ram[4080]), .S(n4279), .Z(n1) );
  MUX2_X1 U9135 ( .A(ram[4032]), .B(ram[4048]), .S(n4279), .Z(n2) );
  MUX2_X1 U9136 ( .A(n2), .B(n1), .S(n4174), .Z(n3) );
  MUX2_X1 U9137 ( .A(ram[4000]), .B(ram[4016]), .S(n4279), .Z(n4) );
  MUX2_X1 U9138 ( .A(ram[3968]), .B(ram[3984]), .S(n4279), .Z(n5) );
  MUX2_X1 U9139 ( .A(n5), .B(n4), .S(n4174), .Z(n6) );
  MUX2_X1 U9140 ( .A(n6), .B(n3), .S(n4120), .Z(n7) );
  MUX2_X1 U9141 ( .A(ram[3936]), .B(ram[3952]), .S(n4279), .Z(n8) );
  MUX2_X1 U9142 ( .A(ram[3904]), .B(ram[3920]), .S(n4279), .Z(n9) );
  MUX2_X1 U9143 ( .A(n9), .B(n8), .S(n4174), .Z(n10) );
  MUX2_X1 U9144 ( .A(ram[3872]), .B(ram[3888]), .S(n4279), .Z(n11) );
  MUX2_X1 U9145 ( .A(ram[3840]), .B(ram[3856]), .S(n4279), .Z(n12) );
  MUX2_X1 U9146 ( .A(n12), .B(n11), .S(n4174), .Z(n13) );
  MUX2_X1 U9147 ( .A(n13), .B(n10), .S(n4120), .Z(n14) );
  MUX2_X1 U9148 ( .A(n14), .B(n7), .S(n4087), .Z(n15) );
  MUX2_X1 U9149 ( .A(ram[3808]), .B(ram[3824]), .S(n4280), .Z(n16) );
  MUX2_X1 U9150 ( .A(ram[3776]), .B(ram[3792]), .S(n4280), .Z(n17) );
  MUX2_X1 U9151 ( .A(n17), .B(n16), .S(n4175), .Z(n18) );
  MUX2_X1 U9152 ( .A(ram[3744]), .B(ram[3760]), .S(n4280), .Z(n19) );
  MUX2_X1 U9153 ( .A(ram[3712]), .B(ram[3728]), .S(n4280), .Z(n20010) );
  MUX2_X1 U9154 ( .A(n20010), .B(n19), .S(n4175), .Z(n21010) );
  MUX2_X1 U9155 ( .A(n21010), .B(n18), .S(n4120), .Z(n22010) );
  MUX2_X1 U9156 ( .A(ram[3680]), .B(ram[3696]), .S(n4280), .Z(n23010) );
  MUX2_X1 U9157 ( .A(ram[3648]), .B(ram[3664]), .S(n4280), .Z(n24010) );
  MUX2_X1 U9158 ( .A(n24010), .B(n23010), .S(n4175), .Z(n25010) );
  MUX2_X1 U9159 ( .A(ram[3616]), .B(ram[3632]), .S(n4280), .Z(n26010) );
  MUX2_X1 U9160 ( .A(ram[3584]), .B(ram[3600]), .S(n4280), .Z(n27010) );
  MUX2_X1 U9161 ( .A(n27010), .B(n26010), .S(n4175), .Z(n28) );
  MUX2_X1 U9162 ( .A(n28), .B(n25010), .S(n4120), .Z(n29) );
  MUX2_X1 U9163 ( .A(n29), .B(n22010), .S(n4087), .Z(n30) );
  MUX2_X1 U9164 ( .A(n30), .B(n15), .S(n4076), .Z(n31) );
  MUX2_X1 U9165 ( .A(ram[3552]), .B(ram[3568]), .S(n4280), .Z(n32) );
  MUX2_X1 U9166 ( .A(ram[3520]), .B(ram[3536]), .S(n4280), .Z(n33) );
  MUX2_X1 U9167 ( .A(n33), .B(n32), .S(n4175), .Z(n34) );
  MUX2_X1 U9168 ( .A(ram[3488]), .B(ram[3504]), .S(n4280), .Z(n35) );
  MUX2_X1 U9169 ( .A(ram[3456]), .B(ram[3472]), .S(n4280), .Z(n36) );
  MUX2_X1 U9170 ( .A(n36), .B(n35), .S(n4175), .Z(n37) );
  MUX2_X1 U9171 ( .A(n37), .B(n34), .S(n4120), .Z(n38) );
  MUX2_X1 U9172 ( .A(ram[3424]), .B(ram[3440]), .S(n4281), .Z(n39) );
  MUX2_X1 U9173 ( .A(ram[3392]), .B(ram[3408]), .S(n4281), .Z(n40) );
  MUX2_X1 U9174 ( .A(n40), .B(n39), .S(n4175), .Z(n41) );
  MUX2_X1 U9175 ( .A(ram[3360]), .B(ram[3376]), .S(n4281), .Z(n42) );
  MUX2_X1 U9176 ( .A(ram[3328]), .B(ram[3344]), .S(n4281), .Z(n43) );
  MUX2_X1 U9177 ( .A(n43), .B(n42), .S(n4175), .Z(n44) );
  MUX2_X1 U9178 ( .A(n44), .B(n41), .S(n4120), .Z(n45) );
  MUX2_X1 U9179 ( .A(n45), .B(n38), .S(n4087), .Z(n46) );
  MUX2_X1 U9180 ( .A(ram[3296]), .B(ram[3312]), .S(n4281), .Z(n47) );
  MUX2_X1 U9181 ( .A(ram[3264]), .B(ram[3280]), .S(n4281), .Z(n48) );
  MUX2_X1 U9182 ( .A(n48), .B(n47), .S(n4175), .Z(n49) );
  MUX2_X1 U9183 ( .A(ram[3232]), .B(ram[3248]), .S(n4281), .Z(n50) );
  MUX2_X1 U9184 ( .A(ram[3200]), .B(ram[3216]), .S(n4281), .Z(n51) );
  MUX2_X1 U9185 ( .A(n51), .B(n50), .S(n4175), .Z(n52) );
  MUX2_X1 U9186 ( .A(n52), .B(n49), .S(n4120), .Z(n53) );
  MUX2_X1 U9187 ( .A(ram[3168]), .B(ram[3184]), .S(n4281), .Z(n54) );
  MUX2_X1 U9188 ( .A(ram[3136]), .B(ram[3152]), .S(n4281), .Z(n55) );
  MUX2_X1 U9189 ( .A(n55), .B(n54), .S(n4175), .Z(n56) );
  MUX2_X1 U9190 ( .A(ram[3104]), .B(ram[3120]), .S(n4281), .Z(n57) );
  MUX2_X1 U9191 ( .A(ram[3072]), .B(ram[3088]), .S(n4281), .Z(n58) );
  MUX2_X1 U9192 ( .A(n58), .B(n57), .S(n4175), .Z(n59) );
  MUX2_X1 U9193 ( .A(n59), .B(n56), .S(n4120), .Z(n60) );
  MUX2_X1 U9194 ( .A(n60), .B(n53), .S(n4087), .Z(n61) );
  MUX2_X1 U9195 ( .A(n61), .B(n46), .S(n4076), .Z(n62) );
  MUX2_X1 U9196 ( .A(n62), .B(n31), .S(n4068), .Z(n63) );
  MUX2_X1 U9197 ( .A(ram[3040]), .B(ram[3056]), .S(n4282), .Z(n64) );
  MUX2_X1 U9198 ( .A(ram[3008]), .B(ram[3024]), .S(n4282), .Z(n65) );
  MUX2_X1 U9199 ( .A(n65), .B(n64), .S(n4176), .Z(n66) );
  MUX2_X1 U9200 ( .A(ram[2976]), .B(ram[2992]), .S(n4282), .Z(n67) );
  MUX2_X1 U9201 ( .A(ram[2944]), .B(ram[2960]), .S(n4282), .Z(n68) );
  MUX2_X1 U9202 ( .A(n68), .B(n67), .S(n4176), .Z(n69) );
  MUX2_X1 U9203 ( .A(n69), .B(n66), .S(n4121), .Z(n70) );
  MUX2_X1 U9204 ( .A(ram[2912]), .B(ram[2928]), .S(n4282), .Z(n71) );
  MUX2_X1 U9205 ( .A(ram[2880]), .B(ram[2896]), .S(n4282), .Z(n72) );
  MUX2_X1 U9206 ( .A(n72), .B(n71), .S(n4176), .Z(n73) );
  MUX2_X1 U9207 ( .A(ram[2848]), .B(ram[2864]), .S(n4282), .Z(n74) );
  MUX2_X1 U9208 ( .A(ram[2816]), .B(ram[2832]), .S(n4282), .Z(n75) );
  MUX2_X1 U9209 ( .A(n75), .B(n74), .S(n4176), .Z(n76) );
  MUX2_X1 U9210 ( .A(n76), .B(n73), .S(n4121), .Z(n77) );
  MUX2_X1 U9211 ( .A(n77), .B(n70), .S(n4088), .Z(n78) );
  MUX2_X1 U9212 ( .A(ram[2784]), .B(ram[2800]), .S(n4282), .Z(n79) );
  MUX2_X1 U9213 ( .A(ram[2752]), .B(ram[2768]), .S(n4282), .Z(n80) );
  MUX2_X1 U9214 ( .A(n80), .B(n79), .S(n4176), .Z(n81) );
  MUX2_X1 U9215 ( .A(ram[2720]), .B(ram[2736]), .S(n4282), .Z(n82) );
  MUX2_X1 U9216 ( .A(ram[2688]), .B(ram[2704]), .S(n4282), .Z(n83) );
  MUX2_X1 U9217 ( .A(n83), .B(n82), .S(n4176), .Z(n84) );
  MUX2_X1 U9218 ( .A(n84), .B(n81), .S(n4121), .Z(n85) );
  MUX2_X1 U9219 ( .A(ram[2656]), .B(ram[2672]), .S(n4283), .Z(n86) );
  MUX2_X1 U9220 ( .A(ram[2624]), .B(ram[2640]), .S(n4283), .Z(n87) );
  MUX2_X1 U9221 ( .A(n87), .B(n86), .S(n4176), .Z(n88) );
  MUX2_X1 U9222 ( .A(ram[2592]), .B(ram[2608]), .S(n4283), .Z(n89) );
  MUX2_X1 U9223 ( .A(ram[2560]), .B(ram[2576]), .S(n4283), .Z(n90) );
  MUX2_X1 U9224 ( .A(n90), .B(n89), .S(n4176), .Z(n91) );
  MUX2_X1 U9225 ( .A(n91), .B(n88), .S(n4121), .Z(n92) );
  MUX2_X1 U9226 ( .A(n92), .B(n85), .S(n4088), .Z(n93) );
  MUX2_X1 U9227 ( .A(n93), .B(n78), .S(n4076), .Z(n94) );
  MUX2_X1 U9228 ( .A(ram[2528]), .B(ram[2544]), .S(n4283), .Z(n95) );
  MUX2_X1 U9229 ( .A(ram[2496]), .B(ram[2512]), .S(n4283), .Z(n96) );
  MUX2_X1 U9230 ( .A(n96), .B(n95), .S(n4176), .Z(n97) );
  MUX2_X1 U9231 ( .A(ram[2464]), .B(ram[2480]), .S(n4283), .Z(n98) );
  MUX2_X1 U9232 ( .A(ram[2432]), .B(ram[2448]), .S(n4283), .Z(n99) );
  MUX2_X1 U9233 ( .A(n99), .B(n98), .S(n4176), .Z(n100) );
  MUX2_X1 U9234 ( .A(n100), .B(n97), .S(n4121), .Z(n101) );
  MUX2_X1 U9235 ( .A(ram[2400]), .B(ram[2416]), .S(n4283), .Z(n102) );
  MUX2_X1 U9236 ( .A(ram[2368]), .B(ram[2384]), .S(n4283), .Z(n103) );
  MUX2_X1 U9237 ( .A(n103), .B(n102), .S(n4176), .Z(n104) );
  MUX2_X1 U9238 ( .A(ram[2336]), .B(ram[2352]), .S(n4283), .Z(n105) );
  MUX2_X1 U9239 ( .A(ram[2304]), .B(ram[2320]), .S(n4283), .Z(n106) );
  MUX2_X1 U9240 ( .A(n106), .B(n105), .S(n4176), .Z(n107) );
  MUX2_X1 U9241 ( .A(n107), .B(n104), .S(n4121), .Z(n108) );
  MUX2_X1 U9242 ( .A(n108), .B(n101), .S(n4088), .Z(n109) );
  MUX2_X1 U9243 ( .A(ram[2272]), .B(ram[2288]), .S(n4284), .Z(n110) );
  MUX2_X1 U9244 ( .A(ram[2240]), .B(ram[2256]), .S(n4284), .Z(n111) );
  MUX2_X1 U9245 ( .A(n111), .B(n110), .S(n4177), .Z(n112) );
  MUX2_X1 U9246 ( .A(ram[2208]), .B(ram[2224]), .S(n4284), .Z(n113) );
  MUX2_X1 U9247 ( .A(ram[2176]), .B(ram[2192]), .S(n4284), .Z(n114) );
  MUX2_X1 U9248 ( .A(n114), .B(n113), .S(n4177), .Z(n115) );
  MUX2_X1 U9249 ( .A(n115), .B(n112), .S(n4121), .Z(n116) );
  MUX2_X1 U9250 ( .A(ram[2144]), .B(ram[2160]), .S(n4284), .Z(n117) );
  MUX2_X1 U9251 ( .A(ram[2112]), .B(ram[2128]), .S(n4284), .Z(n118) );
  MUX2_X1 U9252 ( .A(n118), .B(n117), .S(n4177), .Z(n119) );
  MUX2_X1 U9253 ( .A(ram[2080]), .B(ram[2096]), .S(n4284), .Z(n120) );
  MUX2_X1 U9254 ( .A(ram[2048]), .B(ram[2064]), .S(n4284), .Z(n121) );
  MUX2_X1 U9255 ( .A(n121), .B(n120), .S(n4177), .Z(n122) );
  MUX2_X1 U9256 ( .A(n122), .B(n119), .S(n4121), .Z(n123) );
  MUX2_X1 U9257 ( .A(n123), .B(n116), .S(n4088), .Z(n124) );
  MUX2_X1 U9258 ( .A(n124), .B(n109), .S(n4076), .Z(n125) );
  MUX2_X1 U9259 ( .A(n125), .B(n94), .S(n4068), .Z(n126) );
  MUX2_X1 U9260 ( .A(n126), .B(n63), .S(n4065), .Z(n127) );
  MUX2_X1 U9261 ( .A(ram[2016]), .B(ram[2032]), .S(n4284), .Z(n128) );
  MUX2_X1 U9262 ( .A(ram[1984]), .B(ram[2000]), .S(n4284), .Z(n129) );
  MUX2_X1 U9263 ( .A(n129), .B(n128), .S(n4177), .Z(n130) );
  MUX2_X1 U9264 ( .A(ram[1952]), .B(ram[1968]), .S(n4284), .Z(n131) );
  MUX2_X1 U9265 ( .A(ram[1920]), .B(ram[1936]), .S(n4284), .Z(n132) );
  MUX2_X1 U9266 ( .A(n132), .B(n131), .S(n4177), .Z(n133) );
  MUX2_X1 U9267 ( .A(n133), .B(n130), .S(n4121), .Z(n134) );
  MUX2_X1 U9268 ( .A(ram[1888]), .B(ram[1904]), .S(n4285), .Z(n135) );
  MUX2_X1 U9269 ( .A(ram[1856]), .B(ram[1872]), .S(n4285), .Z(n136) );
  MUX2_X1 U9270 ( .A(n136), .B(n135), .S(n4177), .Z(n137) );
  MUX2_X1 U9271 ( .A(ram[1824]), .B(ram[1840]), .S(n4285), .Z(n138) );
  MUX2_X1 U9272 ( .A(ram[1792]), .B(ram[1808]), .S(n4285), .Z(n139) );
  MUX2_X1 U9273 ( .A(n139), .B(n138), .S(n4177), .Z(n140) );
  MUX2_X1 U9274 ( .A(n140), .B(n137), .S(n4121), .Z(n141) );
  MUX2_X1 U9275 ( .A(n141), .B(n134), .S(n4088), .Z(n142) );
  MUX2_X1 U9276 ( .A(ram[1760]), .B(ram[1776]), .S(n4285), .Z(n143) );
  MUX2_X1 U9277 ( .A(ram[1728]), .B(ram[1744]), .S(n4285), .Z(n144) );
  MUX2_X1 U9278 ( .A(n144), .B(n143), .S(n4177), .Z(n145) );
  MUX2_X1 U9279 ( .A(ram[1696]), .B(ram[1712]), .S(n4285), .Z(n146) );
  MUX2_X1 U9280 ( .A(ram[1664]), .B(ram[1680]), .S(n4285), .Z(n147) );
  MUX2_X1 U9281 ( .A(n147), .B(n146), .S(n4177), .Z(n148) );
  MUX2_X1 U9282 ( .A(n148), .B(n145), .S(n4121), .Z(n149) );
  MUX2_X1 U9283 ( .A(ram[1632]), .B(ram[1648]), .S(n4285), .Z(n150) );
  MUX2_X1 U9284 ( .A(ram[1600]), .B(ram[1616]), .S(n4285), .Z(n151) );
  MUX2_X1 U9285 ( .A(n151), .B(n150), .S(n4177), .Z(n152) );
  MUX2_X1 U9286 ( .A(ram[1568]), .B(ram[1584]), .S(n4285), .Z(n153) );
  MUX2_X1 U9287 ( .A(ram[1536]), .B(ram[1552]), .S(n4285), .Z(n154) );
  MUX2_X1 U9288 ( .A(n154), .B(n153), .S(n4177), .Z(n155) );
  MUX2_X1 U9289 ( .A(n155), .B(n152), .S(n4121), .Z(n156) );
  MUX2_X1 U9290 ( .A(n156), .B(n149), .S(n4088), .Z(n157) );
  MUX2_X1 U9291 ( .A(n157), .B(n142), .S(n4076), .Z(n158) );
  MUX2_X1 U9292 ( .A(ram[1504]), .B(ram[1520]), .S(n4286), .Z(n159) );
  MUX2_X1 U9293 ( .A(ram[1472]), .B(ram[1488]), .S(n4286), .Z(n160) );
  MUX2_X1 U9294 ( .A(n160), .B(n159), .S(n4178), .Z(n161) );
  MUX2_X1 U9295 ( .A(ram[1440]), .B(ram[1456]), .S(n4286), .Z(n162) );
  MUX2_X1 U9296 ( .A(ram[1408]), .B(ram[1424]), .S(n4286), .Z(n163) );
  MUX2_X1 U9297 ( .A(n163), .B(n162), .S(n4178), .Z(n164) );
  MUX2_X1 U9298 ( .A(n164), .B(n161), .S(n4122), .Z(n165) );
  MUX2_X1 U9299 ( .A(ram[1376]), .B(ram[1392]), .S(n4286), .Z(n166) );
  MUX2_X1 U9300 ( .A(ram[1344]), .B(ram[1360]), .S(n4286), .Z(n167) );
  MUX2_X1 U9301 ( .A(n167), .B(n166), .S(n4178), .Z(n168) );
  MUX2_X1 U9302 ( .A(ram[1312]), .B(ram[1328]), .S(n4286), .Z(n169) );
  MUX2_X1 U9303 ( .A(ram[1280]), .B(ram[1296]), .S(n4286), .Z(n170) );
  MUX2_X1 U9304 ( .A(n170), .B(n169), .S(n4178), .Z(n171) );
  MUX2_X1 U9305 ( .A(n171), .B(n168), .S(n4122), .Z(n172) );
  MUX2_X1 U9306 ( .A(n172), .B(n165), .S(n4088), .Z(n173) );
  MUX2_X1 U9307 ( .A(ram[1248]), .B(ram[1264]), .S(n4286), .Z(n174) );
  MUX2_X1 U9308 ( .A(ram[1216]), .B(ram[1232]), .S(n4286), .Z(n175) );
  MUX2_X1 U9309 ( .A(n175), .B(n174), .S(n4178), .Z(n176) );
  MUX2_X1 U9310 ( .A(ram[1184]), .B(ram[1200]), .S(n4286), .Z(n177) );
  MUX2_X1 U9311 ( .A(ram[1152]), .B(ram[1168]), .S(n4286), .Z(n178) );
  MUX2_X1 U9312 ( .A(n178), .B(n177), .S(n4178), .Z(n179) );
  MUX2_X1 U9313 ( .A(n179), .B(n176), .S(n4122), .Z(n180) );
  MUX2_X1 U9314 ( .A(ram[1120]), .B(ram[1136]), .S(n4287), .Z(n181) );
  MUX2_X1 U9315 ( .A(ram[1088]), .B(ram[1104]), .S(n4287), .Z(n182) );
  MUX2_X1 U9316 ( .A(n182), .B(n181), .S(n4178), .Z(n183) );
  MUX2_X1 U9317 ( .A(ram[1056]), .B(ram[1072]), .S(n4287), .Z(n184) );
  MUX2_X1 U9318 ( .A(ram[1024]), .B(ram[1040]), .S(n4287), .Z(n185) );
  MUX2_X1 U9319 ( .A(n185), .B(n184), .S(n4178), .Z(n186) );
  MUX2_X1 U9320 ( .A(n186), .B(n183), .S(n4122), .Z(n187) );
  MUX2_X1 U9321 ( .A(n187), .B(n180), .S(n4088), .Z(n188) );
  MUX2_X1 U9322 ( .A(n188), .B(n173), .S(n4076), .Z(n189) );
  MUX2_X1 U9323 ( .A(n189), .B(n158), .S(n4068), .Z(n190) );
  MUX2_X1 U9324 ( .A(ram[992]), .B(ram[1008]), .S(n4287), .Z(n191) );
  MUX2_X1 U9325 ( .A(ram[960]), .B(ram[976]), .S(n4287), .Z(n192) );
  MUX2_X1 U9326 ( .A(n192), .B(n191), .S(n4178), .Z(n193) );
  MUX2_X1 U9327 ( .A(ram[928]), .B(ram[944]), .S(n4287), .Z(n194) );
  MUX2_X1 U9328 ( .A(ram[896]), .B(ram[912]), .S(n4287), .Z(n195) );
  MUX2_X1 U9329 ( .A(n195), .B(n194), .S(n4178), .Z(n196) );
  MUX2_X1 U9330 ( .A(n196), .B(n193), .S(n4122), .Z(n197) );
  MUX2_X1 U9331 ( .A(ram[864]), .B(ram[880]), .S(n4287), .Z(n198) );
  MUX2_X1 U9332 ( .A(ram[832]), .B(ram[848]), .S(n4287), .Z(n199) );
  MUX2_X1 U9333 ( .A(n199), .B(n198), .S(n4178), .Z(n20000) );
  MUX2_X1 U9334 ( .A(ram[800]), .B(ram[816]), .S(n4287), .Z(n201) );
  MUX2_X1 U9335 ( .A(ram[768]), .B(ram[784]), .S(n4287), .Z(n202) );
  MUX2_X1 U9336 ( .A(n202), .B(n201), .S(n4178), .Z(n203) );
  MUX2_X1 U9337 ( .A(n203), .B(n20000), .S(n4122), .Z(n204) );
  MUX2_X1 U9338 ( .A(n204), .B(n197), .S(n4088), .Z(n205) );
  MUX2_X1 U9339 ( .A(ram[736]), .B(ram[752]), .S(n4288), .Z(n206) );
  MUX2_X1 U9340 ( .A(ram[704]), .B(ram[720]), .S(n4288), .Z(n207) );
  MUX2_X1 U9341 ( .A(n207), .B(n206), .S(n4179), .Z(n208) );
  MUX2_X1 U9342 ( .A(ram[672]), .B(ram[688]), .S(n4288), .Z(n209) );
  MUX2_X1 U9343 ( .A(ram[640]), .B(ram[656]), .S(n4288), .Z(n21000) );
  MUX2_X1 U9344 ( .A(n21000), .B(n209), .S(n4179), .Z(n211) );
  MUX2_X1 U9345 ( .A(n211), .B(n208), .S(n4122), .Z(n212) );
  MUX2_X1 U9346 ( .A(ram[608]), .B(ram[624]), .S(n4288), .Z(n213) );
  MUX2_X1 U9347 ( .A(ram[576]), .B(ram[592]), .S(n4288), .Z(n214) );
  MUX2_X1 U9348 ( .A(n214), .B(n213), .S(n4179), .Z(n215) );
  MUX2_X1 U9349 ( .A(ram[544]), .B(ram[560]), .S(n4288), .Z(n216) );
  MUX2_X1 U9350 ( .A(ram[512]), .B(ram[528]), .S(n4288), .Z(n217) );
  MUX2_X1 U9351 ( .A(n217), .B(n216), .S(n4179), .Z(n218) );
  MUX2_X1 U9352 ( .A(n218), .B(n215), .S(n4122), .Z(n219) );
  MUX2_X1 U9353 ( .A(n219), .B(n212), .S(n4088), .Z(n22000) );
  MUX2_X1 U9354 ( .A(n22000), .B(n205), .S(n4076), .Z(n221) );
  MUX2_X1 U9355 ( .A(ram[480]), .B(ram[496]), .S(n4288), .Z(n222) );
  MUX2_X1 U9356 ( .A(ram[448]), .B(ram[464]), .S(n4288), .Z(n223) );
  MUX2_X1 U9357 ( .A(n223), .B(n222), .S(n4179), .Z(n224) );
  MUX2_X1 U9358 ( .A(ram[416]), .B(ram[432]), .S(n4288), .Z(n225) );
  MUX2_X1 U9359 ( .A(ram[384]), .B(ram[400]), .S(n4288), .Z(n226) );
  MUX2_X1 U9360 ( .A(n226), .B(n225), .S(n4179), .Z(n227) );
  MUX2_X1 U9361 ( .A(n227), .B(n224), .S(n4122), .Z(n228) );
  MUX2_X1 U9362 ( .A(ram[352]), .B(ram[368]), .S(n4289), .Z(n229) );
  MUX2_X1 U9363 ( .A(ram[320]), .B(ram[336]), .S(n4289), .Z(n23000) );
  MUX2_X1 U9364 ( .A(n23000), .B(n229), .S(n4179), .Z(n231) );
  MUX2_X1 U9365 ( .A(ram[288]), .B(ram[304]), .S(n4289), .Z(n232) );
  MUX2_X1 U9366 ( .A(ram[256]), .B(ram[272]), .S(n4289), .Z(n233) );
  MUX2_X1 U9367 ( .A(n233), .B(n232), .S(n4179), .Z(n234) );
  MUX2_X1 U9368 ( .A(n234), .B(n231), .S(n4122), .Z(n235) );
  MUX2_X1 U9369 ( .A(n235), .B(n228), .S(n4088), .Z(n236) );
  MUX2_X1 U9370 ( .A(ram[224]), .B(ram[240]), .S(n4289), .Z(n237) );
  MUX2_X1 U9371 ( .A(ram[192]), .B(ram[208]), .S(n4289), .Z(n238) );
  MUX2_X1 U9372 ( .A(n238), .B(n237), .S(n4179), .Z(n239) );
  MUX2_X1 U9373 ( .A(ram[160]), .B(ram[176]), .S(n4289), .Z(n24000) );
  MUX2_X1 U9374 ( .A(ram[128]), .B(ram[144]), .S(n4289), .Z(n241) );
  MUX2_X1 U9375 ( .A(n241), .B(n24000), .S(n4179), .Z(n242) );
  MUX2_X1 U9376 ( .A(n242), .B(n239), .S(n4122), .Z(n243) );
  MUX2_X1 U9377 ( .A(ram[96]), .B(ram[112]), .S(n4289), .Z(n244) );
  MUX2_X1 U9378 ( .A(ram[64]), .B(ram[80]), .S(n4289), .Z(n245) );
  MUX2_X1 U9379 ( .A(n245), .B(n244), .S(n4179), .Z(n246) );
  MUX2_X1 U9380 ( .A(ram[32]), .B(ram[48]), .S(n4289), .Z(n247) );
  MUX2_X1 U9381 ( .A(ram[0]), .B(ram[16]), .S(n4289), .Z(n248) );
  MUX2_X1 U9382 ( .A(n248), .B(n247), .S(n4179), .Z(n249) );
  MUX2_X1 U9383 ( .A(n249), .B(n246), .S(n4122), .Z(n25000) );
  MUX2_X1 U9384 ( .A(n25000), .B(n243), .S(n4088), .Z(n251) );
  MUX2_X1 U9385 ( .A(n251), .B(n236), .S(n4076), .Z(n252) );
  MUX2_X1 U9386 ( .A(n252), .B(n221), .S(n4068), .Z(n253) );
  MUX2_X1 U9387 ( .A(n253), .B(n190), .S(n4065), .Z(n254) );
  MUX2_X1 U9388 ( .A(n254), .B(n127), .S(mem_access_addr[9]), .Z(N301) );
  MUX2_X1 U9389 ( .A(ram[4065]), .B(ram[4081]), .S(n4290), .Z(n255) );
  MUX2_X1 U9390 ( .A(ram[4033]), .B(ram[4049]), .S(n4290), .Z(n256) );
  MUX2_X1 U9391 ( .A(n256), .B(n255), .S(n4180), .Z(n257) );
  MUX2_X1 U9392 ( .A(ram[4001]), .B(ram[4017]), .S(n4290), .Z(n258) );
  MUX2_X1 U9393 ( .A(ram[3969]), .B(ram[3985]), .S(n4290), .Z(n259) );
  MUX2_X1 U9394 ( .A(n259), .B(n258), .S(n4180), .Z(n26000) );
  MUX2_X1 U9395 ( .A(n26000), .B(n257), .S(n4123), .Z(n261) );
  MUX2_X1 U9396 ( .A(ram[3937]), .B(ram[3953]), .S(n4290), .Z(n262) );
  MUX2_X1 U9397 ( .A(ram[3905]), .B(ram[3921]), .S(n4290), .Z(n263) );
  MUX2_X1 U9398 ( .A(n263), .B(n262), .S(n4180), .Z(n264) );
  MUX2_X1 U9399 ( .A(ram[3873]), .B(ram[3889]), .S(n4290), .Z(n265) );
  MUX2_X1 U9400 ( .A(ram[3841]), .B(ram[3857]), .S(n4290), .Z(n266) );
  MUX2_X1 U9401 ( .A(n266), .B(n265), .S(n4180), .Z(n267) );
  MUX2_X1 U9402 ( .A(n267), .B(n264), .S(n4123), .Z(n268) );
  MUX2_X1 U9403 ( .A(n268), .B(n261), .S(n4089), .Z(n269) );
  MUX2_X1 U9404 ( .A(ram[3809]), .B(ram[3825]), .S(n4290), .Z(n27000) );
  MUX2_X1 U9405 ( .A(ram[3777]), .B(ram[3793]), .S(n4290), .Z(n271) );
  MUX2_X1 U9406 ( .A(n271), .B(n27000), .S(n4180), .Z(n272) );
  MUX2_X1 U9407 ( .A(ram[3745]), .B(ram[3761]), .S(n4290), .Z(n273) );
  MUX2_X1 U9408 ( .A(ram[3713]), .B(ram[3729]), .S(n4290), .Z(n274) );
  MUX2_X1 U9409 ( .A(n274), .B(n273), .S(n4180), .Z(n275) );
  MUX2_X1 U9410 ( .A(n275), .B(n272), .S(n4123), .Z(n276) );
  MUX2_X1 U9411 ( .A(ram[3681]), .B(ram[3697]), .S(n4291), .Z(n277) );
  MUX2_X1 U9412 ( .A(ram[3649]), .B(ram[3665]), .S(n4291), .Z(n278) );
  MUX2_X1 U9413 ( .A(n278), .B(n277), .S(n4180), .Z(n279) );
  MUX2_X1 U9414 ( .A(ram[3617]), .B(ram[3633]), .S(n4291), .Z(n280) );
  MUX2_X1 U9415 ( .A(ram[3585]), .B(ram[3601]), .S(n4291), .Z(n281) );
  MUX2_X1 U9416 ( .A(n281), .B(n280), .S(n4180), .Z(n282) );
  MUX2_X1 U9417 ( .A(n282), .B(n279), .S(n4123), .Z(n283) );
  MUX2_X1 U9418 ( .A(n283), .B(n276), .S(n4089), .Z(n284) );
  MUX2_X1 U9419 ( .A(n284), .B(n269), .S(n4077), .Z(n285) );
  MUX2_X1 U9420 ( .A(ram[3553]), .B(ram[3569]), .S(n4291), .Z(n28600) );
  MUX2_X1 U9421 ( .A(ram[3521]), .B(ram[3537]), .S(n4291), .Z(n28700) );
  MUX2_X1 U9422 ( .A(n28700), .B(n28600), .S(n4180), .Z(n28800) );
  MUX2_X1 U9423 ( .A(ram[3489]), .B(ram[3505]), .S(n4291), .Z(n28900) );
  MUX2_X1 U9424 ( .A(ram[3457]), .B(ram[3473]), .S(n4291), .Z(n29000) );
  MUX2_X1 U9425 ( .A(n29000), .B(n28900), .S(n4180), .Z(n29100) );
  MUX2_X1 U9426 ( .A(n29100), .B(n28800), .S(n4123), .Z(n29200) );
  MUX2_X1 U9427 ( .A(ram[3425]), .B(ram[3441]), .S(n4291), .Z(n29300) );
  MUX2_X1 U9428 ( .A(ram[3393]), .B(ram[3409]), .S(n4291), .Z(n29400) );
  MUX2_X1 U9429 ( .A(n29400), .B(n29300), .S(n4180), .Z(n29500) );
  MUX2_X1 U9430 ( .A(ram[3361]), .B(ram[3377]), .S(n4291), .Z(n29600) );
  MUX2_X1 U9431 ( .A(ram[3329]), .B(ram[3345]), .S(n4291), .Z(n29700) );
  MUX2_X1 U9432 ( .A(n29700), .B(n29600), .S(n4180), .Z(n29800) );
  MUX2_X1 U9433 ( .A(n29800), .B(n29500), .S(n4123), .Z(n29900) );
  MUX2_X1 U9434 ( .A(n29900), .B(n29200), .S(n4089), .Z(n30000) );
  MUX2_X1 U9435 ( .A(ram[3297]), .B(ram[3313]), .S(n4292), .Z(n30100) );
  MUX2_X1 U9436 ( .A(ram[3265]), .B(ram[3281]), .S(n4292), .Z(n302) );
  MUX2_X1 U9437 ( .A(n302), .B(n30100), .S(n4181), .Z(n303) );
  MUX2_X1 U9438 ( .A(ram[3233]), .B(ram[3249]), .S(n4292), .Z(n304) );
  MUX2_X1 U9439 ( .A(ram[3201]), .B(ram[3217]), .S(n4292), .Z(n305) );
  MUX2_X1 U9440 ( .A(n305), .B(n304), .S(n4181), .Z(n306) );
  MUX2_X1 U9441 ( .A(n306), .B(n303), .S(n4123), .Z(n307) );
  MUX2_X1 U9442 ( .A(ram[3169]), .B(ram[3185]), .S(n4292), .Z(n308) );
  MUX2_X1 U9443 ( .A(ram[3137]), .B(ram[3153]), .S(n4292), .Z(n309) );
  MUX2_X1 U9444 ( .A(n309), .B(n308), .S(n4181), .Z(n310) );
  MUX2_X1 U9445 ( .A(ram[3105]), .B(ram[3121]), .S(n4292), .Z(n311) );
  MUX2_X1 U9446 ( .A(ram[3073]), .B(ram[3089]), .S(n4292), .Z(n312) );
  MUX2_X1 U9447 ( .A(n312), .B(n311), .S(n4181), .Z(n313) );
  MUX2_X1 U9448 ( .A(n313), .B(n310), .S(n4123), .Z(n314) );
  MUX2_X1 U9449 ( .A(n314), .B(n307), .S(n4089), .Z(n315) );
  MUX2_X1 U9450 ( .A(n315), .B(n30000), .S(n4077), .Z(n316) );
  MUX2_X1 U9451 ( .A(n316), .B(n285), .S(n4069), .Z(n317) );
  MUX2_X1 U9452 ( .A(ram[3041]), .B(ram[3057]), .S(n4292), .Z(n318) );
  MUX2_X1 U9453 ( .A(ram[3009]), .B(ram[3025]), .S(n4292), .Z(n319) );
  MUX2_X1 U9454 ( .A(n319), .B(n318), .S(n4181), .Z(n320) );
  MUX2_X1 U9455 ( .A(ram[2977]), .B(ram[2993]), .S(n4292), .Z(n321) );
  MUX2_X1 U9456 ( .A(ram[2945]), .B(ram[2961]), .S(n4292), .Z(n322) );
  MUX2_X1 U9457 ( .A(n322), .B(n321), .S(n4181), .Z(n323) );
  MUX2_X1 U9458 ( .A(n323), .B(n320), .S(n4123), .Z(n324) );
  MUX2_X1 U9459 ( .A(ram[2913]), .B(ram[2929]), .S(n4293), .Z(n325) );
  MUX2_X1 U9460 ( .A(ram[2881]), .B(ram[2897]), .S(n4293), .Z(n326) );
  MUX2_X1 U9461 ( .A(n326), .B(n325), .S(n4181), .Z(n327) );
  MUX2_X1 U9462 ( .A(ram[2849]), .B(ram[2865]), .S(n4293), .Z(n328) );
  MUX2_X1 U9463 ( .A(ram[2817]), .B(ram[2833]), .S(n4293), .Z(n329) );
  MUX2_X1 U9464 ( .A(n329), .B(n328), .S(n4181), .Z(n330) );
  MUX2_X1 U9465 ( .A(n330), .B(n327), .S(n4123), .Z(n331) );
  MUX2_X1 U9466 ( .A(n331), .B(n324), .S(n4089), .Z(n332) );
  MUX2_X1 U9467 ( .A(ram[2785]), .B(ram[2801]), .S(n4293), .Z(n333) );
  MUX2_X1 U9468 ( .A(ram[2753]), .B(ram[2769]), .S(n4293), .Z(n334) );
  MUX2_X1 U9469 ( .A(n334), .B(n333), .S(n4181), .Z(n335) );
  MUX2_X1 U9470 ( .A(ram[2721]), .B(ram[2737]), .S(n4293), .Z(n336) );
  MUX2_X1 U9471 ( .A(ram[2689]), .B(ram[2705]), .S(n4293), .Z(n337) );
  MUX2_X1 U9472 ( .A(n337), .B(n336), .S(n4181), .Z(n338) );
  MUX2_X1 U9473 ( .A(n338), .B(n335), .S(n4123), .Z(n339) );
  MUX2_X1 U9474 ( .A(ram[2657]), .B(ram[2673]), .S(n4293), .Z(n340) );
  MUX2_X1 U9475 ( .A(ram[2625]), .B(ram[2641]), .S(n4293), .Z(n341) );
  MUX2_X1 U9476 ( .A(n341), .B(n340), .S(n4181), .Z(n342) );
  MUX2_X1 U9477 ( .A(ram[2593]), .B(ram[2609]), .S(n4293), .Z(n343) );
  MUX2_X1 U9478 ( .A(ram[2561]), .B(ram[2577]), .S(n4293), .Z(n344) );
  MUX2_X1 U9479 ( .A(n344), .B(n343), .S(n4181), .Z(n345) );
  MUX2_X1 U9480 ( .A(n345), .B(n342), .S(n4123), .Z(n346) );
  MUX2_X1 U9481 ( .A(n346), .B(n339), .S(n4089), .Z(n347) );
  MUX2_X1 U9482 ( .A(n347), .B(n332), .S(n4077), .Z(n348) );
  MUX2_X1 U9483 ( .A(ram[2529]), .B(ram[2545]), .S(n4294), .Z(n349) );
  MUX2_X1 U9484 ( .A(ram[2497]), .B(ram[2513]), .S(n4294), .Z(n350) );
  MUX2_X1 U9485 ( .A(n350), .B(n349), .S(n4182), .Z(n351) );
  MUX2_X1 U9486 ( .A(ram[2465]), .B(ram[2481]), .S(n4294), .Z(n352) );
  MUX2_X1 U9487 ( .A(ram[2433]), .B(ram[2449]), .S(n4294), .Z(n353) );
  MUX2_X1 U9488 ( .A(n353), .B(n352), .S(n4182), .Z(n354) );
  MUX2_X1 U9489 ( .A(n354), .B(n351), .S(n4124), .Z(n355) );
  MUX2_X1 U9490 ( .A(ram[2401]), .B(ram[2417]), .S(n4294), .Z(n356) );
  MUX2_X1 U9491 ( .A(ram[2369]), .B(ram[2385]), .S(n4294), .Z(n357) );
  MUX2_X1 U9492 ( .A(n357), .B(n356), .S(n4182), .Z(n358) );
  MUX2_X1 U9493 ( .A(ram[2337]), .B(ram[2353]), .S(n4294), .Z(n359) );
  MUX2_X1 U9494 ( .A(ram[2305]), .B(ram[2321]), .S(n4294), .Z(n360) );
  MUX2_X1 U9495 ( .A(n360), .B(n359), .S(n4182), .Z(n361) );
  MUX2_X1 U9496 ( .A(n361), .B(n358), .S(n4124), .Z(n362) );
  MUX2_X1 U9497 ( .A(n362), .B(n355), .S(n4089), .Z(n363) );
  MUX2_X1 U9498 ( .A(ram[2273]), .B(ram[2289]), .S(n4294), .Z(n364) );
  MUX2_X1 U9499 ( .A(ram[2241]), .B(ram[2257]), .S(n4294), .Z(n365) );
  MUX2_X1 U9500 ( .A(n365), .B(n364), .S(n4182), .Z(n366) );
  MUX2_X1 U9501 ( .A(ram[2209]), .B(ram[2225]), .S(n4294), .Z(n367) );
  MUX2_X1 U9502 ( .A(ram[2177]), .B(ram[2193]), .S(n4294), .Z(n368) );
  MUX2_X1 U9503 ( .A(n368), .B(n367), .S(n4182), .Z(n369) );
  MUX2_X1 U9504 ( .A(n369), .B(n366), .S(n4124), .Z(n370) );
  MUX2_X1 U9505 ( .A(ram[2145]), .B(ram[2161]), .S(n4295), .Z(n371) );
  MUX2_X1 U9506 ( .A(ram[2113]), .B(ram[2129]), .S(n4295), .Z(n372) );
  MUX2_X1 U9507 ( .A(n372), .B(n371), .S(n4182), .Z(n373) );
  MUX2_X1 U9508 ( .A(ram[2081]), .B(ram[2097]), .S(n4295), .Z(n374) );
  MUX2_X1 U9509 ( .A(ram[2049]), .B(ram[2065]), .S(n4295), .Z(n375) );
  MUX2_X1 U9510 ( .A(n375), .B(n374), .S(n4182), .Z(n376) );
  MUX2_X1 U9511 ( .A(n376), .B(n373), .S(n4124), .Z(n377) );
  MUX2_X1 U9512 ( .A(n377), .B(n370), .S(n4089), .Z(n378) );
  MUX2_X1 U9513 ( .A(n378), .B(n363), .S(n4077), .Z(n379) );
  MUX2_X1 U9514 ( .A(n379), .B(n348), .S(n4069), .Z(n380) );
  MUX2_X1 U9515 ( .A(n380), .B(n317), .S(n4065), .Z(n381) );
  MUX2_X1 U9516 ( .A(ram[2017]), .B(ram[2033]), .S(n4295), .Z(n382) );
  MUX2_X1 U9517 ( .A(ram[1985]), .B(ram[2001]), .S(n4295), .Z(n383) );
  MUX2_X1 U9518 ( .A(n383), .B(n382), .S(n4182), .Z(n384) );
  MUX2_X1 U9519 ( .A(ram[1953]), .B(ram[1969]), .S(n4295), .Z(n385) );
  MUX2_X1 U9520 ( .A(ram[1921]), .B(ram[1937]), .S(n4295), .Z(n386) );
  MUX2_X1 U9521 ( .A(n386), .B(n385), .S(n4182), .Z(n387) );
  MUX2_X1 U9522 ( .A(n387), .B(n384), .S(n4124), .Z(n388) );
  MUX2_X1 U9523 ( .A(ram[1889]), .B(ram[1905]), .S(n4295), .Z(n389) );
  MUX2_X1 U9524 ( .A(ram[1857]), .B(ram[1873]), .S(n4295), .Z(n390) );
  MUX2_X1 U9525 ( .A(n390), .B(n389), .S(n4182), .Z(n391) );
  MUX2_X1 U9526 ( .A(ram[1825]), .B(ram[1841]), .S(n4295), .Z(n392) );
  MUX2_X1 U9527 ( .A(ram[1793]), .B(ram[1809]), .S(n4295), .Z(n393) );
  MUX2_X1 U9528 ( .A(n393), .B(n392), .S(n4182), .Z(n394) );
  MUX2_X1 U9529 ( .A(n394), .B(n391), .S(n4124), .Z(n395) );
  MUX2_X1 U9530 ( .A(n395), .B(n388), .S(n4089), .Z(n396) );
  MUX2_X1 U9531 ( .A(ram[1761]), .B(ram[1777]), .S(n4296), .Z(n397) );
  MUX2_X1 U9532 ( .A(ram[1729]), .B(ram[1745]), .S(n4296), .Z(n398) );
  MUX2_X1 U9533 ( .A(n398), .B(n397), .S(n4183), .Z(n399) );
  MUX2_X1 U9534 ( .A(ram[1697]), .B(ram[1713]), .S(n4296), .Z(n400) );
  MUX2_X1 U9535 ( .A(ram[1665]), .B(ram[1681]), .S(n4296), .Z(n401) );
  MUX2_X1 U9536 ( .A(n401), .B(n400), .S(n4183), .Z(n402) );
  MUX2_X1 U9537 ( .A(n402), .B(n399), .S(n4124), .Z(n403) );
  MUX2_X1 U9538 ( .A(ram[1633]), .B(ram[1649]), .S(n4296), .Z(n404) );
  MUX2_X1 U9539 ( .A(ram[1601]), .B(ram[1617]), .S(n4296), .Z(n405) );
  MUX2_X1 U9540 ( .A(n405), .B(n404), .S(n4183), .Z(n406) );
  MUX2_X1 U9541 ( .A(ram[1569]), .B(ram[1585]), .S(n4296), .Z(n407) );
  MUX2_X1 U9542 ( .A(ram[1537]), .B(ram[1553]), .S(n4296), .Z(n408) );
  MUX2_X1 U9543 ( .A(n408), .B(n407), .S(n4183), .Z(n409) );
  MUX2_X1 U9544 ( .A(n409), .B(n406), .S(n4124), .Z(n410) );
  MUX2_X1 U9545 ( .A(n410), .B(n403), .S(n4089), .Z(n411) );
  MUX2_X1 U9546 ( .A(n411), .B(n396), .S(n4077), .Z(n412) );
  MUX2_X1 U9547 ( .A(ram[1505]), .B(ram[1521]), .S(n4296), .Z(n413) );
  MUX2_X1 U9548 ( .A(ram[1473]), .B(ram[1489]), .S(n4296), .Z(n414) );
  MUX2_X1 U9549 ( .A(n414), .B(n413), .S(n4183), .Z(n415) );
  MUX2_X1 U9550 ( .A(ram[1441]), .B(ram[1457]), .S(n4296), .Z(n416) );
  MUX2_X1 U9551 ( .A(ram[1409]), .B(ram[1425]), .S(n4296), .Z(n417) );
  MUX2_X1 U9552 ( .A(n417), .B(n416), .S(n4183), .Z(n418) );
  MUX2_X1 U9553 ( .A(n418), .B(n415), .S(n4124), .Z(n419) );
  MUX2_X1 U9554 ( .A(ram[1377]), .B(ram[1393]), .S(n4297), .Z(n420) );
  MUX2_X1 U9555 ( .A(ram[1345]), .B(ram[1361]), .S(n4297), .Z(n421) );
  MUX2_X1 U9556 ( .A(n421), .B(n420), .S(n4183), .Z(n422) );
  MUX2_X1 U9557 ( .A(ram[1313]), .B(ram[1329]), .S(n4297), .Z(n423) );
  MUX2_X1 U9558 ( .A(ram[1281]), .B(ram[1297]), .S(n4297), .Z(n424) );
  MUX2_X1 U9559 ( .A(n424), .B(n423), .S(n4183), .Z(n425) );
  MUX2_X1 U9560 ( .A(n425), .B(n422), .S(n4124), .Z(n426) );
  MUX2_X1 U9561 ( .A(n426), .B(n419), .S(n4089), .Z(n427) );
  MUX2_X1 U9562 ( .A(ram[1249]), .B(ram[1265]), .S(n4297), .Z(n428) );
  MUX2_X1 U9563 ( .A(ram[1217]), .B(ram[1233]), .S(n4297), .Z(n429) );
  MUX2_X1 U9564 ( .A(n429), .B(n428), .S(n4183), .Z(n430) );
  MUX2_X1 U9565 ( .A(ram[1185]), .B(ram[1201]), .S(n4297), .Z(n431) );
  MUX2_X1 U9566 ( .A(ram[1153]), .B(ram[1169]), .S(n4297), .Z(n432) );
  MUX2_X1 U9567 ( .A(n432), .B(n431), .S(n4183), .Z(n433) );
  MUX2_X1 U9568 ( .A(n433), .B(n430), .S(n4124), .Z(n434) );
  MUX2_X1 U9569 ( .A(ram[1121]), .B(ram[1137]), .S(n4297), .Z(n435) );
  MUX2_X1 U9570 ( .A(ram[1089]), .B(ram[1105]), .S(n4297), .Z(n436) );
  MUX2_X1 U9571 ( .A(n436), .B(n435), .S(n4183), .Z(n437) );
  MUX2_X1 U9572 ( .A(ram[1057]), .B(ram[1073]), .S(n4297), .Z(n438) );
  MUX2_X1 U9573 ( .A(ram[1025]), .B(ram[1041]), .S(n4297), .Z(n439) );
  MUX2_X1 U9574 ( .A(n439), .B(n438), .S(n4183), .Z(n440) );
  MUX2_X1 U9575 ( .A(n440), .B(n437), .S(n4124), .Z(n441) );
  MUX2_X1 U9576 ( .A(n441), .B(n434), .S(n4089), .Z(n442) );
  MUX2_X1 U9577 ( .A(n442), .B(n427), .S(n4077), .Z(n443) );
  MUX2_X1 U9578 ( .A(n443), .B(n412), .S(n4069), .Z(n444) );
  MUX2_X1 U9579 ( .A(ram[993]), .B(ram[1009]), .S(n4298), .Z(n445) );
  MUX2_X1 U9580 ( .A(ram[961]), .B(ram[977]), .S(n4298), .Z(n446) );
  MUX2_X1 U9581 ( .A(n446), .B(n445), .S(n4184), .Z(n447) );
  MUX2_X1 U9582 ( .A(ram[929]), .B(ram[945]), .S(n4298), .Z(n448) );
  MUX2_X1 U9583 ( .A(ram[897]), .B(ram[913]), .S(n4298), .Z(n449) );
  MUX2_X1 U9584 ( .A(n449), .B(n448), .S(n4184), .Z(n450) );
  MUX2_X1 U9585 ( .A(n450), .B(n447), .S(n4125), .Z(n451) );
  MUX2_X1 U9586 ( .A(ram[865]), .B(ram[881]), .S(n4298), .Z(n452) );
  MUX2_X1 U9587 ( .A(ram[833]), .B(ram[849]), .S(n4298), .Z(n453) );
  MUX2_X1 U9588 ( .A(n453), .B(n452), .S(n4184), .Z(n454) );
  MUX2_X1 U9589 ( .A(ram[801]), .B(ram[817]), .S(n4298), .Z(n455) );
  MUX2_X1 U9590 ( .A(ram[769]), .B(ram[785]), .S(n4298), .Z(n456) );
  MUX2_X1 U9591 ( .A(n456), .B(n455), .S(n4184), .Z(n457) );
  MUX2_X1 U9592 ( .A(n457), .B(n454), .S(n4125), .Z(n458) );
  MUX2_X1 U9593 ( .A(n458), .B(n451), .S(n4090), .Z(n459) );
  MUX2_X1 U9594 ( .A(ram[737]), .B(ram[753]), .S(n4298), .Z(n460) );
  MUX2_X1 U9595 ( .A(ram[705]), .B(ram[721]), .S(n4298), .Z(n461) );
  MUX2_X1 U9596 ( .A(n461), .B(n460), .S(n4184), .Z(n462) );
  MUX2_X1 U9597 ( .A(ram[673]), .B(ram[689]), .S(n4298), .Z(n463) );
  MUX2_X1 U9598 ( .A(ram[641]), .B(ram[657]), .S(n4298), .Z(n464) );
  MUX2_X1 U9599 ( .A(n464), .B(n463), .S(n4184), .Z(n465) );
  MUX2_X1 U9600 ( .A(n465), .B(n462), .S(n4125), .Z(n466) );
  MUX2_X1 U9601 ( .A(ram[609]), .B(ram[625]), .S(n4299), .Z(n467) );
  MUX2_X1 U9602 ( .A(ram[577]), .B(ram[593]), .S(n4299), .Z(n468) );
  MUX2_X1 U9603 ( .A(n468), .B(n467), .S(n4184), .Z(n469) );
  MUX2_X1 U9604 ( .A(ram[545]), .B(ram[561]), .S(n4299), .Z(n470) );
  MUX2_X1 U9605 ( .A(ram[513]), .B(ram[529]), .S(n4299), .Z(n471) );
  MUX2_X1 U9606 ( .A(n471), .B(n470), .S(n4184), .Z(n472) );
  MUX2_X1 U9607 ( .A(n472), .B(n469), .S(n4125), .Z(n473) );
  MUX2_X1 U9608 ( .A(n473), .B(n466), .S(n4090), .Z(n474) );
  MUX2_X1 U9609 ( .A(n474), .B(n459), .S(n4077), .Z(n475) );
  MUX2_X1 U9610 ( .A(ram[481]), .B(ram[497]), .S(n4299), .Z(n476) );
  MUX2_X1 U9611 ( .A(ram[449]), .B(ram[465]), .S(n4299), .Z(n477) );
  MUX2_X1 U9612 ( .A(n477), .B(n476), .S(n4184), .Z(n478) );
  MUX2_X1 U9613 ( .A(ram[417]), .B(ram[433]), .S(n4299), .Z(n479) );
  MUX2_X1 U9614 ( .A(ram[385]), .B(ram[401]), .S(n4299), .Z(n480) );
  MUX2_X1 U9615 ( .A(n480), .B(n479), .S(n4184), .Z(n481) );
  MUX2_X1 U9616 ( .A(n481), .B(n478), .S(n4125), .Z(n482) );
  MUX2_X1 U9617 ( .A(ram[353]), .B(ram[369]), .S(n4299), .Z(n483) );
  MUX2_X1 U9618 ( .A(ram[321]), .B(ram[337]), .S(n4299), .Z(n484) );
  MUX2_X1 U9619 ( .A(n484), .B(n483), .S(n4184), .Z(n485) );
  MUX2_X1 U9620 ( .A(ram[289]), .B(ram[305]), .S(n4299), .Z(n486) );
  MUX2_X1 U9621 ( .A(ram[257]), .B(ram[273]), .S(n4299), .Z(n487) );
  MUX2_X1 U9622 ( .A(n487), .B(n486), .S(n4184), .Z(n488) );
  MUX2_X1 U9623 ( .A(n488), .B(n485), .S(n4125), .Z(n489) );
  MUX2_X1 U9624 ( .A(n489), .B(n482), .S(n4090), .Z(n490) );
  MUX2_X1 U9625 ( .A(ram[225]), .B(ram[241]), .S(n4300), .Z(n491) );
  MUX2_X1 U9626 ( .A(ram[193]), .B(ram[209]), .S(n4300), .Z(n492) );
  MUX2_X1 U9627 ( .A(n492), .B(n491), .S(n4185), .Z(n493) );
  MUX2_X1 U9628 ( .A(ram[161]), .B(ram[177]), .S(n4300), .Z(n494) );
  MUX2_X1 U9629 ( .A(ram[129]), .B(ram[145]), .S(n4300), .Z(n495) );
  MUX2_X1 U9630 ( .A(n495), .B(n494), .S(n4185), .Z(n496) );
  MUX2_X1 U9631 ( .A(n496), .B(n493), .S(n4125), .Z(n497) );
  MUX2_X1 U9632 ( .A(ram[97]), .B(ram[113]), .S(n4300), .Z(n498) );
  MUX2_X1 U9633 ( .A(ram[65]), .B(ram[81]), .S(n4300), .Z(n499) );
  MUX2_X1 U9634 ( .A(n499), .B(n498), .S(n4185), .Z(n500) );
  MUX2_X1 U9635 ( .A(ram[33]), .B(ram[49]), .S(n4300), .Z(n501) );
  MUX2_X1 U9636 ( .A(ram[1]), .B(ram[17]), .S(n4300), .Z(n502) );
  MUX2_X1 U9637 ( .A(n502), .B(n501), .S(n4185), .Z(n503) );
  MUX2_X1 U9638 ( .A(n503), .B(n500), .S(n4125), .Z(n504) );
  MUX2_X1 U9639 ( .A(n504), .B(n497), .S(n4090), .Z(n505) );
  MUX2_X1 U9640 ( .A(n505), .B(n490), .S(n4077), .Z(n506) );
  MUX2_X1 U9641 ( .A(n506), .B(n475), .S(n4069), .Z(n507) );
  MUX2_X1 U9642 ( .A(n507), .B(n444), .S(n4065), .Z(n508) );
  MUX2_X1 U9643 ( .A(n508), .B(n381), .S(mem_access_addr[9]), .Z(N300) );
  MUX2_X1 U9644 ( .A(ram[4066]), .B(ram[4082]), .S(n4300), .Z(n509) );
  MUX2_X1 U9645 ( .A(ram[4034]), .B(ram[4050]), .S(n4300), .Z(n510) );
  MUX2_X1 U9646 ( .A(n510), .B(n509), .S(n4185), .Z(n511) );
  MUX2_X1 U9647 ( .A(ram[4002]), .B(ram[4018]), .S(n4300), .Z(n512) );
  MUX2_X1 U9648 ( .A(ram[3970]), .B(ram[3986]), .S(n4300), .Z(n513) );
  MUX2_X1 U9649 ( .A(n513), .B(n512), .S(n4185), .Z(n514) );
  MUX2_X1 U9650 ( .A(n514), .B(n511), .S(n4125), .Z(n515) );
  MUX2_X1 U9651 ( .A(ram[3938]), .B(ram[3954]), .S(n4301), .Z(n516) );
  MUX2_X1 U9652 ( .A(ram[3906]), .B(ram[3922]), .S(n4301), .Z(n517) );
  MUX2_X1 U9653 ( .A(n517), .B(n516), .S(n4185), .Z(n518) );
  MUX2_X1 U9654 ( .A(ram[3874]), .B(ram[3890]), .S(n4301), .Z(n519) );
  MUX2_X1 U9655 ( .A(ram[3842]), .B(ram[3858]), .S(n4301), .Z(n520) );
  MUX2_X1 U9656 ( .A(n520), .B(n519), .S(n4185), .Z(n521) );
  MUX2_X1 U9657 ( .A(n521), .B(n518), .S(n4125), .Z(n522) );
  MUX2_X1 U9658 ( .A(n522), .B(n515), .S(n4090), .Z(n523) );
  MUX2_X1 U9659 ( .A(ram[3810]), .B(ram[3826]), .S(n4301), .Z(n524) );
  MUX2_X1 U9660 ( .A(ram[3778]), .B(ram[3794]), .S(n4301), .Z(n525) );
  MUX2_X1 U9661 ( .A(n525), .B(n524), .S(n4185), .Z(n526) );
  MUX2_X1 U9662 ( .A(ram[3746]), .B(ram[3762]), .S(n4301), .Z(n527) );
  MUX2_X1 U9663 ( .A(ram[3714]), .B(ram[3730]), .S(n4301), .Z(n528) );
  MUX2_X1 U9664 ( .A(n528), .B(n527), .S(n4185), .Z(n529) );
  MUX2_X1 U9665 ( .A(n529), .B(n526), .S(n4125), .Z(n530) );
  MUX2_X1 U9666 ( .A(ram[3682]), .B(ram[3698]), .S(n4301), .Z(n531) );
  MUX2_X1 U9667 ( .A(ram[3650]), .B(ram[3666]), .S(n4301), .Z(n532) );
  MUX2_X1 U9668 ( .A(n532), .B(n531), .S(n4185), .Z(n533) );
  MUX2_X1 U9669 ( .A(ram[3618]), .B(ram[3634]), .S(n4301), .Z(n534) );
  MUX2_X1 U9670 ( .A(ram[3586]), .B(ram[3602]), .S(n4301), .Z(n535) );
  MUX2_X1 U9671 ( .A(n535), .B(n534), .S(n4185), .Z(n536) );
  MUX2_X1 U9672 ( .A(n536), .B(n533), .S(n4125), .Z(n537) );
  MUX2_X1 U9673 ( .A(n537), .B(n530), .S(n4090), .Z(n538) );
  MUX2_X1 U9674 ( .A(n538), .B(n523), .S(n4077), .Z(n539) );
  MUX2_X1 U9675 ( .A(ram[3554]), .B(ram[3570]), .S(n4302), .Z(n540) );
  MUX2_X1 U9676 ( .A(ram[3522]), .B(ram[3538]), .S(n4302), .Z(n541) );
  MUX2_X1 U9677 ( .A(n541), .B(n540), .S(n4186), .Z(n542) );
  MUX2_X1 U9678 ( .A(ram[3490]), .B(ram[3506]), .S(n4302), .Z(n543) );
  MUX2_X1 U9679 ( .A(ram[3458]), .B(ram[3474]), .S(n4302), .Z(n544) );
  MUX2_X1 U9680 ( .A(n544), .B(n543), .S(n4186), .Z(n545) );
  MUX2_X1 U9681 ( .A(n545), .B(n542), .S(n4126), .Z(n546) );
  MUX2_X1 U9682 ( .A(ram[3426]), .B(ram[3442]), .S(n4302), .Z(n547) );
  MUX2_X1 U9683 ( .A(ram[3394]), .B(ram[3410]), .S(n4302), .Z(n548) );
  MUX2_X1 U9684 ( .A(n548), .B(n547), .S(n4186), .Z(n549) );
  MUX2_X1 U9685 ( .A(ram[3362]), .B(ram[3378]), .S(n4302), .Z(n550) );
  MUX2_X1 U9686 ( .A(ram[3330]), .B(ram[3346]), .S(n4302), .Z(n551) );
  MUX2_X1 U9687 ( .A(n551), .B(n550), .S(n4186), .Z(n552) );
  MUX2_X1 U9688 ( .A(n552), .B(n549), .S(n4126), .Z(n553) );
  MUX2_X1 U9689 ( .A(n553), .B(n546), .S(n4090), .Z(n554) );
  MUX2_X1 U9690 ( .A(ram[3298]), .B(ram[3314]), .S(n4302), .Z(n555) );
  MUX2_X1 U9691 ( .A(ram[3266]), .B(ram[3282]), .S(n4302), .Z(n556) );
  MUX2_X1 U9692 ( .A(n556), .B(n555), .S(n4186), .Z(n557) );
  MUX2_X1 U9693 ( .A(ram[3234]), .B(ram[3250]), .S(n4302), .Z(n558) );
  MUX2_X1 U9694 ( .A(ram[3202]), .B(ram[3218]), .S(n4302), .Z(n559) );
  MUX2_X1 U9695 ( .A(n559), .B(n558), .S(n4186), .Z(n560) );
  MUX2_X1 U9696 ( .A(n560), .B(n557), .S(n4126), .Z(n561) );
  MUX2_X1 U9697 ( .A(ram[3170]), .B(ram[3186]), .S(n4303), .Z(n562) );
  MUX2_X1 U9698 ( .A(ram[3138]), .B(ram[3154]), .S(n4303), .Z(n563) );
  MUX2_X1 U9699 ( .A(n563), .B(n562), .S(n4186), .Z(n564) );
  MUX2_X1 U9700 ( .A(ram[3106]), .B(ram[3122]), .S(n4303), .Z(n565) );
  MUX2_X1 U9701 ( .A(ram[3074]), .B(ram[3090]), .S(n4303), .Z(n566) );
  MUX2_X1 U9702 ( .A(n566), .B(n565), .S(n4186), .Z(n567) );
  MUX2_X1 U9703 ( .A(n567), .B(n564), .S(n4126), .Z(n568) );
  MUX2_X1 U9704 ( .A(n568), .B(n561), .S(n4090), .Z(n569) );
  MUX2_X1 U9705 ( .A(n569), .B(n554), .S(n4077), .Z(n570) );
  MUX2_X1 U9706 ( .A(n570), .B(n539), .S(n4069), .Z(n571) );
  MUX2_X1 U9707 ( .A(ram[3042]), .B(ram[3058]), .S(n4303), .Z(n572) );
  MUX2_X1 U9708 ( .A(ram[3010]), .B(ram[3026]), .S(n4303), .Z(n573) );
  MUX2_X1 U9709 ( .A(n573), .B(n572), .S(n4186), .Z(n574) );
  MUX2_X1 U9710 ( .A(ram[2978]), .B(ram[2994]), .S(n4303), .Z(n575) );
  MUX2_X1 U9711 ( .A(ram[2946]), .B(ram[2962]), .S(n4303), .Z(n576) );
  MUX2_X1 U9712 ( .A(n576), .B(n575), .S(n4186), .Z(n577) );
  MUX2_X1 U9713 ( .A(n577), .B(n574), .S(n4126), .Z(n578) );
  MUX2_X1 U9714 ( .A(ram[2914]), .B(ram[2930]), .S(n4303), .Z(n579) );
  MUX2_X1 U9715 ( .A(ram[2882]), .B(ram[2898]), .S(n4303), .Z(n580) );
  MUX2_X1 U9716 ( .A(n580), .B(n579), .S(n4186), .Z(n581) );
  MUX2_X1 U9717 ( .A(ram[2850]), .B(ram[2866]), .S(n4303), .Z(n582) );
  MUX2_X1 U9718 ( .A(ram[2818]), .B(ram[2834]), .S(n4303), .Z(n583) );
  MUX2_X1 U9719 ( .A(n583), .B(n582), .S(n4186), .Z(n584) );
  MUX2_X1 U9720 ( .A(n584), .B(n581), .S(n4126), .Z(n585) );
  MUX2_X1 U9721 ( .A(n585), .B(n578), .S(n4090), .Z(n586) );
  MUX2_X1 U9722 ( .A(ram[2786]), .B(ram[2802]), .S(n4304), .Z(n587) );
  MUX2_X1 U9723 ( .A(ram[2754]), .B(ram[2770]), .S(n4304), .Z(n588) );
  MUX2_X1 U9724 ( .A(n588), .B(n587), .S(n4187), .Z(n589) );
  MUX2_X1 U9725 ( .A(ram[2722]), .B(ram[2738]), .S(n4304), .Z(n590) );
  MUX2_X1 U9726 ( .A(ram[2690]), .B(ram[2706]), .S(n4304), .Z(n591) );
  MUX2_X1 U9727 ( .A(n591), .B(n590), .S(n4187), .Z(n592) );
  MUX2_X1 U9728 ( .A(n592), .B(n589), .S(n4126), .Z(n593) );
  MUX2_X1 U9729 ( .A(ram[2658]), .B(ram[2674]), .S(n4304), .Z(n594) );
  MUX2_X1 U9730 ( .A(ram[2626]), .B(ram[2642]), .S(n4304), .Z(n595) );
  MUX2_X1 U9731 ( .A(n595), .B(n594), .S(n4187), .Z(n596) );
  MUX2_X1 U9732 ( .A(ram[2594]), .B(ram[2610]), .S(n4304), .Z(n597) );
  MUX2_X1 U9733 ( .A(ram[2562]), .B(ram[2578]), .S(n4304), .Z(n598) );
  MUX2_X1 U9734 ( .A(n598), .B(n597), .S(n4187), .Z(n599) );
  MUX2_X1 U9735 ( .A(n599), .B(n596), .S(n4126), .Z(n600) );
  MUX2_X1 U9736 ( .A(n600), .B(n593), .S(n4090), .Z(n601) );
  MUX2_X1 U9737 ( .A(n601), .B(n586), .S(n4077), .Z(n602) );
  MUX2_X1 U9738 ( .A(ram[2530]), .B(ram[2546]), .S(n4304), .Z(n603) );
  MUX2_X1 U9739 ( .A(ram[2498]), .B(ram[2514]), .S(n4304), .Z(n604) );
  MUX2_X1 U9740 ( .A(n604), .B(n603), .S(n4187), .Z(n605) );
  MUX2_X1 U9741 ( .A(ram[2466]), .B(ram[2482]), .S(n4304), .Z(n606) );
  MUX2_X1 U9742 ( .A(ram[2434]), .B(ram[2450]), .S(n4304), .Z(n607) );
  MUX2_X1 U9743 ( .A(n607), .B(n606), .S(n4187), .Z(n608) );
  MUX2_X1 U9744 ( .A(n608), .B(n605), .S(n4126), .Z(n609) );
  MUX2_X1 U9745 ( .A(ram[2402]), .B(ram[2418]), .S(n4305), .Z(n610) );
  MUX2_X1 U9746 ( .A(ram[2370]), .B(ram[2386]), .S(n4305), .Z(n611) );
  MUX2_X1 U9747 ( .A(n611), .B(n610), .S(n4187), .Z(n612) );
  MUX2_X1 U9748 ( .A(ram[2338]), .B(ram[2354]), .S(n4305), .Z(n613) );
  MUX2_X1 U9749 ( .A(ram[2306]), .B(ram[2322]), .S(n4305), .Z(n614) );
  MUX2_X1 U9750 ( .A(n614), .B(n613), .S(n4187), .Z(n615) );
  MUX2_X1 U9751 ( .A(n615), .B(n612), .S(n4126), .Z(n616) );
  MUX2_X1 U9752 ( .A(n616), .B(n609), .S(n4090), .Z(n617) );
  MUX2_X1 U9753 ( .A(ram[2274]), .B(ram[2290]), .S(n4305), .Z(n618) );
  MUX2_X1 U9754 ( .A(ram[2242]), .B(ram[2258]), .S(n4305), .Z(n619) );
  MUX2_X1 U9755 ( .A(n619), .B(n618), .S(n4187), .Z(n620) );
  MUX2_X1 U9756 ( .A(ram[2210]), .B(ram[2226]), .S(n4305), .Z(n621) );
  MUX2_X1 U9757 ( .A(ram[2178]), .B(ram[2194]), .S(n4305), .Z(n622) );
  MUX2_X1 U9758 ( .A(n622), .B(n621), .S(n4187), .Z(n623) );
  MUX2_X1 U9759 ( .A(n623), .B(n620), .S(n4126), .Z(n624) );
  MUX2_X1 U9760 ( .A(ram[2146]), .B(ram[2162]), .S(n4305), .Z(n625) );
  MUX2_X1 U9761 ( .A(ram[2114]), .B(ram[2130]), .S(n4305), .Z(n626) );
  MUX2_X1 U9762 ( .A(n626), .B(n625), .S(n4187), .Z(n627) );
  MUX2_X1 U9763 ( .A(ram[2082]), .B(ram[2098]), .S(n4305), .Z(n628) );
  MUX2_X1 U9764 ( .A(ram[2050]), .B(ram[2066]), .S(n4305), .Z(n629) );
  MUX2_X1 U9765 ( .A(n629), .B(n628), .S(n4187), .Z(n630) );
  MUX2_X1 U9766 ( .A(n630), .B(n627), .S(n4126), .Z(n631) );
  MUX2_X1 U9767 ( .A(n631), .B(n624), .S(n4090), .Z(n632) );
  MUX2_X1 U9768 ( .A(n632), .B(n617), .S(n4077), .Z(n633) );
  MUX2_X1 U9769 ( .A(n633), .B(n602), .S(n4069), .Z(n634) );
  MUX2_X1 U9770 ( .A(n634), .B(n571), .S(n4065), .Z(n635) );
  MUX2_X1 U9771 ( .A(ram[2018]), .B(ram[2034]), .S(n4306), .Z(n636) );
  MUX2_X1 U9772 ( .A(ram[1986]), .B(ram[2002]), .S(n4306), .Z(n637) );
  MUX2_X1 U9773 ( .A(n637), .B(n636), .S(n4188), .Z(n638) );
  MUX2_X1 U9774 ( .A(ram[1954]), .B(ram[1970]), .S(n4306), .Z(n639) );
  MUX2_X1 U9775 ( .A(ram[1922]), .B(ram[1938]), .S(n4306), .Z(n640) );
  MUX2_X1 U9776 ( .A(n640), .B(n639), .S(n4188), .Z(n641) );
  MUX2_X1 U9777 ( .A(n641), .B(n638), .S(n4127), .Z(n642) );
  MUX2_X1 U9778 ( .A(ram[1890]), .B(ram[1906]), .S(n4306), .Z(n643) );
  MUX2_X1 U9779 ( .A(ram[1858]), .B(ram[1874]), .S(n4306), .Z(n644) );
  MUX2_X1 U9780 ( .A(n644), .B(n643), .S(n4188), .Z(n645) );
  MUX2_X1 U9781 ( .A(ram[1826]), .B(ram[1842]), .S(n4306), .Z(n646) );
  MUX2_X1 U9782 ( .A(ram[1794]), .B(ram[1810]), .S(n4306), .Z(n647) );
  MUX2_X1 U9783 ( .A(n647), .B(n646), .S(n4188), .Z(n648) );
  MUX2_X1 U9784 ( .A(n648), .B(n645), .S(n4127), .Z(n649) );
  MUX2_X1 U9785 ( .A(n649), .B(n642), .S(n4091), .Z(n650) );
  MUX2_X1 U9786 ( .A(ram[1762]), .B(ram[1778]), .S(n4306), .Z(n651) );
  MUX2_X1 U9787 ( .A(ram[1730]), .B(ram[1746]), .S(n4306), .Z(n652) );
  MUX2_X1 U9788 ( .A(n652), .B(n651), .S(n4188), .Z(n653) );
  MUX2_X1 U9789 ( .A(ram[1698]), .B(ram[1714]), .S(n4306), .Z(n654) );
  MUX2_X1 U9790 ( .A(ram[1666]), .B(ram[1682]), .S(n4306), .Z(n655) );
  MUX2_X1 U9791 ( .A(n655), .B(n654), .S(n4188), .Z(n656) );
  MUX2_X1 U9792 ( .A(n656), .B(n653), .S(n4127), .Z(n657) );
  MUX2_X1 U9793 ( .A(ram[1634]), .B(ram[1650]), .S(n4307), .Z(n658) );
  MUX2_X1 U9794 ( .A(ram[1602]), .B(ram[1618]), .S(n4307), .Z(n659) );
  MUX2_X1 U9795 ( .A(n659), .B(n658), .S(n4188), .Z(n660) );
  MUX2_X1 U9796 ( .A(ram[1570]), .B(ram[1586]), .S(n4307), .Z(n661) );
  MUX2_X1 U9797 ( .A(ram[1538]), .B(ram[1554]), .S(n4307), .Z(n662) );
  MUX2_X1 U9798 ( .A(n662), .B(n661), .S(n4188), .Z(n663) );
  MUX2_X1 U9799 ( .A(n663), .B(n660), .S(n4127), .Z(n664) );
  MUX2_X1 U9800 ( .A(n664), .B(n657), .S(n4091), .Z(n665) );
  MUX2_X1 U9801 ( .A(n665), .B(n650), .S(n4078), .Z(n666) );
  MUX2_X1 U9802 ( .A(ram[1506]), .B(ram[1522]), .S(n4307), .Z(n667) );
  MUX2_X1 U9803 ( .A(ram[1474]), .B(ram[1490]), .S(n4307), .Z(n668) );
  MUX2_X1 U9804 ( .A(n668), .B(n667), .S(n4188), .Z(n669) );
  MUX2_X1 U9805 ( .A(ram[1442]), .B(ram[1458]), .S(n4307), .Z(n670) );
  MUX2_X1 U9806 ( .A(ram[1410]), .B(ram[1426]), .S(n4307), .Z(n671) );
  MUX2_X1 U9807 ( .A(n671), .B(n670), .S(n4188), .Z(n672) );
  MUX2_X1 U9808 ( .A(n672), .B(n669), .S(n4127), .Z(n673) );
  MUX2_X1 U9809 ( .A(ram[1378]), .B(ram[1394]), .S(n4307), .Z(n674) );
  MUX2_X1 U9810 ( .A(ram[1346]), .B(ram[1362]), .S(n4307), .Z(n675) );
  MUX2_X1 U9811 ( .A(n675), .B(n674), .S(n4188), .Z(n676) );
  MUX2_X1 U9812 ( .A(ram[1314]), .B(ram[1330]), .S(n4307), .Z(n677) );
  MUX2_X1 U9813 ( .A(ram[1282]), .B(ram[1298]), .S(n4307), .Z(n678) );
  MUX2_X1 U9814 ( .A(n678), .B(n677), .S(n4188), .Z(n679) );
  MUX2_X1 U9815 ( .A(n679), .B(n676), .S(n4127), .Z(n680) );
  MUX2_X1 U9816 ( .A(n680), .B(n673), .S(n4091), .Z(n681) );
  MUX2_X1 U9817 ( .A(ram[1250]), .B(ram[1266]), .S(n4308), .Z(n682) );
  MUX2_X1 U9818 ( .A(ram[1218]), .B(ram[1234]), .S(n4308), .Z(n683) );
  MUX2_X1 U9819 ( .A(n683), .B(n682), .S(n4189), .Z(n684) );
  MUX2_X1 U9820 ( .A(ram[1186]), .B(ram[1202]), .S(n4308), .Z(n685) );
  MUX2_X1 U9821 ( .A(ram[1154]), .B(ram[1170]), .S(n4308), .Z(n686) );
  MUX2_X1 U9822 ( .A(n686), .B(n685), .S(n4189), .Z(n687) );
  MUX2_X1 U9823 ( .A(n687), .B(n684), .S(n4127), .Z(n688) );
  MUX2_X1 U9824 ( .A(ram[1122]), .B(ram[1138]), .S(n4308), .Z(n689) );
  MUX2_X1 U9825 ( .A(ram[1090]), .B(ram[1106]), .S(n4308), .Z(n690) );
  MUX2_X1 U9826 ( .A(n690), .B(n689), .S(n4189), .Z(n691) );
  MUX2_X1 U9827 ( .A(ram[1058]), .B(ram[1074]), .S(n4308), .Z(n692) );
  MUX2_X1 U9828 ( .A(ram[1026]), .B(ram[1042]), .S(n4308), .Z(n693) );
  MUX2_X1 U9829 ( .A(n693), .B(n692), .S(n4189), .Z(n694) );
  MUX2_X1 U9830 ( .A(n694), .B(n691), .S(n4127), .Z(n695) );
  MUX2_X1 U9831 ( .A(n695), .B(n688), .S(n4091), .Z(n696) );
  MUX2_X1 U9832 ( .A(n696), .B(n681), .S(n4078), .Z(n697) );
  MUX2_X1 U9833 ( .A(n697), .B(n666), .S(n4069), .Z(n698) );
  MUX2_X1 U9834 ( .A(ram[994]), .B(ram[1010]), .S(n4308), .Z(n699) );
  MUX2_X1 U9835 ( .A(ram[962]), .B(ram[978]), .S(n4308), .Z(n700) );
  MUX2_X1 U9836 ( .A(n700), .B(n699), .S(n4189), .Z(n701) );
  MUX2_X1 U9837 ( .A(ram[930]), .B(ram[946]), .S(n4308), .Z(n702) );
  MUX2_X1 U9838 ( .A(ram[898]), .B(ram[914]), .S(n4308), .Z(n703) );
  MUX2_X1 U9839 ( .A(n703), .B(n702), .S(n4189), .Z(n704) );
  MUX2_X1 U9840 ( .A(n704), .B(n701), .S(n4127), .Z(n705) );
  MUX2_X1 U9841 ( .A(ram[866]), .B(ram[882]), .S(n4309), .Z(n706) );
  MUX2_X1 U9842 ( .A(ram[834]), .B(ram[850]), .S(n4309), .Z(n707) );
  MUX2_X1 U9843 ( .A(n707), .B(n706), .S(n4189), .Z(n708) );
  MUX2_X1 U9844 ( .A(ram[802]), .B(ram[818]), .S(n4309), .Z(n709) );
  MUX2_X1 U9845 ( .A(ram[770]), .B(ram[786]), .S(n4309), .Z(n710) );
  MUX2_X1 U9846 ( .A(n710), .B(n709), .S(n4189), .Z(n711) );
  MUX2_X1 U9847 ( .A(n711), .B(n708), .S(n4127), .Z(n712) );
  MUX2_X1 U9848 ( .A(n712), .B(n705), .S(n4091), .Z(n713) );
  MUX2_X1 U9849 ( .A(ram[738]), .B(ram[754]), .S(n4309), .Z(n714) );
  MUX2_X1 U9850 ( .A(ram[706]), .B(ram[722]), .S(n4309), .Z(n715) );
  MUX2_X1 U9851 ( .A(n715), .B(n714), .S(n4189), .Z(n716) );
  MUX2_X1 U9852 ( .A(ram[674]), .B(ram[690]), .S(n4309), .Z(n717) );
  MUX2_X1 U9853 ( .A(ram[642]), .B(ram[658]), .S(n4309), .Z(n718) );
  MUX2_X1 U9854 ( .A(n718), .B(n717), .S(n4189), .Z(n719) );
  MUX2_X1 U9855 ( .A(n719), .B(n716), .S(n4127), .Z(n720) );
  MUX2_X1 U9856 ( .A(ram[610]), .B(ram[626]), .S(n4309), .Z(n721) );
  MUX2_X1 U9857 ( .A(ram[578]), .B(ram[594]), .S(n4309), .Z(n722) );
  MUX2_X1 U9858 ( .A(n722), .B(n721), .S(n4189), .Z(n723) );
  MUX2_X1 U9859 ( .A(ram[546]), .B(ram[562]), .S(n4309), .Z(n724) );
  MUX2_X1 U9860 ( .A(ram[514]), .B(ram[530]), .S(n4309), .Z(n725) );
  MUX2_X1 U9861 ( .A(n725), .B(n724), .S(n4189), .Z(n726) );
  MUX2_X1 U9862 ( .A(n726), .B(n723), .S(n4127), .Z(n727) );
  MUX2_X1 U9863 ( .A(n727), .B(n720), .S(n4091), .Z(n728) );
  MUX2_X1 U9864 ( .A(n728), .B(n713), .S(n4078), .Z(n729) );
  MUX2_X1 U9865 ( .A(ram[482]), .B(ram[498]), .S(n4310), .Z(n730) );
  MUX2_X1 U9866 ( .A(ram[450]), .B(ram[466]), .S(n4310), .Z(n731) );
  MUX2_X1 U9867 ( .A(n731), .B(n730), .S(n4190), .Z(n732) );
  MUX2_X1 U9868 ( .A(ram[418]), .B(ram[434]), .S(n4310), .Z(n733) );
  MUX2_X1 U9869 ( .A(ram[386]), .B(ram[402]), .S(n4310), .Z(n734) );
  MUX2_X1 U9870 ( .A(n734), .B(n733), .S(n4190), .Z(n735) );
  MUX2_X1 U9871 ( .A(n735), .B(n732), .S(n4128), .Z(n736) );
  MUX2_X1 U9872 ( .A(ram[354]), .B(ram[370]), .S(n4310), .Z(n737) );
  MUX2_X1 U9873 ( .A(ram[322]), .B(ram[338]), .S(n4310), .Z(n738) );
  MUX2_X1 U9874 ( .A(n738), .B(n737), .S(n4190), .Z(n739) );
  MUX2_X1 U9875 ( .A(ram[290]), .B(ram[306]), .S(n4310), .Z(n740) );
  MUX2_X1 U9876 ( .A(ram[258]), .B(ram[274]), .S(n4310), .Z(n741) );
  MUX2_X1 U9877 ( .A(n741), .B(n740), .S(n4190), .Z(n742) );
  MUX2_X1 U9878 ( .A(n742), .B(n739), .S(n4128), .Z(n743) );
  MUX2_X1 U9879 ( .A(n743), .B(n736), .S(n4091), .Z(n744) );
  MUX2_X1 U9880 ( .A(ram[226]), .B(ram[242]), .S(n4310), .Z(n745) );
  MUX2_X1 U9881 ( .A(ram[194]), .B(ram[210]), .S(n4310), .Z(n746) );
  MUX2_X1 U9882 ( .A(n746), .B(n745), .S(n4190), .Z(n747) );
  MUX2_X1 U9883 ( .A(ram[162]), .B(ram[178]), .S(n4310), .Z(n748) );
  MUX2_X1 U9884 ( .A(ram[130]), .B(ram[146]), .S(n4310), .Z(n749) );
  MUX2_X1 U9885 ( .A(n749), .B(n748), .S(n4190), .Z(n750) );
  MUX2_X1 U9886 ( .A(n750), .B(n747), .S(n4128), .Z(n751) );
  MUX2_X1 U9887 ( .A(ram[98]), .B(ram[114]), .S(n4311), .Z(n752) );
  MUX2_X1 U9888 ( .A(ram[66]), .B(ram[82]), .S(n4311), .Z(n753) );
  MUX2_X1 U9889 ( .A(n753), .B(n752), .S(n4190), .Z(n754) );
  MUX2_X1 U9890 ( .A(ram[34]), .B(ram[50]), .S(n4311), .Z(n755) );
  MUX2_X1 U9891 ( .A(ram[2]), .B(ram[18]), .S(n4311), .Z(n756) );
  MUX2_X1 U9892 ( .A(n756), .B(n755), .S(n4190), .Z(n757) );
  MUX2_X1 U9893 ( .A(n757), .B(n754), .S(n4128), .Z(n758) );
  MUX2_X1 U9894 ( .A(n758), .B(n751), .S(n4091), .Z(n759) );
  MUX2_X1 U9895 ( .A(n759), .B(n744), .S(n4078), .Z(n760) );
  MUX2_X1 U9896 ( .A(n760), .B(n729), .S(n4069), .Z(n761) );
  MUX2_X1 U9897 ( .A(n761), .B(n698), .S(n4065), .Z(n762) );
  MUX2_X1 U9898 ( .A(n762), .B(n635), .S(mem_access_addr[9]), .Z(N299) );
  MUX2_X1 U9899 ( .A(ram[4067]), .B(ram[4083]), .S(n4311), .Z(n763) );
  MUX2_X1 U9900 ( .A(ram[4035]), .B(ram[4051]), .S(n4311), .Z(n764) );
  MUX2_X1 U9901 ( .A(n764), .B(n763), .S(n4190), .Z(n765) );
  MUX2_X1 U9902 ( .A(ram[4003]), .B(ram[4019]), .S(n4311), .Z(n766) );
  MUX2_X1 U9903 ( .A(ram[3971]), .B(ram[3987]), .S(n4311), .Z(n767) );
  MUX2_X1 U9904 ( .A(n767), .B(n766), .S(n4190), .Z(n768) );
  MUX2_X1 U9905 ( .A(n768), .B(n765), .S(n4128), .Z(n769) );
  MUX2_X1 U9906 ( .A(ram[3939]), .B(ram[3955]), .S(n4311), .Z(n770) );
  MUX2_X1 U9907 ( .A(ram[3907]), .B(ram[3923]), .S(n4311), .Z(n771) );
  MUX2_X1 U9908 ( .A(n771), .B(n770), .S(n4190), .Z(n772) );
  MUX2_X1 U9909 ( .A(ram[3875]), .B(ram[3891]), .S(n4311), .Z(n773) );
  MUX2_X1 U9910 ( .A(ram[3843]), .B(ram[3859]), .S(n4311), .Z(n774) );
  MUX2_X1 U9911 ( .A(n774), .B(n773), .S(n4190), .Z(n775) );
  MUX2_X1 U9912 ( .A(n775), .B(n772), .S(n4128), .Z(n776) );
  MUX2_X1 U9913 ( .A(n776), .B(n769), .S(n4091), .Z(n777) );
  MUX2_X1 U9914 ( .A(ram[3811]), .B(ram[3827]), .S(n4312), .Z(n778) );
  MUX2_X1 U9915 ( .A(ram[3779]), .B(ram[3795]), .S(n4312), .Z(n779) );
  MUX2_X1 U9916 ( .A(n779), .B(n778), .S(n4191), .Z(n780) );
  MUX2_X1 U9917 ( .A(ram[3747]), .B(ram[3763]), .S(n4312), .Z(n781) );
  MUX2_X1 U9918 ( .A(ram[3715]), .B(ram[3731]), .S(n4312), .Z(n782) );
  MUX2_X1 U9919 ( .A(n782), .B(n781), .S(n4191), .Z(n783) );
  MUX2_X1 U9920 ( .A(n783), .B(n780), .S(n4128), .Z(n784) );
  MUX2_X1 U9921 ( .A(ram[3683]), .B(ram[3699]), .S(n4312), .Z(n785) );
  MUX2_X1 U9922 ( .A(ram[3651]), .B(ram[3667]), .S(n4312), .Z(n786) );
  MUX2_X1 U9923 ( .A(n786), .B(n785), .S(n4191), .Z(n787) );
  MUX2_X1 U9924 ( .A(ram[3619]), .B(ram[3635]), .S(n4312), .Z(n788) );
  MUX2_X1 U9925 ( .A(ram[3587]), .B(ram[3603]), .S(n4312), .Z(n789) );
  MUX2_X1 U9926 ( .A(n789), .B(n788), .S(n4191), .Z(n790) );
  MUX2_X1 U9927 ( .A(n790), .B(n787), .S(n4128), .Z(n791) );
  MUX2_X1 U9928 ( .A(n791), .B(n784), .S(n4091), .Z(n792) );
  MUX2_X1 U9929 ( .A(n792), .B(n777), .S(n4078), .Z(n793) );
  MUX2_X1 U9930 ( .A(ram[3555]), .B(ram[3571]), .S(n4312), .Z(n794) );
  MUX2_X1 U9931 ( .A(ram[3523]), .B(ram[3539]), .S(n4312), .Z(n795) );
  MUX2_X1 U9932 ( .A(n795), .B(n794), .S(n4191), .Z(n796) );
  MUX2_X1 U9933 ( .A(ram[3491]), .B(ram[3507]), .S(n4312), .Z(n797) );
  MUX2_X1 U9934 ( .A(ram[3459]), .B(ram[3475]), .S(n4312), .Z(n798) );
  MUX2_X1 U9935 ( .A(n798), .B(n797), .S(n4191), .Z(n799) );
  MUX2_X1 U9936 ( .A(n799), .B(n796), .S(n4128), .Z(n800) );
  MUX2_X1 U9937 ( .A(ram[3427]), .B(ram[3443]), .S(n4313), .Z(n801) );
  MUX2_X1 U9938 ( .A(ram[3395]), .B(ram[3411]), .S(n4313), .Z(n802) );
  MUX2_X1 U9939 ( .A(n802), .B(n801), .S(n4191), .Z(n803) );
  MUX2_X1 U9940 ( .A(ram[3363]), .B(ram[3379]), .S(n4313), .Z(n804) );
  MUX2_X1 U9941 ( .A(ram[3331]), .B(ram[3347]), .S(n4313), .Z(n805) );
  MUX2_X1 U9942 ( .A(n805), .B(n804), .S(n4191), .Z(n806) );
  MUX2_X1 U9943 ( .A(n806), .B(n803), .S(n4128), .Z(n807) );
  MUX2_X1 U9944 ( .A(n807), .B(n800), .S(n4091), .Z(n808) );
  MUX2_X1 U9945 ( .A(ram[3299]), .B(ram[3315]), .S(n4313), .Z(n809) );
  MUX2_X1 U9946 ( .A(ram[3267]), .B(ram[3283]), .S(n4313), .Z(n810) );
  MUX2_X1 U9947 ( .A(n810), .B(n809), .S(n4191), .Z(n811) );
  MUX2_X1 U9948 ( .A(ram[3235]), .B(ram[3251]), .S(n4313), .Z(n812) );
  MUX2_X1 U9949 ( .A(ram[3203]), .B(ram[3219]), .S(n4313), .Z(n813) );
  MUX2_X1 U9950 ( .A(n813), .B(n812), .S(n4191), .Z(n814) );
  MUX2_X1 U9951 ( .A(n814), .B(n811), .S(n4128), .Z(n815) );
  MUX2_X1 U9952 ( .A(ram[3171]), .B(ram[3187]), .S(n4313), .Z(n816) );
  MUX2_X1 U9953 ( .A(ram[3139]), .B(ram[3155]), .S(n4313), .Z(n817) );
  MUX2_X1 U9954 ( .A(n817), .B(n816), .S(n4191), .Z(n818) );
  MUX2_X1 U9955 ( .A(ram[3107]), .B(ram[3123]), .S(n4313), .Z(n819) );
  MUX2_X1 U9956 ( .A(ram[3075]), .B(ram[3091]), .S(n4313), .Z(n820) );
  MUX2_X1 U9957 ( .A(n820), .B(n819), .S(n4191), .Z(n821) );
  MUX2_X1 U9958 ( .A(n821), .B(n818), .S(n4128), .Z(n822) );
  MUX2_X1 U9959 ( .A(n822), .B(n815), .S(n4091), .Z(n823) );
  MUX2_X1 U9960 ( .A(n823), .B(n808), .S(n4078), .Z(n824) );
  MUX2_X1 U9961 ( .A(n824), .B(n793), .S(n4069), .Z(n825) );
  MUX2_X1 U9962 ( .A(ram[3043]), .B(ram[3059]), .S(n4314), .Z(n826) );
  MUX2_X1 U9963 ( .A(ram[3011]), .B(ram[3027]), .S(n4314), .Z(n827) );
  MUX2_X1 U9964 ( .A(n827), .B(n826), .S(n4192), .Z(n828) );
  MUX2_X1 U9965 ( .A(ram[2979]), .B(ram[2995]), .S(n4314), .Z(n829) );
  MUX2_X1 U9966 ( .A(ram[2947]), .B(ram[2963]), .S(n4314), .Z(n830) );
  MUX2_X1 U9967 ( .A(n830), .B(n829), .S(n4192), .Z(n831) );
  MUX2_X1 U9968 ( .A(n831), .B(n828), .S(n4129), .Z(n832) );
  MUX2_X1 U9969 ( .A(ram[2915]), .B(ram[2931]), .S(n4314), .Z(n833) );
  MUX2_X1 U9970 ( .A(ram[2883]), .B(ram[2899]), .S(n4314), .Z(n834) );
  MUX2_X1 U9971 ( .A(n834), .B(n833), .S(n4192), .Z(n835) );
  MUX2_X1 U9972 ( .A(ram[2851]), .B(ram[2867]), .S(n4314), .Z(n836) );
  MUX2_X1 U9973 ( .A(ram[2819]), .B(ram[2835]), .S(n4314), .Z(n837) );
  MUX2_X1 U9974 ( .A(n837), .B(n836), .S(n4192), .Z(n838) );
  MUX2_X1 U9975 ( .A(n838), .B(n835), .S(n4129), .Z(n839) );
  MUX2_X1 U9976 ( .A(n839), .B(n832), .S(n4092), .Z(n840) );
  MUX2_X1 U9977 ( .A(ram[2787]), .B(ram[2803]), .S(n4314), .Z(n841) );
  MUX2_X1 U9978 ( .A(ram[2755]), .B(ram[2771]), .S(n4314), .Z(n842) );
  MUX2_X1 U9979 ( .A(n842), .B(n841), .S(n4192), .Z(n843) );
  MUX2_X1 U9980 ( .A(ram[2723]), .B(ram[2739]), .S(n4314), .Z(n844) );
  MUX2_X1 U9981 ( .A(ram[2691]), .B(ram[2707]), .S(n4314), .Z(n845) );
  MUX2_X1 U9982 ( .A(n845), .B(n844), .S(n4192), .Z(n846) );
  MUX2_X1 U9983 ( .A(n846), .B(n843), .S(n4129), .Z(n847) );
  MUX2_X1 U9984 ( .A(ram[2659]), .B(ram[2675]), .S(n4315), .Z(n848) );
  MUX2_X1 U9985 ( .A(ram[2627]), .B(ram[2643]), .S(n4315), .Z(n849) );
  MUX2_X1 U9986 ( .A(n849), .B(n848), .S(n4192), .Z(n850) );
  MUX2_X1 U9987 ( .A(ram[2595]), .B(ram[2611]), .S(n4315), .Z(n851) );
  MUX2_X1 U9988 ( .A(ram[2563]), .B(ram[2579]), .S(n4315), .Z(n852) );
  MUX2_X1 U9989 ( .A(n852), .B(n851), .S(n4192), .Z(n853) );
  MUX2_X1 U9990 ( .A(n853), .B(n850), .S(n4129), .Z(n854) );
  MUX2_X1 U9991 ( .A(n854), .B(n847), .S(n4092), .Z(n855) );
  MUX2_X1 U9992 ( .A(n855), .B(n840), .S(n4078), .Z(n856) );
  MUX2_X1 U9993 ( .A(ram[2531]), .B(ram[2547]), .S(n4315), .Z(n857) );
  MUX2_X1 U9994 ( .A(ram[2499]), .B(ram[2515]), .S(n4315), .Z(n858) );
  MUX2_X1 U9995 ( .A(n858), .B(n857), .S(n4192), .Z(n859) );
  MUX2_X1 U9996 ( .A(ram[2467]), .B(ram[2483]), .S(n4315), .Z(n860) );
  MUX2_X1 U9997 ( .A(ram[2435]), .B(ram[2451]), .S(n4315), .Z(n861) );
  MUX2_X1 U9998 ( .A(n861), .B(n860), .S(n4192), .Z(n862) );
  MUX2_X1 U9999 ( .A(n862), .B(n859), .S(n4129), .Z(n863) );
  MUX2_X1 U10000 ( .A(ram[2403]), .B(ram[2419]), .S(n4315), .Z(n864) );
  MUX2_X1 U10001 ( .A(ram[2371]), .B(ram[2387]), .S(n4315), .Z(n865) );
  MUX2_X1 U10002 ( .A(n865), .B(n864), .S(n4192), .Z(n866) );
  MUX2_X1 U10003 ( .A(ram[2339]), .B(ram[2355]), .S(n4315), .Z(n867) );
  MUX2_X1 U10004 ( .A(ram[2307]), .B(ram[2323]), .S(n4315), .Z(n868) );
  MUX2_X1 U10005 ( .A(n868), .B(n867), .S(n4192), .Z(n869) );
  MUX2_X1 U10006 ( .A(n869), .B(n866), .S(n4129), .Z(n870) );
  MUX2_X1 U10007 ( .A(n870), .B(n863), .S(n4092), .Z(n871) );
  MUX2_X1 U10008 ( .A(ram[2275]), .B(ram[2291]), .S(n4316), .Z(n872) );
  MUX2_X1 U10009 ( .A(ram[2243]), .B(ram[2259]), .S(n4316), .Z(n873) );
  MUX2_X1 U10010 ( .A(n873), .B(n872), .S(n4193), .Z(n874) );
  MUX2_X1 U10011 ( .A(ram[2211]), .B(ram[2227]), .S(n4316), .Z(n875) );
  MUX2_X1 U10012 ( .A(ram[2179]), .B(ram[2195]), .S(n4316), .Z(n876) );
  MUX2_X1 U10013 ( .A(n876), .B(n875), .S(n4193), .Z(n877) );
  MUX2_X1 U10014 ( .A(n877), .B(n874), .S(n4129), .Z(n878) );
  MUX2_X1 U10015 ( .A(ram[2147]), .B(ram[2163]), .S(n4316), .Z(n879) );
  MUX2_X1 U10016 ( .A(ram[2115]), .B(ram[2131]), .S(n4316), .Z(n880) );
  MUX2_X1 U10017 ( .A(n880), .B(n879), .S(n4193), .Z(n881) );
  MUX2_X1 U10018 ( .A(ram[2083]), .B(ram[2099]), .S(n4316), .Z(n882) );
  MUX2_X1 U10019 ( .A(ram[2051]), .B(ram[2067]), .S(n4316), .Z(n883) );
  MUX2_X1 U10020 ( .A(n883), .B(n882), .S(n4193), .Z(n884) );
  MUX2_X1 U10021 ( .A(n884), .B(n881), .S(n4129), .Z(n885) );
  MUX2_X1 U10022 ( .A(n885), .B(n878), .S(n4092), .Z(n886) );
  MUX2_X1 U10023 ( .A(n886), .B(n871), .S(n4078), .Z(n887) );
  MUX2_X1 U10024 ( .A(n887), .B(n856), .S(n4069), .Z(n888) );
  MUX2_X1 U10025 ( .A(n888), .B(n825), .S(n4065), .Z(n889) );
  MUX2_X1 U10026 ( .A(ram[2019]), .B(ram[2035]), .S(n4316), .Z(n890) );
  MUX2_X1 U10027 ( .A(ram[1987]), .B(ram[2003]), .S(n4316), .Z(n891) );
  MUX2_X1 U10028 ( .A(n891), .B(n890), .S(n4193), .Z(n892) );
  MUX2_X1 U10029 ( .A(ram[1955]), .B(ram[1971]), .S(n4316), .Z(n893) );
  MUX2_X1 U10030 ( .A(ram[1923]), .B(ram[1939]), .S(n4316), .Z(n894) );
  MUX2_X1 U10031 ( .A(n894), .B(n893), .S(n4193), .Z(n895) );
  MUX2_X1 U10032 ( .A(n895), .B(n892), .S(n4129), .Z(n896) );
  MUX2_X1 U10033 ( .A(ram[1891]), .B(ram[1907]), .S(n4317), .Z(n897) );
  MUX2_X1 U10034 ( .A(ram[1859]), .B(ram[1875]), .S(n4317), .Z(n898) );
  MUX2_X1 U10035 ( .A(n898), .B(n897), .S(n4193), .Z(n899) );
  MUX2_X1 U10036 ( .A(ram[1827]), .B(ram[1843]), .S(n4317), .Z(n900) );
  MUX2_X1 U10037 ( .A(ram[1795]), .B(ram[1811]), .S(n4317), .Z(n901) );
  MUX2_X1 U10038 ( .A(n901), .B(n900), .S(n4193), .Z(n902) );
  MUX2_X1 U10039 ( .A(n902), .B(n899), .S(n4129), .Z(n903) );
  MUX2_X1 U10040 ( .A(n903), .B(n896), .S(n4092), .Z(n904) );
  MUX2_X1 U10041 ( .A(ram[1763]), .B(ram[1779]), .S(n4317), .Z(n905) );
  MUX2_X1 U10042 ( .A(ram[1731]), .B(ram[1747]), .S(n4317), .Z(n906) );
  MUX2_X1 U10043 ( .A(n906), .B(n905), .S(n4193), .Z(n907) );
  MUX2_X1 U10044 ( .A(ram[1699]), .B(ram[1715]), .S(n4317), .Z(n908) );
  MUX2_X1 U10045 ( .A(ram[1667]), .B(ram[1683]), .S(n4317), .Z(n909) );
  MUX2_X1 U10046 ( .A(n909), .B(n908), .S(n4193), .Z(n910) );
  MUX2_X1 U10047 ( .A(n910), .B(n907), .S(n4129), .Z(n911) );
  MUX2_X1 U10048 ( .A(ram[1635]), .B(ram[1651]), .S(n4317), .Z(n912) );
  MUX2_X1 U10049 ( .A(ram[1603]), .B(ram[1619]), .S(n4317), .Z(n913) );
  MUX2_X1 U10050 ( .A(n913), .B(n912), .S(n4193), .Z(n914) );
  MUX2_X1 U10051 ( .A(ram[1571]), .B(ram[1587]), .S(n4317), .Z(n915) );
  MUX2_X1 U10052 ( .A(ram[1539]), .B(ram[1555]), .S(n4317), .Z(n916) );
  MUX2_X1 U10053 ( .A(n916), .B(n915), .S(n4193), .Z(n917) );
  MUX2_X1 U10054 ( .A(n917), .B(n914), .S(n4129), .Z(n918) );
  MUX2_X1 U10055 ( .A(n918), .B(n911), .S(n4092), .Z(n919) );
  MUX2_X1 U10056 ( .A(n919), .B(n904), .S(n4078), .Z(n920) );
  MUX2_X1 U10057 ( .A(ram[1507]), .B(ram[1523]), .S(n4318), .Z(n921) );
  MUX2_X1 U10058 ( .A(ram[1475]), .B(ram[1491]), .S(n4318), .Z(n922) );
  MUX2_X1 U10059 ( .A(n922), .B(n921), .S(n4194), .Z(n923) );
  MUX2_X1 U10060 ( .A(ram[1443]), .B(ram[1459]), .S(n4318), .Z(n924) );
  MUX2_X1 U10061 ( .A(ram[1411]), .B(ram[1427]), .S(n4318), .Z(n925) );
  MUX2_X1 U10062 ( .A(n925), .B(n924), .S(n4194), .Z(n926) );
  MUX2_X1 U10063 ( .A(n926), .B(n923), .S(n4130), .Z(n927) );
  MUX2_X1 U10064 ( .A(ram[1379]), .B(ram[1395]), .S(n4318), .Z(n928) );
  MUX2_X1 U10065 ( .A(ram[1347]), .B(ram[1363]), .S(n4318), .Z(n929) );
  MUX2_X1 U10066 ( .A(n929), .B(n928), .S(n4194), .Z(n930) );
  MUX2_X1 U10067 ( .A(ram[1315]), .B(ram[1331]), .S(n4318), .Z(n931) );
  MUX2_X1 U10068 ( .A(ram[1283]), .B(ram[1299]), .S(n4318), .Z(n932) );
  MUX2_X1 U10069 ( .A(n932), .B(n931), .S(n4194), .Z(n933) );
  MUX2_X1 U10070 ( .A(n933), .B(n930), .S(n4130), .Z(n934) );
  MUX2_X1 U10071 ( .A(n934), .B(n927), .S(n4092), .Z(n935) );
  MUX2_X1 U10072 ( .A(ram[1251]), .B(ram[1267]), .S(n4318), .Z(n936) );
  MUX2_X1 U10073 ( .A(ram[1219]), .B(ram[1235]), .S(n4318), .Z(n937) );
  MUX2_X1 U10074 ( .A(n937), .B(n936), .S(n4194), .Z(n938) );
  MUX2_X1 U10075 ( .A(ram[1187]), .B(ram[1203]), .S(n4318), .Z(n939) );
  MUX2_X1 U10076 ( .A(ram[1155]), .B(ram[1171]), .S(n4318), .Z(n940) );
  MUX2_X1 U10077 ( .A(n940), .B(n939), .S(n4194), .Z(n941) );
  MUX2_X1 U10078 ( .A(n941), .B(n938), .S(n4130), .Z(n942) );
  MUX2_X1 U10079 ( .A(ram[1123]), .B(ram[1139]), .S(n4319), .Z(n943) );
  MUX2_X1 U10080 ( .A(ram[1091]), .B(ram[1107]), .S(n4319), .Z(n944) );
  MUX2_X1 U10081 ( .A(n944), .B(n943), .S(n4194), .Z(n945) );
  MUX2_X1 U10082 ( .A(ram[1059]), .B(ram[1075]), .S(n4319), .Z(n946) );
  MUX2_X1 U10083 ( .A(ram[1027]), .B(ram[1043]), .S(n4319), .Z(n947) );
  MUX2_X1 U10084 ( .A(n947), .B(n946), .S(n4194), .Z(n948) );
  MUX2_X1 U10085 ( .A(n948), .B(n945), .S(n4130), .Z(n949) );
  MUX2_X1 U10086 ( .A(n949), .B(n942), .S(n4092), .Z(n950) );
  MUX2_X1 U10087 ( .A(n950), .B(n935), .S(n4078), .Z(n951) );
  MUX2_X1 U10088 ( .A(n951), .B(n920), .S(n4069), .Z(n952) );
  MUX2_X1 U10089 ( .A(ram[995]), .B(ram[1011]), .S(n4319), .Z(n953) );
  MUX2_X1 U10090 ( .A(ram[963]), .B(ram[979]), .S(n4319), .Z(n954) );
  MUX2_X1 U10091 ( .A(n954), .B(n953), .S(n4194), .Z(n955) );
  MUX2_X1 U10092 ( .A(ram[931]), .B(ram[947]), .S(n4319), .Z(n956) );
  MUX2_X1 U10093 ( .A(ram[899]), .B(ram[915]), .S(n4319), .Z(n957) );
  MUX2_X1 U10094 ( .A(n957), .B(n956), .S(n4194), .Z(n958) );
  MUX2_X1 U10095 ( .A(n958), .B(n955), .S(n4130), .Z(n959) );
  MUX2_X1 U10096 ( .A(ram[867]), .B(ram[883]), .S(n4319), .Z(n960) );
  MUX2_X1 U10097 ( .A(ram[835]), .B(ram[851]), .S(n4319), .Z(n961) );
  MUX2_X1 U10098 ( .A(n961), .B(n960), .S(n4194), .Z(n962) );
  MUX2_X1 U10099 ( .A(ram[803]), .B(ram[819]), .S(n4319), .Z(n963) );
  MUX2_X1 U10100 ( .A(ram[771]), .B(ram[787]), .S(n4319), .Z(n964) );
  MUX2_X1 U10101 ( .A(n964), .B(n963), .S(n4194), .Z(n965) );
  MUX2_X1 U10102 ( .A(n965), .B(n962), .S(n4130), .Z(n966) );
  MUX2_X1 U10103 ( .A(n966), .B(n959), .S(n4092), .Z(n967) );
  MUX2_X1 U10104 ( .A(ram[739]), .B(ram[755]), .S(n4320), .Z(n968) );
  MUX2_X1 U10105 ( .A(ram[707]), .B(ram[723]), .S(n4320), .Z(n969) );
  MUX2_X1 U10106 ( .A(n969), .B(n968), .S(n4195), .Z(n970) );
  MUX2_X1 U10107 ( .A(ram[675]), .B(ram[691]), .S(n4320), .Z(n971) );
  MUX2_X1 U10108 ( .A(ram[643]), .B(ram[659]), .S(n4320), .Z(n972) );
  MUX2_X1 U10109 ( .A(n972), .B(n971), .S(n4195), .Z(n973) );
  MUX2_X1 U10110 ( .A(n973), .B(n970), .S(n4130), .Z(n974) );
  MUX2_X1 U10111 ( .A(ram[611]), .B(ram[627]), .S(n4320), .Z(n975) );
  MUX2_X1 U10112 ( .A(ram[579]), .B(ram[595]), .S(n4320), .Z(n976) );
  MUX2_X1 U10113 ( .A(n976), .B(n975), .S(n4195), .Z(n977) );
  MUX2_X1 U10114 ( .A(ram[547]), .B(ram[563]), .S(n4320), .Z(n978) );
  MUX2_X1 U10115 ( .A(ram[515]), .B(ram[531]), .S(n4320), .Z(n979) );
  MUX2_X1 U10116 ( .A(n979), .B(n978), .S(n4195), .Z(n980) );
  MUX2_X1 U10117 ( .A(n980), .B(n977), .S(n4130), .Z(n981) );
  MUX2_X1 U10118 ( .A(n981), .B(n974), .S(n4092), .Z(n982) );
  MUX2_X1 U10119 ( .A(n982), .B(n967), .S(n4078), .Z(n983) );
  MUX2_X1 U10120 ( .A(ram[483]), .B(ram[499]), .S(n4320), .Z(n984) );
  MUX2_X1 U10121 ( .A(ram[451]), .B(ram[467]), .S(n4320), .Z(n985) );
  MUX2_X1 U10122 ( .A(n985), .B(n984), .S(n4195), .Z(n986) );
  MUX2_X1 U10123 ( .A(ram[419]), .B(ram[435]), .S(n4320), .Z(n987) );
  MUX2_X1 U10124 ( .A(ram[387]), .B(ram[403]), .S(n4320), .Z(n988) );
  MUX2_X1 U10125 ( .A(n988), .B(n987), .S(n4195), .Z(n989) );
  MUX2_X1 U10126 ( .A(n989), .B(n986), .S(n4130), .Z(n990) );
  MUX2_X1 U10127 ( .A(ram[355]), .B(ram[371]), .S(n4321), .Z(n991) );
  MUX2_X1 U10128 ( .A(ram[323]), .B(ram[339]), .S(n4321), .Z(n992) );
  MUX2_X1 U10129 ( .A(n992), .B(n991), .S(n4195), .Z(n993) );
  MUX2_X1 U10130 ( .A(ram[291]), .B(ram[307]), .S(n4321), .Z(n994) );
  MUX2_X1 U10131 ( .A(ram[259]), .B(ram[275]), .S(n4321), .Z(n995) );
  MUX2_X1 U10132 ( .A(n995), .B(n994), .S(n4195), .Z(n996) );
  MUX2_X1 U10133 ( .A(n996), .B(n993), .S(n4130), .Z(n997) );
  MUX2_X1 U10134 ( .A(n997), .B(n990), .S(n4092), .Z(n998) );
  MUX2_X1 U10135 ( .A(ram[227]), .B(ram[243]), .S(n4321), .Z(n999) );
  MUX2_X1 U10136 ( .A(ram[195]), .B(ram[211]), .S(n4321), .Z(n1000) );
  MUX2_X1 U10137 ( .A(n1000), .B(n999), .S(n4195), .Z(n1001) );
  MUX2_X1 U10138 ( .A(ram[163]), .B(ram[179]), .S(n4321), .Z(n1002) );
  MUX2_X1 U10139 ( .A(ram[131]), .B(ram[147]), .S(n4321), .Z(n1003) );
  MUX2_X1 U10140 ( .A(n1003), .B(n1002), .S(n4195), .Z(n1004) );
  MUX2_X1 U10141 ( .A(n1004), .B(n1001), .S(n4130), .Z(n1005) );
  MUX2_X1 U10142 ( .A(ram[99]), .B(ram[115]), .S(n4321), .Z(n1006) );
  MUX2_X1 U10143 ( .A(ram[67]), .B(ram[83]), .S(n4321), .Z(n1007) );
  MUX2_X1 U10144 ( .A(n1007), .B(n1006), .S(n4195), .Z(n1008) );
  MUX2_X1 U10145 ( .A(ram[35]), .B(ram[51]), .S(n4321), .Z(n1009) );
  MUX2_X1 U10146 ( .A(ram[3]), .B(ram[19]), .S(n4321), .Z(n1010) );
  MUX2_X1 U10147 ( .A(n1010), .B(n1009), .S(n4195), .Z(n1011) );
  MUX2_X1 U10148 ( .A(n1011), .B(n1008), .S(n4130), .Z(n1012) );
  MUX2_X1 U10149 ( .A(n1012), .B(n1005), .S(n4092), .Z(n1013) );
  MUX2_X1 U10150 ( .A(n1013), .B(n998), .S(n4078), .Z(n1014) );
  MUX2_X1 U10151 ( .A(n1014), .B(n983), .S(n4069), .Z(n1015) );
  MUX2_X1 U10152 ( .A(n1015), .B(n952), .S(n4065), .Z(n1016) );
  MUX2_X1 U10153 ( .A(n1016), .B(n889), .S(mem_access_addr[9]), .Z(N298) );
  MUX2_X1 U10154 ( .A(ram[4068]), .B(ram[4084]), .S(n4322), .Z(n1017) );
  MUX2_X1 U10155 ( .A(ram[4036]), .B(ram[4052]), .S(n4322), .Z(n1018) );
  MUX2_X1 U10156 ( .A(n1018), .B(n1017), .S(n4196), .Z(n1019) );
  MUX2_X1 U10157 ( .A(ram[4004]), .B(ram[4020]), .S(n4322), .Z(n1020) );
  MUX2_X1 U10158 ( .A(ram[3972]), .B(ram[3988]), .S(n4322), .Z(n1021) );
  MUX2_X1 U10159 ( .A(n1021), .B(n1020), .S(n4196), .Z(n1022) );
  MUX2_X1 U10160 ( .A(n1022), .B(n1019), .S(n4131), .Z(n1023) );
  MUX2_X1 U10161 ( .A(ram[3940]), .B(ram[3956]), .S(n4322), .Z(n1024) );
  MUX2_X1 U10162 ( .A(ram[3908]), .B(ram[3924]), .S(n4322), .Z(n1025) );
  MUX2_X1 U10163 ( .A(n1025), .B(n1024), .S(n4196), .Z(n1026) );
  MUX2_X1 U10164 ( .A(ram[3876]), .B(ram[3892]), .S(n4322), .Z(n1027) );
  MUX2_X1 U10165 ( .A(ram[3844]), .B(ram[3860]), .S(n4322), .Z(n1028) );
  MUX2_X1 U10166 ( .A(n1028), .B(n1027), .S(n4196), .Z(n1029) );
  MUX2_X1 U10167 ( .A(n1029), .B(n1026), .S(n4131), .Z(n1030) );
  MUX2_X1 U10168 ( .A(n1030), .B(n1023), .S(n4093), .Z(n1031) );
  MUX2_X1 U10169 ( .A(ram[3812]), .B(ram[3828]), .S(n4322), .Z(n1032) );
  MUX2_X1 U10170 ( .A(ram[3780]), .B(ram[3796]), .S(n4322), .Z(n1033) );
  MUX2_X1 U10171 ( .A(n1033), .B(n1032), .S(n4196), .Z(n1034) );
  MUX2_X1 U10172 ( .A(ram[3748]), .B(ram[3764]), .S(n4322), .Z(n1035) );
  MUX2_X1 U10173 ( .A(ram[3716]), .B(ram[3732]), .S(n4322), .Z(n1036) );
  MUX2_X1 U10174 ( .A(n1036), .B(n1035), .S(n4196), .Z(n1037) );
  MUX2_X1 U10175 ( .A(n1037), .B(n1034), .S(n4131), .Z(n1038) );
  MUX2_X1 U10176 ( .A(ram[3684]), .B(ram[3700]), .S(n4323), .Z(n1039) );
  MUX2_X1 U10177 ( .A(ram[3652]), .B(ram[3668]), .S(n4323), .Z(n1040) );
  MUX2_X1 U10178 ( .A(n1040), .B(n1039), .S(n4196), .Z(n1041) );
  MUX2_X1 U10179 ( .A(ram[3620]), .B(ram[3636]), .S(n4323), .Z(n1042) );
  MUX2_X1 U10180 ( .A(ram[3588]), .B(ram[3604]), .S(n4323), .Z(n1043) );
  MUX2_X1 U10181 ( .A(n1043), .B(n1042), .S(n4196), .Z(n1044) );
  MUX2_X1 U10182 ( .A(n1044), .B(n1041), .S(n4131), .Z(n1045) );
  MUX2_X1 U10183 ( .A(n1045), .B(n1038), .S(n4093), .Z(n1046) );
  MUX2_X1 U10184 ( .A(n1046), .B(n1031), .S(n4079), .Z(n1047) );
  MUX2_X1 U10185 ( .A(ram[3556]), .B(ram[3572]), .S(n4323), .Z(n1048) );
  MUX2_X1 U10186 ( .A(ram[3524]), .B(ram[3540]), .S(n4323), .Z(n1049) );
  MUX2_X1 U10187 ( .A(n1049), .B(n1048), .S(n4196), .Z(n1050) );
  MUX2_X1 U10188 ( .A(ram[3492]), .B(ram[3508]), .S(n4323), .Z(n1051) );
  MUX2_X1 U10189 ( .A(ram[3460]), .B(ram[3476]), .S(n4323), .Z(n1052) );
  MUX2_X1 U10190 ( .A(n1052), .B(n1051), .S(n4196), .Z(n1053) );
  MUX2_X1 U10191 ( .A(n1053), .B(n1050), .S(n4131), .Z(n1054) );
  MUX2_X1 U10192 ( .A(ram[3428]), .B(ram[3444]), .S(n4323), .Z(n1055) );
  MUX2_X1 U10193 ( .A(ram[3396]), .B(ram[3412]), .S(n4323), .Z(n1056) );
  MUX2_X1 U10194 ( .A(n1056), .B(n1055), .S(n4196), .Z(n1057) );
  MUX2_X1 U10195 ( .A(ram[3364]), .B(ram[3380]), .S(n4323), .Z(n1058) );
  MUX2_X1 U10196 ( .A(ram[3332]), .B(ram[3348]), .S(n4323), .Z(n1059) );
  MUX2_X1 U10197 ( .A(n1059), .B(n1058), .S(n4196), .Z(n1060) );
  MUX2_X1 U10198 ( .A(n1060), .B(n1057), .S(n4131), .Z(n1061) );
  MUX2_X1 U10199 ( .A(n1061), .B(n1054), .S(n4093), .Z(n1062) );
  MUX2_X1 U10200 ( .A(ram[3300]), .B(ram[3316]), .S(n4324), .Z(n1063) );
  MUX2_X1 U10201 ( .A(ram[3268]), .B(ram[3284]), .S(n4324), .Z(n1064) );
  MUX2_X1 U10202 ( .A(n1064), .B(n1063), .S(n4197), .Z(n1065) );
  MUX2_X1 U10203 ( .A(ram[3236]), .B(ram[3252]), .S(n4324), .Z(n1066) );
  MUX2_X1 U10204 ( .A(ram[3204]), .B(ram[3220]), .S(n4324), .Z(n1067) );
  MUX2_X1 U10205 ( .A(n1067), .B(n1066), .S(n4197), .Z(n1068) );
  MUX2_X1 U10206 ( .A(n1068), .B(n1065), .S(n4131), .Z(n1069) );
  MUX2_X1 U10207 ( .A(ram[3172]), .B(ram[3188]), .S(n4324), .Z(n1070) );
  MUX2_X1 U10208 ( .A(ram[3140]), .B(ram[3156]), .S(n4324), .Z(n1071) );
  MUX2_X1 U10209 ( .A(n1071), .B(n1070), .S(n4197), .Z(n1072) );
  MUX2_X1 U10210 ( .A(ram[3108]), .B(ram[3124]), .S(n4324), .Z(n1073) );
  MUX2_X1 U10211 ( .A(ram[3076]), .B(ram[3092]), .S(n4324), .Z(n1074) );
  MUX2_X1 U10212 ( .A(n1074), .B(n1073), .S(n4197), .Z(n1075) );
  MUX2_X1 U10213 ( .A(n1075), .B(n1072), .S(n4131), .Z(n1076) );
  MUX2_X1 U10214 ( .A(n1076), .B(n1069), .S(n4093), .Z(n1077) );
  MUX2_X1 U10215 ( .A(n1077), .B(n1062), .S(n4079), .Z(n1078) );
  MUX2_X1 U10216 ( .A(n1078), .B(n1047), .S(n4070), .Z(n1079) );
  MUX2_X1 U10217 ( .A(ram[3044]), .B(ram[3060]), .S(n4324), .Z(n1080) );
  MUX2_X1 U10218 ( .A(ram[3012]), .B(ram[3028]), .S(n4324), .Z(n1081) );
  MUX2_X1 U10219 ( .A(n1081), .B(n1080), .S(n4197), .Z(n1082) );
  MUX2_X1 U10220 ( .A(ram[2980]), .B(ram[2996]), .S(n4324), .Z(n1083) );
  MUX2_X1 U10221 ( .A(ram[2948]), .B(ram[2964]), .S(n4324), .Z(n1084) );
  MUX2_X1 U10222 ( .A(n1084), .B(n1083), .S(n4197), .Z(n1085) );
  MUX2_X1 U10223 ( .A(n1085), .B(n1082), .S(n4131), .Z(n1086) );
  MUX2_X1 U10224 ( .A(ram[2916]), .B(ram[2932]), .S(n4325), .Z(n1087) );
  MUX2_X1 U10225 ( .A(ram[2884]), .B(ram[2900]), .S(n4325), .Z(n1088) );
  MUX2_X1 U10226 ( .A(n1088), .B(n1087), .S(n4197), .Z(n1089) );
  MUX2_X1 U10227 ( .A(ram[2852]), .B(ram[2868]), .S(n4325), .Z(n1090) );
  MUX2_X1 U10228 ( .A(ram[2820]), .B(ram[2836]), .S(n4325), .Z(n1091) );
  MUX2_X1 U10229 ( .A(n1091), .B(n1090), .S(n4197), .Z(n1092) );
  MUX2_X1 U10230 ( .A(n1092), .B(n1089), .S(n4131), .Z(n1093) );
  MUX2_X1 U10231 ( .A(n1093), .B(n1086), .S(n4093), .Z(n1094) );
  MUX2_X1 U10232 ( .A(ram[2788]), .B(ram[2804]), .S(n4325), .Z(n1095) );
  MUX2_X1 U10233 ( .A(ram[2756]), .B(ram[2772]), .S(n4325), .Z(n1096) );
  MUX2_X1 U10234 ( .A(n1096), .B(n1095), .S(n4197), .Z(n1097) );
  MUX2_X1 U10235 ( .A(ram[2724]), .B(ram[2740]), .S(n4325), .Z(n1098) );
  MUX2_X1 U10236 ( .A(ram[2692]), .B(ram[2708]), .S(n4325), .Z(n1099) );
  MUX2_X1 U10237 ( .A(n1099), .B(n1098), .S(n4197), .Z(n1100) );
  MUX2_X1 U10238 ( .A(n1100), .B(n1097), .S(n4131), .Z(n1101) );
  MUX2_X1 U10239 ( .A(ram[2660]), .B(ram[2676]), .S(n4325), .Z(n1102) );
  MUX2_X1 U10240 ( .A(ram[2628]), .B(ram[2644]), .S(n4325), .Z(n1103) );
  MUX2_X1 U10241 ( .A(n1103), .B(n1102), .S(n4197), .Z(n1104) );
  MUX2_X1 U10242 ( .A(ram[2596]), .B(ram[2612]), .S(n4325), .Z(n1105) );
  MUX2_X1 U10243 ( .A(ram[2564]), .B(ram[2580]), .S(n4325), .Z(n1106) );
  MUX2_X1 U10244 ( .A(n1106), .B(n1105), .S(n4197), .Z(n1107) );
  MUX2_X1 U10245 ( .A(n1107), .B(n1104), .S(n4131), .Z(n1108) );
  MUX2_X1 U10246 ( .A(n1108), .B(n1101), .S(n4093), .Z(n1109) );
  MUX2_X1 U10247 ( .A(n1109), .B(n1094), .S(n4079), .Z(n1110) );
  MUX2_X1 U10248 ( .A(ram[2532]), .B(ram[2548]), .S(n4326), .Z(n1111) );
  MUX2_X1 U10249 ( .A(ram[2500]), .B(ram[2516]), .S(n4326), .Z(n1112) );
  MUX2_X1 U10250 ( .A(n1112), .B(n1111), .S(n4198), .Z(n1113) );
  MUX2_X1 U10251 ( .A(ram[2468]), .B(ram[2484]), .S(n4326), .Z(n1114) );
  MUX2_X1 U10252 ( .A(ram[2436]), .B(ram[2452]), .S(n4326), .Z(n1115) );
  MUX2_X1 U10253 ( .A(n1115), .B(n1114), .S(n4198), .Z(n1116) );
  MUX2_X1 U10254 ( .A(n1116), .B(n1113), .S(n4132), .Z(n1117) );
  MUX2_X1 U10255 ( .A(ram[2404]), .B(ram[2420]), .S(n4326), .Z(n1118) );
  MUX2_X1 U10256 ( .A(ram[2372]), .B(ram[2388]), .S(n4326), .Z(n1119) );
  MUX2_X1 U10257 ( .A(n1119), .B(n1118), .S(n4198), .Z(n1120) );
  MUX2_X1 U10258 ( .A(ram[2340]), .B(ram[2356]), .S(n4326), .Z(n1121) );
  MUX2_X1 U10259 ( .A(ram[2308]), .B(ram[2324]), .S(n4326), .Z(n1122) );
  MUX2_X1 U10260 ( .A(n1122), .B(n1121), .S(n4198), .Z(n1123) );
  MUX2_X1 U10261 ( .A(n1123), .B(n1120), .S(n4132), .Z(n1124) );
  MUX2_X1 U10262 ( .A(n1124), .B(n1117), .S(n4093), .Z(n1125) );
  MUX2_X1 U10263 ( .A(ram[2276]), .B(ram[2292]), .S(n4326), .Z(n1126) );
  MUX2_X1 U10264 ( .A(ram[2244]), .B(ram[2260]), .S(n4326), .Z(n1127) );
  MUX2_X1 U10265 ( .A(n1127), .B(n1126), .S(n4198), .Z(n1128) );
  MUX2_X1 U10266 ( .A(ram[2212]), .B(ram[2228]), .S(n4326), .Z(n1129) );
  MUX2_X1 U10267 ( .A(ram[2180]), .B(ram[2196]), .S(n4326), .Z(n1130) );
  MUX2_X1 U10268 ( .A(n1130), .B(n1129), .S(n4198), .Z(n1131) );
  MUX2_X1 U10269 ( .A(n1131), .B(n1128), .S(n4132), .Z(n1132) );
  MUX2_X1 U10270 ( .A(ram[2148]), .B(ram[2164]), .S(n4327), .Z(n1133) );
  MUX2_X1 U10271 ( .A(ram[2116]), .B(ram[2132]), .S(n4327), .Z(n1134) );
  MUX2_X1 U10272 ( .A(n1134), .B(n1133), .S(n4198), .Z(n1135) );
  MUX2_X1 U10273 ( .A(ram[2084]), .B(ram[2100]), .S(n4327), .Z(n1136) );
  MUX2_X1 U10274 ( .A(ram[2052]), .B(ram[2068]), .S(n4327), .Z(n1137) );
  MUX2_X1 U10275 ( .A(n1137), .B(n1136), .S(n4198), .Z(n1138) );
  MUX2_X1 U10276 ( .A(n1138), .B(n1135), .S(n4132), .Z(n1139) );
  MUX2_X1 U10277 ( .A(n1139), .B(n1132), .S(n4093), .Z(n1140) );
  MUX2_X1 U10278 ( .A(n1140), .B(n1125), .S(n4079), .Z(n1141) );
  MUX2_X1 U10279 ( .A(n1141), .B(n1110), .S(n4070), .Z(n1142) );
  MUX2_X1 U10280 ( .A(n1142), .B(n1079), .S(n4066), .Z(n1143) );
  MUX2_X1 U10281 ( .A(ram[2020]), .B(ram[2036]), .S(n4327), .Z(n1144) );
  MUX2_X1 U10282 ( .A(ram[1988]), .B(ram[2004]), .S(n4327), .Z(n1145) );
  MUX2_X1 U10283 ( .A(n1145), .B(n1144), .S(n4198), .Z(n1146) );
  MUX2_X1 U10284 ( .A(ram[1956]), .B(ram[1972]), .S(n4327), .Z(n1147) );
  MUX2_X1 U10285 ( .A(ram[1924]), .B(ram[1940]), .S(n4327), .Z(n1148) );
  MUX2_X1 U10286 ( .A(n1148), .B(n1147), .S(n4198), .Z(n1149) );
  MUX2_X1 U10287 ( .A(n1149), .B(n1146), .S(n4132), .Z(n1150) );
  MUX2_X1 U10288 ( .A(ram[1892]), .B(ram[1908]), .S(n4327), .Z(n1151) );
  MUX2_X1 U10289 ( .A(ram[1860]), .B(ram[1876]), .S(n4327), .Z(n1152) );
  MUX2_X1 U10290 ( .A(n1152), .B(n1151), .S(n4198), .Z(n1153) );
  MUX2_X1 U10291 ( .A(ram[1828]), .B(ram[1844]), .S(n4327), .Z(n1154) );
  MUX2_X1 U10292 ( .A(ram[1796]), .B(ram[1812]), .S(n4327), .Z(n1155) );
  MUX2_X1 U10293 ( .A(n1155), .B(n1154), .S(n4198), .Z(n1156) );
  MUX2_X1 U10294 ( .A(n1156), .B(n1153), .S(n4132), .Z(n1157) );
  MUX2_X1 U10295 ( .A(n1157), .B(n1150), .S(n4093), .Z(n1158) );
  MUX2_X1 U10296 ( .A(ram[1764]), .B(ram[1780]), .S(n4328), .Z(n1159) );
  MUX2_X1 U10297 ( .A(ram[1732]), .B(ram[1748]), .S(n4328), .Z(n1160) );
  MUX2_X1 U10298 ( .A(n1160), .B(n1159), .S(n4199), .Z(n1161) );
  MUX2_X1 U10299 ( .A(ram[1700]), .B(ram[1716]), .S(n4328), .Z(n1162) );
  MUX2_X1 U10300 ( .A(ram[1668]), .B(ram[1684]), .S(n4328), .Z(n1163) );
  MUX2_X1 U10301 ( .A(n1163), .B(n1162), .S(n4199), .Z(n1164) );
  MUX2_X1 U10302 ( .A(n1164), .B(n1161), .S(n4132), .Z(n1165) );
  MUX2_X1 U10303 ( .A(ram[1636]), .B(ram[1652]), .S(n4328), .Z(n1166) );
  MUX2_X1 U10304 ( .A(ram[1604]), .B(ram[1620]), .S(n4328), .Z(n1167) );
  MUX2_X1 U10305 ( .A(n1167), .B(n1166), .S(n4199), .Z(n1168) );
  MUX2_X1 U10306 ( .A(ram[1572]), .B(ram[1588]), .S(n4328), .Z(n1169) );
  MUX2_X1 U10307 ( .A(ram[1540]), .B(ram[1556]), .S(n4328), .Z(n1170) );
  MUX2_X1 U10308 ( .A(n1170), .B(n1169), .S(n4199), .Z(n1171) );
  MUX2_X1 U10309 ( .A(n1171), .B(n1168), .S(n4132), .Z(n1172) );
  MUX2_X1 U10310 ( .A(n1172), .B(n1165), .S(n4093), .Z(n1173) );
  MUX2_X1 U10311 ( .A(n1173), .B(n1158), .S(n4079), .Z(n1174) );
  MUX2_X1 U10312 ( .A(ram[1508]), .B(ram[1524]), .S(n4328), .Z(n1175) );
  MUX2_X1 U10313 ( .A(ram[1476]), .B(ram[1492]), .S(n4328), .Z(n1176) );
  MUX2_X1 U10314 ( .A(n1176), .B(n1175), .S(n4199), .Z(n1177) );
  MUX2_X1 U10315 ( .A(ram[1444]), .B(ram[1460]), .S(n4328), .Z(n1178) );
  MUX2_X1 U10316 ( .A(ram[1412]), .B(ram[1428]), .S(n4328), .Z(n1179) );
  MUX2_X1 U10317 ( .A(n1179), .B(n1178), .S(n4199), .Z(n1180) );
  MUX2_X1 U10318 ( .A(n1180), .B(n1177), .S(n4132), .Z(n1181) );
  MUX2_X1 U10319 ( .A(ram[1380]), .B(ram[1396]), .S(n4329), .Z(n1182) );
  MUX2_X1 U10320 ( .A(ram[1348]), .B(ram[1364]), .S(n4329), .Z(n1183) );
  MUX2_X1 U10321 ( .A(n1183), .B(n1182), .S(n4199), .Z(n1184) );
  MUX2_X1 U10322 ( .A(ram[1316]), .B(ram[1332]), .S(n4329), .Z(n1185) );
  MUX2_X1 U10323 ( .A(ram[1284]), .B(ram[1300]), .S(n4329), .Z(n1186) );
  MUX2_X1 U10324 ( .A(n1186), .B(n1185), .S(n4199), .Z(n1187) );
  MUX2_X1 U10325 ( .A(n1187), .B(n1184), .S(n4132), .Z(n1188) );
  MUX2_X1 U10326 ( .A(n1188), .B(n1181), .S(n4093), .Z(n1189) );
  MUX2_X1 U10327 ( .A(ram[1252]), .B(ram[1268]), .S(n4329), .Z(n1190) );
  MUX2_X1 U10328 ( .A(ram[1220]), .B(ram[1236]), .S(n4329), .Z(n1191) );
  MUX2_X1 U10329 ( .A(n1191), .B(n1190), .S(n4199), .Z(n1192) );
  MUX2_X1 U10330 ( .A(ram[1188]), .B(ram[1204]), .S(n4329), .Z(n1193) );
  MUX2_X1 U10331 ( .A(ram[1156]), .B(ram[1172]), .S(n4329), .Z(n1194) );
  MUX2_X1 U10332 ( .A(n1194), .B(n1193), .S(n4199), .Z(n1195) );
  MUX2_X1 U10333 ( .A(n1195), .B(n1192), .S(n4132), .Z(n1196) );
  MUX2_X1 U10334 ( .A(ram[1124]), .B(ram[1140]), .S(n4329), .Z(n1197) );
  MUX2_X1 U10335 ( .A(ram[1092]), .B(ram[1108]), .S(n4329), .Z(n1198) );
  MUX2_X1 U10336 ( .A(n1198), .B(n1197), .S(n4199), .Z(n1199) );
  MUX2_X1 U10337 ( .A(ram[1060]), .B(ram[1076]), .S(n4329), .Z(n1200) );
  MUX2_X1 U10338 ( .A(ram[1028]), .B(ram[1044]), .S(n4329), .Z(n1201) );
  MUX2_X1 U10339 ( .A(n1201), .B(n1200), .S(n4199), .Z(n1202) );
  MUX2_X1 U10340 ( .A(n1202), .B(n1199), .S(n4132), .Z(n1203) );
  MUX2_X1 U10341 ( .A(n1203), .B(n1196), .S(n4093), .Z(n1204) );
  MUX2_X1 U10342 ( .A(n1204), .B(n1189), .S(n4079), .Z(n1205) );
  MUX2_X1 U10343 ( .A(n1205), .B(n1174), .S(n4070), .Z(n1206) );
  MUX2_X1 U10344 ( .A(ram[996]), .B(ram[1012]), .S(n4330), .Z(n1207) );
  MUX2_X1 U10345 ( .A(ram[964]), .B(ram[980]), .S(n4330), .Z(n1208) );
  MUX2_X1 U10346 ( .A(n1208), .B(n1207), .S(n4200), .Z(n1209) );
  MUX2_X1 U10347 ( .A(ram[932]), .B(ram[948]), .S(n4330), .Z(n1210) );
  MUX2_X1 U10348 ( .A(ram[900]), .B(ram[916]), .S(n4330), .Z(n1211) );
  MUX2_X1 U10349 ( .A(n1211), .B(n1210), .S(n4200), .Z(n1212) );
  MUX2_X1 U10350 ( .A(n1212), .B(n1209), .S(n4133), .Z(n1213) );
  MUX2_X1 U10351 ( .A(ram[868]), .B(ram[884]), .S(n4330), .Z(n1214) );
  MUX2_X1 U10352 ( .A(ram[836]), .B(ram[852]), .S(n4330), .Z(n1215) );
  MUX2_X1 U10353 ( .A(n1215), .B(n1214), .S(n4200), .Z(n1216) );
  MUX2_X1 U10354 ( .A(ram[804]), .B(ram[820]), .S(n4330), .Z(n1217) );
  MUX2_X1 U10355 ( .A(ram[772]), .B(ram[788]), .S(n4330), .Z(n1218) );
  MUX2_X1 U10356 ( .A(n1218), .B(n1217), .S(n4200), .Z(n1219) );
  MUX2_X1 U10357 ( .A(n1219), .B(n1216), .S(n4133), .Z(n1220) );
  MUX2_X1 U10358 ( .A(n1220), .B(n1213), .S(n4094), .Z(n1221) );
  MUX2_X1 U10359 ( .A(ram[740]), .B(ram[756]), .S(n4330), .Z(n1222) );
  MUX2_X1 U10360 ( .A(ram[708]), .B(ram[724]), .S(n4330), .Z(n1223) );
  MUX2_X1 U10361 ( .A(n1223), .B(n1222), .S(n4200), .Z(n1224) );
  MUX2_X1 U10362 ( .A(ram[676]), .B(ram[692]), .S(n4330), .Z(n1225) );
  MUX2_X1 U10363 ( .A(ram[644]), .B(ram[660]), .S(n4330), .Z(n1226) );
  MUX2_X1 U10364 ( .A(n1226), .B(n1225), .S(n4200), .Z(n1227) );
  MUX2_X1 U10365 ( .A(n1227), .B(n1224), .S(n4133), .Z(n1228) );
  MUX2_X1 U10366 ( .A(ram[612]), .B(ram[628]), .S(n4331), .Z(n1229) );
  MUX2_X1 U10367 ( .A(ram[580]), .B(ram[596]), .S(n4331), .Z(n1230) );
  MUX2_X1 U10368 ( .A(n1230), .B(n1229), .S(n4200), .Z(n1231) );
  MUX2_X1 U10369 ( .A(ram[548]), .B(ram[564]), .S(n4331), .Z(n1232) );
  MUX2_X1 U10370 ( .A(ram[516]), .B(ram[532]), .S(n4331), .Z(n1233) );
  MUX2_X1 U10371 ( .A(n1233), .B(n1232), .S(n4200), .Z(n1234) );
  MUX2_X1 U10372 ( .A(n1234), .B(n1231), .S(n4133), .Z(n1235) );
  MUX2_X1 U10373 ( .A(n1235), .B(n1228), .S(n4094), .Z(n1236) );
  MUX2_X1 U10374 ( .A(n1236), .B(n1221), .S(n4079), .Z(n1237) );
  MUX2_X1 U10375 ( .A(ram[484]), .B(ram[500]), .S(n4331), .Z(n1238) );
  MUX2_X1 U10376 ( .A(ram[452]), .B(ram[468]), .S(n4331), .Z(n1239) );
  MUX2_X1 U10377 ( .A(n1239), .B(n1238), .S(n4200), .Z(n1240) );
  MUX2_X1 U10378 ( .A(ram[420]), .B(ram[436]), .S(n4331), .Z(n1241) );
  MUX2_X1 U10379 ( .A(ram[388]), .B(ram[404]), .S(n4331), .Z(n1242) );
  MUX2_X1 U10380 ( .A(n1242), .B(n1241), .S(n4200), .Z(n1243) );
  MUX2_X1 U10381 ( .A(n1243), .B(n1240), .S(n4133), .Z(n1244) );
  MUX2_X1 U10382 ( .A(ram[356]), .B(ram[372]), .S(n4331), .Z(n1245) );
  MUX2_X1 U10383 ( .A(ram[324]), .B(ram[340]), .S(n4331), .Z(n1246) );
  MUX2_X1 U10384 ( .A(n1246), .B(n1245), .S(n4200), .Z(n1247) );
  MUX2_X1 U10385 ( .A(ram[292]), .B(ram[308]), .S(n4331), .Z(n1248) );
  MUX2_X1 U10386 ( .A(ram[260]), .B(ram[276]), .S(n4331), .Z(n1249) );
  MUX2_X1 U10387 ( .A(n1249), .B(n1248), .S(n4200), .Z(n1250) );
  MUX2_X1 U10388 ( .A(n1250), .B(n1247), .S(n4133), .Z(n1251) );
  MUX2_X1 U10389 ( .A(n1251), .B(n1244), .S(n4094), .Z(n1252) );
  MUX2_X1 U10390 ( .A(ram[228]), .B(ram[244]), .S(n4332), .Z(n1253) );
  MUX2_X1 U10391 ( .A(ram[196]), .B(ram[212]), .S(n4332), .Z(n1254) );
  MUX2_X1 U10392 ( .A(n1254), .B(n1253), .S(n4201), .Z(n1255) );
  MUX2_X1 U10393 ( .A(ram[164]), .B(ram[180]), .S(n4332), .Z(n1256) );
  MUX2_X1 U10394 ( .A(ram[132]), .B(ram[148]), .S(n4332), .Z(n1257) );
  MUX2_X1 U10395 ( .A(n1257), .B(n1256), .S(n4201), .Z(n1258) );
  MUX2_X1 U10396 ( .A(n1258), .B(n1255), .S(n4133), .Z(n1259) );
  MUX2_X1 U10397 ( .A(ram[100]), .B(ram[116]), .S(n4332), .Z(n1260) );
  MUX2_X1 U10398 ( .A(ram[68]), .B(ram[84]), .S(n4332), .Z(n1261) );
  MUX2_X1 U10399 ( .A(n1261), .B(n1260), .S(n4201), .Z(n1262) );
  MUX2_X1 U10400 ( .A(ram[36]), .B(ram[52]), .S(n4332), .Z(n1263) );
  MUX2_X1 U10401 ( .A(ram[4]), .B(ram[20]), .S(n4332), .Z(n1264) );
  MUX2_X1 U10402 ( .A(n1264), .B(n1263), .S(n4201), .Z(n1265) );
  MUX2_X1 U10403 ( .A(n1265), .B(n1262), .S(n4133), .Z(n1266) );
  MUX2_X1 U10404 ( .A(n1266), .B(n1259), .S(n4094), .Z(n1267) );
  MUX2_X1 U10405 ( .A(n1267), .B(n1252), .S(n4079), .Z(n1268) );
  MUX2_X1 U10406 ( .A(n1268), .B(n1237), .S(n4070), .Z(n1269) );
  MUX2_X1 U10407 ( .A(n1269), .B(n1206), .S(n4066), .Z(n1270) );
  MUX2_X1 U10408 ( .A(n1270), .B(n1143), .S(mem_access_addr[9]), .Z(N297) );
  MUX2_X1 U10409 ( .A(ram[4069]), .B(ram[4085]), .S(n4332), .Z(n1271) );
  MUX2_X1 U10410 ( .A(ram[4037]), .B(ram[4053]), .S(n4332), .Z(n1272) );
  MUX2_X1 U10411 ( .A(n1272), .B(n1271), .S(n4201), .Z(n1273) );
  MUX2_X1 U10412 ( .A(ram[4005]), .B(ram[4021]), .S(n4332), .Z(n1274) );
  MUX2_X1 U10413 ( .A(ram[3973]), .B(ram[3989]), .S(n4332), .Z(n1275) );
  MUX2_X1 U10414 ( .A(n1275), .B(n1274), .S(n4201), .Z(n1276) );
  MUX2_X1 U10415 ( .A(n1276), .B(n1273), .S(n4133), .Z(n1277) );
  MUX2_X1 U10416 ( .A(ram[3941]), .B(ram[3957]), .S(n4333), .Z(n1278) );
  MUX2_X1 U10417 ( .A(ram[3909]), .B(ram[3925]), .S(n4333), .Z(n1279) );
  MUX2_X1 U10418 ( .A(n1279), .B(n1278), .S(n4201), .Z(n1280) );
  MUX2_X1 U10419 ( .A(ram[3877]), .B(ram[3893]), .S(n4333), .Z(n1281) );
  MUX2_X1 U10420 ( .A(ram[3845]), .B(ram[3861]), .S(n4333), .Z(n1282) );
  MUX2_X1 U10421 ( .A(n1282), .B(n1281), .S(n4201), .Z(n1283) );
  MUX2_X1 U10422 ( .A(n1283), .B(n1280), .S(n4133), .Z(n1284) );
  MUX2_X1 U10423 ( .A(n1284), .B(n1277), .S(n4094), .Z(n1285) );
  MUX2_X1 U10424 ( .A(ram[3813]), .B(ram[3829]), .S(n4333), .Z(n1286) );
  MUX2_X1 U10425 ( .A(ram[3781]), .B(ram[3797]), .S(n4333), .Z(n1287) );
  MUX2_X1 U10426 ( .A(n1287), .B(n1286), .S(n4201), .Z(n1288) );
  MUX2_X1 U10427 ( .A(ram[3749]), .B(ram[3765]), .S(n4333), .Z(n1289) );
  MUX2_X1 U10428 ( .A(ram[3717]), .B(ram[3733]), .S(n4333), .Z(n1290) );
  MUX2_X1 U10429 ( .A(n1290), .B(n1289), .S(n4201), .Z(n1291) );
  MUX2_X1 U10430 ( .A(n1291), .B(n1288), .S(n4133), .Z(n1292) );
  MUX2_X1 U10431 ( .A(ram[3685]), .B(ram[3701]), .S(n4333), .Z(n1293) );
  MUX2_X1 U10432 ( .A(ram[3653]), .B(ram[3669]), .S(n4333), .Z(n1294) );
  MUX2_X1 U10433 ( .A(n1294), .B(n1293), .S(n4201), .Z(n1295) );
  MUX2_X1 U10434 ( .A(ram[3621]), .B(ram[3637]), .S(n4333), .Z(n1296) );
  MUX2_X1 U10435 ( .A(ram[3589]), .B(ram[3605]), .S(n4333), .Z(n1297) );
  MUX2_X1 U10436 ( .A(n1297), .B(n1296), .S(n4201), .Z(n1298) );
  MUX2_X1 U10437 ( .A(n1298), .B(n1295), .S(n4133), .Z(n1299) );
  MUX2_X1 U10438 ( .A(n1299), .B(n1292), .S(n4094), .Z(n1300) );
  MUX2_X1 U10439 ( .A(n1300), .B(n1285), .S(n4079), .Z(n1301) );
  MUX2_X1 U10440 ( .A(ram[3557]), .B(ram[3573]), .S(n4334), .Z(n1302) );
  MUX2_X1 U10441 ( .A(ram[3525]), .B(ram[3541]), .S(n4334), .Z(n1303) );
  MUX2_X1 U10442 ( .A(n1303), .B(n1302), .S(n4202), .Z(n1304) );
  MUX2_X1 U10443 ( .A(ram[3493]), .B(ram[3509]), .S(n4334), .Z(n1305) );
  MUX2_X1 U10444 ( .A(ram[3461]), .B(ram[3477]), .S(n4334), .Z(n1306) );
  MUX2_X1 U10445 ( .A(n1306), .B(n1305), .S(n4202), .Z(n1307) );
  MUX2_X1 U10446 ( .A(n1307), .B(n1304), .S(n4134), .Z(n1308) );
  MUX2_X1 U10447 ( .A(ram[3429]), .B(ram[3445]), .S(n4334), .Z(n1309) );
  MUX2_X1 U10448 ( .A(ram[3397]), .B(ram[3413]), .S(n4334), .Z(n1310) );
  MUX2_X1 U10449 ( .A(n1310), .B(n1309), .S(n4202), .Z(n1311) );
  MUX2_X1 U10450 ( .A(ram[3365]), .B(ram[3381]), .S(n4334), .Z(n1312) );
  MUX2_X1 U10451 ( .A(ram[3333]), .B(ram[3349]), .S(n4334), .Z(n1313) );
  MUX2_X1 U10452 ( .A(n1313), .B(n1312), .S(n4202), .Z(n1314) );
  MUX2_X1 U10453 ( .A(n1314), .B(n1311), .S(n4134), .Z(n1315) );
  MUX2_X1 U10454 ( .A(n1315), .B(n1308), .S(n4094), .Z(n1316) );
  MUX2_X1 U10455 ( .A(ram[3301]), .B(ram[3317]), .S(n4334), .Z(n1317) );
  MUX2_X1 U10456 ( .A(ram[3269]), .B(ram[3285]), .S(n4334), .Z(n1318) );
  MUX2_X1 U10457 ( .A(n1318), .B(n1317), .S(n4202), .Z(n1319) );
  MUX2_X1 U10458 ( .A(ram[3237]), .B(ram[3253]), .S(n4334), .Z(n1320) );
  MUX2_X1 U10459 ( .A(ram[3205]), .B(ram[3221]), .S(n4334), .Z(n1321) );
  MUX2_X1 U10460 ( .A(n1321), .B(n1320), .S(n4202), .Z(n1322) );
  MUX2_X1 U10461 ( .A(n1322), .B(n1319), .S(n4134), .Z(n1323) );
  MUX2_X1 U10462 ( .A(ram[3173]), .B(ram[3189]), .S(n4335), .Z(n1324) );
  MUX2_X1 U10463 ( .A(ram[3141]), .B(ram[3157]), .S(n4335), .Z(n1325) );
  MUX2_X1 U10464 ( .A(n1325), .B(n1324), .S(n4202), .Z(n1326) );
  MUX2_X1 U10465 ( .A(ram[3109]), .B(ram[3125]), .S(n4335), .Z(n1327) );
  MUX2_X1 U10466 ( .A(ram[3077]), .B(ram[3093]), .S(n4335), .Z(n1328) );
  MUX2_X1 U10467 ( .A(n1328), .B(n1327), .S(n4202), .Z(n1329) );
  MUX2_X1 U10468 ( .A(n1329), .B(n1326), .S(n4134), .Z(n1330) );
  MUX2_X1 U10469 ( .A(n1330), .B(n1323), .S(n4094), .Z(n1331) );
  MUX2_X1 U10470 ( .A(n1331), .B(n1316), .S(n4079), .Z(n1332) );
  MUX2_X1 U10471 ( .A(n1332), .B(n1301), .S(n4070), .Z(n1333) );
  MUX2_X1 U10472 ( .A(ram[3045]), .B(ram[3061]), .S(n4335), .Z(n1334) );
  MUX2_X1 U10473 ( .A(ram[3013]), .B(ram[3029]), .S(n4335), .Z(n1335) );
  MUX2_X1 U10474 ( .A(n1335), .B(n1334), .S(n4202), .Z(n1336) );
  MUX2_X1 U10475 ( .A(ram[2981]), .B(ram[2997]), .S(n4335), .Z(n1337) );
  MUX2_X1 U10476 ( .A(ram[2949]), .B(ram[2965]), .S(n4335), .Z(n1338) );
  MUX2_X1 U10477 ( .A(n1338), .B(n1337), .S(n4202), .Z(n1339) );
  MUX2_X1 U10478 ( .A(n1339), .B(n1336), .S(n4134), .Z(n1340) );
  MUX2_X1 U10479 ( .A(ram[2917]), .B(ram[2933]), .S(n4335), .Z(n1341) );
  MUX2_X1 U10480 ( .A(ram[2885]), .B(ram[2901]), .S(n4335), .Z(n1342) );
  MUX2_X1 U10481 ( .A(n1342), .B(n1341), .S(n4202), .Z(n1343) );
  MUX2_X1 U10482 ( .A(ram[2853]), .B(ram[2869]), .S(n4335), .Z(n1344) );
  MUX2_X1 U10483 ( .A(ram[2821]), .B(ram[2837]), .S(n4335), .Z(n1345) );
  MUX2_X1 U10484 ( .A(n1345), .B(n1344), .S(n4202), .Z(n1346) );
  MUX2_X1 U10485 ( .A(n1346), .B(n1343), .S(n4134), .Z(n1347) );
  MUX2_X1 U10486 ( .A(n1347), .B(n1340), .S(n4094), .Z(n1348) );
  MUX2_X1 U10487 ( .A(ram[2789]), .B(ram[2805]), .S(n4336), .Z(n1349) );
  MUX2_X1 U10488 ( .A(ram[2757]), .B(ram[2773]), .S(n4336), .Z(n1350) );
  MUX2_X1 U10489 ( .A(n1350), .B(n1349), .S(n4203), .Z(n1351) );
  MUX2_X1 U10490 ( .A(ram[2725]), .B(ram[2741]), .S(n4336), .Z(n1352) );
  MUX2_X1 U10491 ( .A(ram[2693]), .B(ram[2709]), .S(n4336), .Z(n1353) );
  MUX2_X1 U10492 ( .A(n1353), .B(n1352), .S(n4203), .Z(n1354) );
  MUX2_X1 U10493 ( .A(n1354), .B(n1351), .S(n4134), .Z(n1355) );
  MUX2_X1 U10494 ( .A(ram[2661]), .B(ram[2677]), .S(n4336), .Z(n1356) );
  MUX2_X1 U10495 ( .A(ram[2629]), .B(ram[2645]), .S(n4336), .Z(n1357) );
  MUX2_X1 U10496 ( .A(n1357), .B(n1356), .S(n4203), .Z(n1358) );
  MUX2_X1 U10497 ( .A(ram[2597]), .B(ram[2613]), .S(n4336), .Z(n1359) );
  MUX2_X1 U10498 ( .A(ram[2565]), .B(ram[2581]), .S(n4336), .Z(n1360) );
  MUX2_X1 U10499 ( .A(n1360), .B(n1359), .S(n4203), .Z(n1361) );
  MUX2_X1 U10500 ( .A(n1361), .B(n1358), .S(n4134), .Z(n1362) );
  MUX2_X1 U10501 ( .A(n1362), .B(n1355), .S(n4094), .Z(n1363) );
  MUX2_X1 U10502 ( .A(n1363), .B(n1348), .S(n4079), .Z(n1364) );
  MUX2_X1 U10503 ( .A(ram[2533]), .B(ram[2549]), .S(n4336), .Z(n1365) );
  MUX2_X1 U10504 ( .A(ram[2501]), .B(ram[2517]), .S(n4336), .Z(n1366) );
  MUX2_X1 U10505 ( .A(n1366), .B(n1365), .S(n4203), .Z(n1367) );
  MUX2_X1 U10506 ( .A(ram[2469]), .B(ram[2485]), .S(n4336), .Z(n1368) );
  MUX2_X1 U10507 ( .A(ram[2437]), .B(ram[2453]), .S(n4336), .Z(n1369) );
  MUX2_X1 U10508 ( .A(n1369), .B(n1368), .S(n4203), .Z(n1370) );
  MUX2_X1 U10509 ( .A(n1370), .B(n1367), .S(n4134), .Z(n1371) );
  MUX2_X1 U10510 ( .A(ram[2405]), .B(ram[2421]), .S(n4337), .Z(n1372) );
  MUX2_X1 U10511 ( .A(ram[2373]), .B(ram[2389]), .S(n4337), .Z(n1373) );
  MUX2_X1 U10512 ( .A(n1373), .B(n1372), .S(n4203), .Z(n1374) );
  MUX2_X1 U10513 ( .A(ram[2341]), .B(ram[2357]), .S(n4337), .Z(n1375) );
  MUX2_X1 U10514 ( .A(ram[2309]), .B(ram[2325]), .S(n4337), .Z(n1376) );
  MUX2_X1 U10515 ( .A(n1376), .B(n1375), .S(n4203), .Z(n1377) );
  MUX2_X1 U10516 ( .A(n1377), .B(n1374), .S(n4134), .Z(n1378) );
  MUX2_X1 U10517 ( .A(n1378), .B(n1371), .S(n4094), .Z(n1379) );
  MUX2_X1 U10518 ( .A(ram[2277]), .B(ram[2293]), .S(n4337), .Z(n1380) );
  MUX2_X1 U10519 ( .A(ram[2245]), .B(ram[2261]), .S(n4337), .Z(n1381) );
  MUX2_X1 U10520 ( .A(n1381), .B(n1380), .S(n4203), .Z(n1382) );
  MUX2_X1 U10521 ( .A(ram[2213]), .B(ram[2229]), .S(n4337), .Z(n1383) );
  MUX2_X1 U10522 ( .A(ram[2181]), .B(ram[2197]), .S(n4337), .Z(n1384) );
  MUX2_X1 U10523 ( .A(n1384), .B(n1383), .S(n4203), .Z(n1385) );
  MUX2_X1 U10524 ( .A(n1385), .B(n1382), .S(n4134), .Z(n1386) );
  MUX2_X1 U10525 ( .A(ram[2149]), .B(ram[2165]), .S(n4337), .Z(n1387) );
  MUX2_X1 U10526 ( .A(ram[2117]), .B(ram[2133]), .S(n4337), .Z(n1388) );
  MUX2_X1 U10527 ( .A(n1388), .B(n1387), .S(n4203), .Z(n1389) );
  MUX2_X1 U10528 ( .A(ram[2085]), .B(ram[2101]), .S(n4337), .Z(n1390) );
  MUX2_X1 U10529 ( .A(ram[2053]), .B(ram[2069]), .S(n4337), .Z(n1391) );
  MUX2_X1 U10530 ( .A(n1391), .B(n1390), .S(n4203), .Z(n1392) );
  MUX2_X1 U10531 ( .A(n1392), .B(n1389), .S(n4134), .Z(n1393) );
  MUX2_X1 U10532 ( .A(n1393), .B(n1386), .S(n4094), .Z(n1394) );
  MUX2_X1 U10533 ( .A(n1394), .B(n1379), .S(n4079), .Z(n1395) );
  MUX2_X1 U10534 ( .A(n1395), .B(n1364), .S(n4070), .Z(n1396) );
  MUX2_X1 U10535 ( .A(n1396), .B(n1333), .S(n4066), .Z(n1397) );
  MUX2_X1 U10536 ( .A(ram[2021]), .B(ram[2037]), .S(n4338), .Z(n1398) );
  MUX2_X1 U10537 ( .A(ram[1989]), .B(ram[2005]), .S(n4338), .Z(n1399) );
  MUX2_X1 U10538 ( .A(n1399), .B(n1398), .S(n4204), .Z(n1400) );
  MUX2_X1 U10539 ( .A(ram[1957]), .B(ram[1973]), .S(n4338), .Z(n1401) );
  MUX2_X1 U10540 ( .A(ram[1925]), .B(ram[1941]), .S(n4338), .Z(n1402) );
  MUX2_X1 U10541 ( .A(n1402), .B(n1401), .S(n4204), .Z(n1403) );
  MUX2_X1 U10542 ( .A(n1403), .B(n1400), .S(n4135), .Z(n1404) );
  MUX2_X1 U10543 ( .A(ram[1893]), .B(ram[1909]), .S(n4338), .Z(n1405) );
  MUX2_X1 U10544 ( .A(ram[1861]), .B(ram[1877]), .S(n4338), .Z(n1406) );
  MUX2_X1 U10545 ( .A(n1406), .B(n1405), .S(n4204), .Z(n1407) );
  MUX2_X1 U10546 ( .A(ram[1829]), .B(ram[1845]), .S(n4338), .Z(n1408) );
  MUX2_X1 U10547 ( .A(ram[1797]), .B(ram[1813]), .S(n4338), .Z(n1409) );
  MUX2_X1 U10548 ( .A(n1409), .B(n1408), .S(n4204), .Z(n1410) );
  MUX2_X1 U10549 ( .A(n1410), .B(n1407), .S(n4135), .Z(n1411) );
  MUX2_X1 U10550 ( .A(n1411), .B(n1404), .S(n4095), .Z(n1412) );
  MUX2_X1 U10551 ( .A(ram[1765]), .B(ram[1781]), .S(n4338), .Z(n1413) );
  MUX2_X1 U10552 ( .A(ram[1733]), .B(ram[1749]), .S(n4338), .Z(n1414) );
  MUX2_X1 U10553 ( .A(n1414), .B(n1413), .S(n4204), .Z(n1415) );
  MUX2_X1 U10554 ( .A(ram[1701]), .B(ram[1717]), .S(n4338), .Z(n1416) );
  MUX2_X1 U10555 ( .A(ram[1669]), .B(ram[1685]), .S(n4338), .Z(n1417) );
  MUX2_X1 U10556 ( .A(n1417), .B(n1416), .S(n4204), .Z(n1418) );
  MUX2_X1 U10557 ( .A(n1418), .B(n1415), .S(n4135), .Z(n1419) );
  MUX2_X1 U10558 ( .A(ram[1637]), .B(ram[1653]), .S(n4339), .Z(n1420) );
  MUX2_X1 U10559 ( .A(ram[1605]), .B(ram[1621]), .S(n4339), .Z(n1421) );
  MUX2_X1 U10560 ( .A(n1421), .B(n1420), .S(n4204), .Z(n1422) );
  MUX2_X1 U10561 ( .A(ram[1573]), .B(ram[1589]), .S(n4339), .Z(n1423) );
  MUX2_X1 U10562 ( .A(ram[1541]), .B(ram[1557]), .S(n4339), .Z(n1424) );
  MUX2_X1 U10563 ( .A(n1424), .B(n1423), .S(n4204), .Z(n1425) );
  MUX2_X1 U10564 ( .A(n1425), .B(n1422), .S(n4135), .Z(n1426) );
  MUX2_X1 U10565 ( .A(n1426), .B(n1419), .S(n4095), .Z(n1427) );
  MUX2_X1 U10566 ( .A(n1427), .B(n1412), .S(n4080), .Z(n1428) );
  MUX2_X1 U10567 ( .A(ram[1509]), .B(ram[1525]), .S(n4339), .Z(n1429) );
  MUX2_X1 U10568 ( .A(ram[1477]), .B(ram[1493]), .S(n4339), .Z(n1430) );
  MUX2_X1 U10569 ( .A(n1430), .B(n1429), .S(n4204), .Z(n1431) );
  MUX2_X1 U10570 ( .A(ram[1445]), .B(ram[1461]), .S(n4339), .Z(n1432) );
  MUX2_X1 U10571 ( .A(ram[1413]), .B(ram[1429]), .S(n4339), .Z(n1433) );
  MUX2_X1 U10572 ( .A(n1433), .B(n1432), .S(n4204), .Z(n1434) );
  MUX2_X1 U10573 ( .A(n1434), .B(n1431), .S(n4135), .Z(n1435) );
  MUX2_X1 U10574 ( .A(ram[1381]), .B(ram[1397]), .S(n4339), .Z(n1436) );
  MUX2_X1 U10575 ( .A(ram[1349]), .B(ram[1365]), .S(n4339), .Z(n1437) );
  MUX2_X1 U10576 ( .A(n1437), .B(n1436), .S(n4204), .Z(n1438) );
  MUX2_X1 U10577 ( .A(ram[1317]), .B(ram[1333]), .S(n4339), .Z(n1439) );
  MUX2_X1 U10578 ( .A(ram[1285]), .B(ram[1301]), .S(n4339), .Z(n1440) );
  MUX2_X1 U10579 ( .A(n1440), .B(n1439), .S(n4204), .Z(n1441) );
  MUX2_X1 U10580 ( .A(n1441), .B(n1438), .S(n4135), .Z(n1442) );
  MUX2_X1 U10581 ( .A(n1442), .B(n1435), .S(n4095), .Z(n1443) );
  MUX2_X1 U10582 ( .A(ram[1253]), .B(ram[1269]), .S(n4340), .Z(n1444) );
  MUX2_X1 U10583 ( .A(ram[1221]), .B(ram[1237]), .S(n4340), .Z(n1445) );
  MUX2_X1 U10584 ( .A(n1445), .B(n1444), .S(n4205), .Z(n1446) );
  MUX2_X1 U10585 ( .A(ram[1189]), .B(ram[1205]), .S(n4340), .Z(n1447) );
  MUX2_X1 U10586 ( .A(ram[1157]), .B(ram[1173]), .S(n4340), .Z(n1448) );
  MUX2_X1 U10587 ( .A(n1448), .B(n1447), .S(n4205), .Z(n1449) );
  MUX2_X1 U10588 ( .A(n1449), .B(n1446), .S(n4135), .Z(n1450) );
  MUX2_X1 U10589 ( .A(ram[1125]), .B(ram[1141]), .S(n4340), .Z(n1451) );
  MUX2_X1 U10590 ( .A(ram[1093]), .B(ram[1109]), .S(n4340), .Z(n1452) );
  MUX2_X1 U10591 ( .A(n1452), .B(n1451), .S(n4205), .Z(n1453) );
  MUX2_X1 U10592 ( .A(ram[1061]), .B(ram[1077]), .S(n4340), .Z(n1454) );
  MUX2_X1 U10593 ( .A(ram[1029]), .B(ram[1045]), .S(n4340), .Z(n1455) );
  MUX2_X1 U10594 ( .A(n1455), .B(n1454), .S(n4205), .Z(n1456) );
  MUX2_X1 U10595 ( .A(n1456), .B(n1453), .S(n4135), .Z(n1457) );
  MUX2_X1 U10596 ( .A(n1457), .B(n1450), .S(n4095), .Z(n1458) );
  MUX2_X1 U10597 ( .A(n1458), .B(n1443), .S(n4080), .Z(n1459) );
  MUX2_X1 U10598 ( .A(n1459), .B(n1428), .S(n4070), .Z(n1460) );
  MUX2_X1 U10599 ( .A(ram[997]), .B(ram[1013]), .S(n4340), .Z(n1461) );
  MUX2_X1 U10600 ( .A(ram[965]), .B(ram[981]), .S(n4340), .Z(n1462) );
  MUX2_X1 U10601 ( .A(n1462), .B(n1461), .S(n4205), .Z(n1463) );
  MUX2_X1 U10602 ( .A(ram[933]), .B(ram[949]), .S(n4340), .Z(n1464) );
  MUX2_X1 U10603 ( .A(ram[901]), .B(ram[917]), .S(n4340), .Z(n1465) );
  MUX2_X1 U10604 ( .A(n1465), .B(n1464), .S(n4205), .Z(n1466) );
  MUX2_X1 U10605 ( .A(n1466), .B(n1463), .S(n4135), .Z(n1467) );
  MUX2_X1 U10606 ( .A(ram[869]), .B(ram[885]), .S(n4341), .Z(n1468) );
  MUX2_X1 U10607 ( .A(ram[837]), .B(ram[853]), .S(n4341), .Z(n1469) );
  MUX2_X1 U10608 ( .A(n1469), .B(n1468), .S(n4205), .Z(n1470) );
  MUX2_X1 U10609 ( .A(ram[805]), .B(ram[821]), .S(n4341), .Z(n1471) );
  MUX2_X1 U10610 ( .A(ram[773]), .B(ram[789]), .S(n4341), .Z(n1472) );
  MUX2_X1 U10611 ( .A(n1472), .B(n1471), .S(n4205), .Z(n1473) );
  MUX2_X1 U10612 ( .A(n1473), .B(n1470), .S(n4135), .Z(n1474) );
  MUX2_X1 U10613 ( .A(n1474), .B(n1467), .S(n4095), .Z(n1475) );
  MUX2_X1 U10614 ( .A(ram[741]), .B(ram[757]), .S(n4341), .Z(n1476) );
  MUX2_X1 U10615 ( .A(ram[709]), .B(ram[725]), .S(n4341), .Z(n1477) );
  MUX2_X1 U10616 ( .A(n1477), .B(n1476), .S(n4205), .Z(n1478) );
  MUX2_X1 U10617 ( .A(ram[677]), .B(ram[693]), .S(n4341), .Z(n1479) );
  MUX2_X1 U10618 ( .A(ram[645]), .B(ram[661]), .S(n4341), .Z(n1480) );
  MUX2_X1 U10619 ( .A(n1480), .B(n1479), .S(n4205), .Z(n1481) );
  MUX2_X1 U10620 ( .A(n1481), .B(n1478), .S(n4135), .Z(n1482) );
  MUX2_X1 U10621 ( .A(ram[613]), .B(ram[629]), .S(n4341), .Z(n1483) );
  MUX2_X1 U10622 ( .A(ram[581]), .B(ram[597]), .S(n4341), .Z(n1484) );
  MUX2_X1 U10623 ( .A(n1484), .B(n1483), .S(n4205), .Z(n1485) );
  MUX2_X1 U10624 ( .A(ram[549]), .B(ram[565]), .S(n4341), .Z(n1486) );
  MUX2_X1 U10625 ( .A(ram[517]), .B(ram[533]), .S(n4341), .Z(n1487) );
  MUX2_X1 U10626 ( .A(n1487), .B(n1486), .S(n4205), .Z(n1488) );
  MUX2_X1 U10627 ( .A(n1488), .B(n1485), .S(n4135), .Z(n1489) );
  MUX2_X1 U10628 ( .A(n1489), .B(n1482), .S(n4095), .Z(n1490) );
  MUX2_X1 U10629 ( .A(n1490), .B(n1475), .S(n4080), .Z(n1491) );
  MUX2_X1 U10630 ( .A(ram[485]), .B(ram[501]), .S(n4342), .Z(n1492) );
  MUX2_X1 U10631 ( .A(ram[453]), .B(ram[469]), .S(n4342), .Z(n1493) );
  MUX2_X1 U10632 ( .A(n1493), .B(n1492), .S(n4206), .Z(n1494) );
  MUX2_X1 U10633 ( .A(ram[421]), .B(ram[437]), .S(n4342), .Z(n1495) );
  MUX2_X1 U10634 ( .A(ram[389]), .B(ram[405]), .S(n4342), .Z(n1496) );
  MUX2_X1 U10635 ( .A(n1496), .B(n1495), .S(n4206), .Z(n1497) );
  MUX2_X1 U10636 ( .A(n1497), .B(n1494), .S(n4136), .Z(n1498) );
  MUX2_X1 U10637 ( .A(ram[357]), .B(ram[373]), .S(n4342), .Z(n1499) );
  MUX2_X1 U10638 ( .A(ram[325]), .B(ram[341]), .S(n4342), .Z(n1500) );
  MUX2_X1 U10639 ( .A(n1500), .B(n1499), .S(n4206), .Z(n1501) );
  MUX2_X1 U10640 ( .A(ram[293]), .B(ram[309]), .S(n4342), .Z(n1502) );
  MUX2_X1 U10641 ( .A(ram[261]), .B(ram[277]), .S(n4342), .Z(n1503) );
  MUX2_X1 U10642 ( .A(n1503), .B(n1502), .S(n4206), .Z(n1504) );
  MUX2_X1 U10643 ( .A(n1504), .B(n1501), .S(n4136), .Z(n1505) );
  MUX2_X1 U10644 ( .A(n1505), .B(n1498), .S(n4095), .Z(n1506) );
  MUX2_X1 U10645 ( .A(ram[229]), .B(ram[245]), .S(n4342), .Z(n1507) );
  MUX2_X1 U10646 ( .A(ram[197]), .B(ram[213]), .S(n4342), .Z(n1508) );
  MUX2_X1 U10647 ( .A(n1508), .B(n1507), .S(n4206), .Z(n1509) );
  MUX2_X1 U10648 ( .A(ram[165]), .B(ram[181]), .S(n4342), .Z(n1510) );
  MUX2_X1 U10649 ( .A(ram[133]), .B(ram[149]), .S(n4342), .Z(n1511) );
  MUX2_X1 U10650 ( .A(n1511), .B(n1510), .S(n4206), .Z(n1512) );
  MUX2_X1 U10651 ( .A(n1512), .B(n1509), .S(n4136), .Z(n1513) );
  MUX2_X1 U10652 ( .A(ram[101]), .B(ram[117]), .S(n4343), .Z(n1514) );
  MUX2_X1 U10653 ( .A(ram[69]), .B(ram[85]), .S(n4343), .Z(n1515) );
  MUX2_X1 U10654 ( .A(n1515), .B(n1514), .S(n4206), .Z(n1516) );
  MUX2_X1 U10655 ( .A(ram[37]), .B(ram[53]), .S(n4343), .Z(n1517) );
  MUX2_X1 U10656 ( .A(ram[5]), .B(ram[21]), .S(n4343), .Z(n1518) );
  MUX2_X1 U10657 ( .A(n1518), .B(n1517), .S(n4206), .Z(n1519) );
  MUX2_X1 U10658 ( .A(n1519), .B(n1516), .S(n4136), .Z(n1520) );
  MUX2_X1 U10659 ( .A(n1520), .B(n1513), .S(n4095), .Z(n1521) );
  MUX2_X1 U10660 ( .A(n1521), .B(n1506), .S(n4080), .Z(n1522) );
  MUX2_X1 U10661 ( .A(n1522), .B(n1491), .S(n4070), .Z(n1523) );
  MUX2_X1 U10662 ( .A(n1523), .B(n1460), .S(n4066), .Z(n1524) );
  MUX2_X1 U10663 ( .A(n1524), .B(n1397), .S(mem_access_addr[9]), .Z(N296) );
  MUX2_X1 U10664 ( .A(ram[4070]), .B(ram[4086]), .S(n4343), .Z(n1525) );
  MUX2_X1 U10665 ( .A(ram[4038]), .B(ram[4054]), .S(n4343), .Z(n1526) );
  MUX2_X1 U10666 ( .A(n1526), .B(n1525), .S(n4206), .Z(n1527) );
  MUX2_X1 U10667 ( .A(ram[4006]), .B(ram[4022]), .S(n4343), .Z(n1528) );
  MUX2_X1 U10668 ( .A(ram[3974]), .B(ram[3990]), .S(n4343), .Z(n1529) );
  MUX2_X1 U10669 ( .A(n1529), .B(n1528), .S(n4206), .Z(n1530) );
  MUX2_X1 U10670 ( .A(n1530), .B(n1527), .S(n4136), .Z(n1531) );
  MUX2_X1 U10671 ( .A(ram[3942]), .B(ram[3958]), .S(n4343), .Z(n1532) );
  MUX2_X1 U10672 ( .A(ram[3910]), .B(ram[3926]), .S(n4343), .Z(n1533) );
  MUX2_X1 U10673 ( .A(n1533), .B(n1532), .S(n4206), .Z(n1534) );
  MUX2_X1 U10674 ( .A(ram[3878]), .B(ram[3894]), .S(n4343), .Z(n1535) );
  MUX2_X1 U10675 ( .A(ram[3846]), .B(ram[3862]), .S(n4343), .Z(n1536) );
  MUX2_X1 U10676 ( .A(n1536), .B(n1535), .S(n4206), .Z(n1537) );
  MUX2_X1 U10677 ( .A(n1537), .B(n1534), .S(n4136), .Z(n1538) );
  MUX2_X1 U10678 ( .A(n1538), .B(n1531), .S(n4095), .Z(n1539) );
  MUX2_X1 U10679 ( .A(ram[3814]), .B(ram[3830]), .S(n4344), .Z(n1540) );
  MUX2_X1 U10680 ( .A(ram[3782]), .B(ram[3798]), .S(n4344), .Z(n1541) );
  MUX2_X1 U10681 ( .A(n1541), .B(n1540), .S(n4207), .Z(n1542) );
  MUX2_X1 U10682 ( .A(ram[3750]), .B(ram[3766]), .S(n4344), .Z(n1543) );
  MUX2_X1 U10683 ( .A(ram[3718]), .B(ram[3734]), .S(n4344), .Z(n1544) );
  MUX2_X1 U10684 ( .A(n1544), .B(n1543), .S(n4207), .Z(n1545) );
  MUX2_X1 U10685 ( .A(n1545), .B(n1542), .S(n4136), .Z(n1546) );
  MUX2_X1 U10686 ( .A(ram[3686]), .B(ram[3702]), .S(n4344), .Z(n1547) );
  MUX2_X1 U10687 ( .A(ram[3654]), .B(ram[3670]), .S(n4344), .Z(n1548) );
  MUX2_X1 U10688 ( .A(n1548), .B(n1547), .S(n4207), .Z(n1549) );
  MUX2_X1 U10689 ( .A(ram[3622]), .B(ram[3638]), .S(n4344), .Z(n1550) );
  MUX2_X1 U10690 ( .A(ram[3590]), .B(ram[3606]), .S(n4344), .Z(n1551) );
  MUX2_X1 U10691 ( .A(n1551), .B(n1550), .S(n4207), .Z(n1552) );
  MUX2_X1 U10692 ( .A(n1552), .B(n1549), .S(n4136), .Z(n1553) );
  MUX2_X1 U10693 ( .A(n1553), .B(n1546), .S(n4095), .Z(n1554) );
  MUX2_X1 U10694 ( .A(n1554), .B(n1539), .S(n4080), .Z(n1555) );
  MUX2_X1 U10695 ( .A(ram[3558]), .B(ram[3574]), .S(n4344), .Z(n1556) );
  MUX2_X1 U10696 ( .A(ram[3526]), .B(ram[3542]), .S(n4344), .Z(n1557) );
  MUX2_X1 U10697 ( .A(n1557), .B(n1556), .S(n4207), .Z(n1558) );
  MUX2_X1 U10698 ( .A(ram[3494]), .B(ram[3510]), .S(n4344), .Z(n1559) );
  MUX2_X1 U10699 ( .A(ram[3462]), .B(ram[3478]), .S(n4344), .Z(n1560) );
  MUX2_X1 U10700 ( .A(n1560), .B(n1559), .S(n4207), .Z(n1561) );
  MUX2_X1 U10701 ( .A(n1561), .B(n1558), .S(n4136), .Z(n1562) );
  MUX2_X1 U10702 ( .A(ram[3430]), .B(ram[3446]), .S(n4345), .Z(n1563) );
  MUX2_X1 U10703 ( .A(ram[3398]), .B(ram[3414]), .S(n4345), .Z(n1564) );
  MUX2_X1 U10704 ( .A(n1564), .B(n1563), .S(n4207), .Z(n1565) );
  MUX2_X1 U10705 ( .A(ram[3366]), .B(ram[3382]), .S(n4345), .Z(n1566) );
  MUX2_X1 U10706 ( .A(ram[3334]), .B(ram[3350]), .S(n4345), .Z(n1567) );
  MUX2_X1 U10707 ( .A(n1567), .B(n1566), .S(n4207), .Z(n1568) );
  MUX2_X1 U10708 ( .A(n1568), .B(n1565), .S(n4136), .Z(n1569) );
  MUX2_X1 U10709 ( .A(n1569), .B(n1562), .S(n4095), .Z(n1570) );
  MUX2_X1 U10710 ( .A(ram[3302]), .B(ram[3318]), .S(n4345), .Z(n1571) );
  MUX2_X1 U10711 ( .A(ram[3270]), .B(ram[3286]), .S(n4345), .Z(n1572) );
  MUX2_X1 U10712 ( .A(n1572), .B(n1571), .S(n4207), .Z(n1573) );
  MUX2_X1 U10713 ( .A(ram[3238]), .B(ram[3254]), .S(n4345), .Z(n1574) );
  MUX2_X1 U10714 ( .A(ram[3206]), .B(ram[3222]), .S(n4345), .Z(n1575) );
  MUX2_X1 U10715 ( .A(n1575), .B(n1574), .S(n4207), .Z(n1576) );
  MUX2_X1 U10716 ( .A(n1576), .B(n1573), .S(n4136), .Z(n1577) );
  MUX2_X1 U10717 ( .A(ram[3174]), .B(ram[3190]), .S(n4345), .Z(n1578) );
  MUX2_X1 U10718 ( .A(ram[3142]), .B(ram[3158]), .S(n4345), .Z(n1579) );
  MUX2_X1 U10719 ( .A(n1579), .B(n1578), .S(n4207), .Z(n1580) );
  MUX2_X1 U10720 ( .A(ram[3110]), .B(ram[3126]), .S(n4345), .Z(n1581) );
  MUX2_X1 U10721 ( .A(ram[3078]), .B(ram[3094]), .S(n4345), .Z(n1582) );
  MUX2_X1 U10722 ( .A(n1582), .B(n1581), .S(n4207), .Z(n1583) );
  MUX2_X1 U10723 ( .A(n1583), .B(n1580), .S(n4136), .Z(n1584) );
  MUX2_X1 U10724 ( .A(n1584), .B(n1577), .S(n4095), .Z(n1585) );
  MUX2_X1 U10725 ( .A(n1585), .B(n1570), .S(n4080), .Z(n1586) );
  MUX2_X1 U10726 ( .A(n1586), .B(n1555), .S(n4070), .Z(n1587) );
  MUX2_X1 U10727 ( .A(ram[3046]), .B(ram[3062]), .S(n4346), .Z(n1588) );
  MUX2_X1 U10728 ( .A(ram[3014]), .B(ram[3030]), .S(n4346), .Z(n1589) );
  MUX2_X1 U10729 ( .A(n1589), .B(n1588), .S(n4208), .Z(n1590) );
  MUX2_X1 U10730 ( .A(ram[2982]), .B(ram[2998]), .S(n4346), .Z(n1591) );
  MUX2_X1 U10731 ( .A(ram[2950]), .B(ram[2966]), .S(n4346), .Z(n1592) );
  MUX2_X1 U10732 ( .A(n1592), .B(n1591), .S(n4208), .Z(n1593) );
  MUX2_X1 U10733 ( .A(n1593), .B(n1590), .S(n4137), .Z(n1594) );
  MUX2_X1 U10734 ( .A(ram[2918]), .B(ram[2934]), .S(n4346), .Z(n1595) );
  MUX2_X1 U10735 ( .A(ram[2886]), .B(ram[2902]), .S(n4346), .Z(n1596) );
  MUX2_X1 U10736 ( .A(n1596), .B(n1595), .S(n4208), .Z(n1597) );
  MUX2_X1 U10737 ( .A(ram[2854]), .B(ram[2870]), .S(n4346), .Z(n1598) );
  MUX2_X1 U10738 ( .A(ram[2822]), .B(ram[2838]), .S(n4346), .Z(n1599) );
  MUX2_X1 U10739 ( .A(n1599), .B(n1598), .S(n4208), .Z(n1600) );
  MUX2_X1 U10740 ( .A(n1600), .B(n1597), .S(n4137), .Z(n1601) );
  MUX2_X1 U10741 ( .A(n1601), .B(n1594), .S(n4096), .Z(n1602) );
  MUX2_X1 U10742 ( .A(ram[2790]), .B(ram[2806]), .S(n4346), .Z(n1603) );
  MUX2_X1 U10743 ( .A(ram[2758]), .B(ram[2774]), .S(n4346), .Z(n1604) );
  MUX2_X1 U10744 ( .A(n1604), .B(n1603), .S(n4208), .Z(n1605) );
  MUX2_X1 U10745 ( .A(ram[2726]), .B(ram[2742]), .S(n4346), .Z(n1606) );
  MUX2_X1 U10746 ( .A(ram[2694]), .B(ram[2710]), .S(n4346), .Z(n1607) );
  MUX2_X1 U10747 ( .A(n1607), .B(n1606), .S(n4208), .Z(n1608) );
  MUX2_X1 U10748 ( .A(n1608), .B(n1605), .S(n4137), .Z(n1609) );
  MUX2_X1 U10749 ( .A(ram[2662]), .B(ram[2678]), .S(n4347), .Z(n1610) );
  MUX2_X1 U10750 ( .A(ram[2630]), .B(ram[2646]), .S(n4347), .Z(n1611) );
  MUX2_X1 U10751 ( .A(n1611), .B(n1610), .S(n4208), .Z(n1612) );
  MUX2_X1 U10752 ( .A(ram[2598]), .B(ram[2614]), .S(n4347), .Z(n1613) );
  MUX2_X1 U10753 ( .A(ram[2566]), .B(ram[2582]), .S(n4347), .Z(n1614) );
  MUX2_X1 U10754 ( .A(n1614), .B(n1613), .S(n4208), .Z(n1615) );
  MUX2_X1 U10755 ( .A(n1615), .B(n1612), .S(n4137), .Z(n1616) );
  MUX2_X1 U10756 ( .A(n1616), .B(n1609), .S(n4096), .Z(n1617) );
  MUX2_X1 U10757 ( .A(n1617), .B(n1602), .S(n4080), .Z(n1618) );
  MUX2_X1 U10758 ( .A(ram[2534]), .B(ram[2550]), .S(n4347), .Z(n1619) );
  MUX2_X1 U10759 ( .A(ram[2502]), .B(ram[2518]), .S(n4347), .Z(n1620) );
  MUX2_X1 U10760 ( .A(n1620), .B(n1619), .S(n4208), .Z(n1621) );
  MUX2_X1 U10761 ( .A(ram[2470]), .B(ram[2486]), .S(n4347), .Z(n1622) );
  MUX2_X1 U10762 ( .A(ram[2438]), .B(ram[2454]), .S(n4347), .Z(n1623) );
  MUX2_X1 U10763 ( .A(n1623), .B(n1622), .S(n4208), .Z(n1624) );
  MUX2_X1 U10764 ( .A(n1624), .B(n1621), .S(n4137), .Z(n1625) );
  MUX2_X1 U10765 ( .A(ram[2406]), .B(ram[2422]), .S(n4347), .Z(n1626) );
  MUX2_X1 U10766 ( .A(ram[2374]), .B(ram[2390]), .S(n4347), .Z(n1627) );
  MUX2_X1 U10767 ( .A(n1627), .B(n1626), .S(n4208), .Z(n1628) );
  MUX2_X1 U10768 ( .A(ram[2342]), .B(ram[2358]), .S(n4347), .Z(n1629) );
  MUX2_X1 U10769 ( .A(ram[2310]), .B(ram[2326]), .S(n4347), .Z(n1630) );
  MUX2_X1 U10770 ( .A(n1630), .B(n1629), .S(n4208), .Z(n1631) );
  MUX2_X1 U10771 ( .A(n1631), .B(n1628), .S(n4137), .Z(n1632) );
  MUX2_X1 U10772 ( .A(n1632), .B(n1625), .S(n4096), .Z(n1633) );
  MUX2_X1 U10773 ( .A(ram[2278]), .B(ram[2294]), .S(n4348), .Z(n1634) );
  MUX2_X1 U10774 ( .A(ram[2246]), .B(ram[2262]), .S(n4348), .Z(n1635) );
  MUX2_X1 U10775 ( .A(n1635), .B(n1634), .S(n4209), .Z(n1636) );
  MUX2_X1 U10776 ( .A(ram[2214]), .B(ram[2230]), .S(n4348), .Z(n1637) );
  MUX2_X1 U10777 ( .A(ram[2182]), .B(ram[2198]), .S(n4348), .Z(n1638) );
  MUX2_X1 U10778 ( .A(n1638), .B(n1637), .S(n4209), .Z(n1639) );
  MUX2_X1 U10779 ( .A(n1639), .B(n1636), .S(n4137), .Z(n1640) );
  MUX2_X1 U10780 ( .A(ram[2150]), .B(ram[2166]), .S(n4348), .Z(n1641) );
  MUX2_X1 U10781 ( .A(ram[2118]), .B(ram[2134]), .S(n4348), .Z(n1642) );
  MUX2_X1 U10782 ( .A(n1642), .B(n1641), .S(n4209), .Z(n1643) );
  MUX2_X1 U10783 ( .A(ram[2086]), .B(ram[2102]), .S(n4348), .Z(n1644) );
  MUX2_X1 U10784 ( .A(ram[2054]), .B(ram[2070]), .S(n4348), .Z(n1645) );
  MUX2_X1 U10785 ( .A(n1645), .B(n1644), .S(n4209), .Z(n1646) );
  MUX2_X1 U10786 ( .A(n1646), .B(n1643), .S(n4137), .Z(n1647) );
  MUX2_X1 U10787 ( .A(n1647), .B(n1640), .S(n4096), .Z(n1648) );
  MUX2_X1 U10788 ( .A(n1648), .B(n1633), .S(n4080), .Z(n1649) );
  MUX2_X1 U10789 ( .A(n1649), .B(n1618), .S(n4070), .Z(n1650) );
  MUX2_X1 U10790 ( .A(n1650), .B(n1587), .S(n4066), .Z(n1651) );
  MUX2_X1 U10791 ( .A(ram[2022]), .B(ram[2038]), .S(n4348), .Z(n1652) );
  MUX2_X1 U10792 ( .A(ram[1990]), .B(ram[2006]), .S(n4348), .Z(n1653) );
  MUX2_X1 U10793 ( .A(n1653), .B(n1652), .S(n4209), .Z(n1654) );
  MUX2_X1 U10794 ( .A(ram[1958]), .B(ram[1974]), .S(n4348), .Z(n1655) );
  MUX2_X1 U10795 ( .A(ram[1926]), .B(ram[1942]), .S(n4348), .Z(n1656) );
  MUX2_X1 U10796 ( .A(n1656), .B(n1655), .S(n4209), .Z(n1657) );
  MUX2_X1 U10797 ( .A(n1657), .B(n1654), .S(n4137), .Z(n1658) );
  MUX2_X1 U10798 ( .A(ram[1894]), .B(ram[1910]), .S(n4349), .Z(n1659) );
  MUX2_X1 U10799 ( .A(ram[1862]), .B(ram[1878]), .S(n4349), .Z(n1660) );
  MUX2_X1 U10800 ( .A(n1660), .B(n1659), .S(n4209), .Z(n1661) );
  MUX2_X1 U10801 ( .A(ram[1830]), .B(ram[1846]), .S(n4349), .Z(n1662) );
  MUX2_X1 U10802 ( .A(ram[1798]), .B(ram[1814]), .S(n4349), .Z(n1663) );
  MUX2_X1 U10803 ( .A(n1663), .B(n1662), .S(n4209), .Z(n1664) );
  MUX2_X1 U10804 ( .A(n1664), .B(n1661), .S(n4137), .Z(n1665) );
  MUX2_X1 U10805 ( .A(n1665), .B(n1658), .S(n4096), .Z(n1666) );
  MUX2_X1 U10806 ( .A(ram[1766]), .B(ram[1782]), .S(n4349), .Z(n1667) );
  MUX2_X1 U10807 ( .A(ram[1734]), .B(ram[1750]), .S(n4349), .Z(n1668) );
  MUX2_X1 U10808 ( .A(n1668), .B(n1667), .S(n4209), .Z(n1669) );
  MUX2_X1 U10809 ( .A(ram[1702]), .B(ram[1718]), .S(n4349), .Z(n1670) );
  MUX2_X1 U10810 ( .A(ram[1670]), .B(ram[1686]), .S(n4349), .Z(n1671) );
  MUX2_X1 U10811 ( .A(n1671), .B(n1670), .S(n4209), .Z(n1672) );
  MUX2_X1 U10812 ( .A(n1672), .B(n1669), .S(n4137), .Z(n1673) );
  MUX2_X1 U10813 ( .A(ram[1638]), .B(ram[1654]), .S(n4349), .Z(n1674) );
  MUX2_X1 U10814 ( .A(ram[1606]), .B(ram[1622]), .S(n4349), .Z(n1675) );
  MUX2_X1 U10815 ( .A(n1675), .B(n1674), .S(n4209), .Z(n1676) );
  MUX2_X1 U10816 ( .A(ram[1574]), .B(ram[1590]), .S(n4349), .Z(n1677) );
  MUX2_X1 U10817 ( .A(ram[1542]), .B(ram[1558]), .S(n4349), .Z(n1678) );
  MUX2_X1 U10818 ( .A(n1678), .B(n1677), .S(n4209), .Z(n1679) );
  MUX2_X1 U10819 ( .A(n1679), .B(n1676), .S(n4137), .Z(n1680) );
  MUX2_X1 U10820 ( .A(n1680), .B(n1673), .S(n4096), .Z(n1681) );
  MUX2_X1 U10821 ( .A(n1681), .B(n1666), .S(n4080), .Z(n1682) );
  MUX2_X1 U10822 ( .A(ram[1510]), .B(ram[1526]), .S(n4350), .Z(n1683) );
  MUX2_X1 U10823 ( .A(ram[1478]), .B(ram[1494]), .S(n4350), .Z(n1684) );
  MUX2_X1 U10824 ( .A(n1684), .B(n1683), .S(n4210), .Z(n1685) );
  MUX2_X1 U10825 ( .A(ram[1446]), .B(ram[1462]), .S(n4350), .Z(n1686) );
  MUX2_X1 U10826 ( .A(ram[1414]), .B(ram[1430]), .S(n4350), .Z(n1687) );
  MUX2_X1 U10827 ( .A(n1687), .B(n1686), .S(n4210), .Z(n1688) );
  MUX2_X1 U10828 ( .A(n1688), .B(n1685), .S(n4138), .Z(n1689) );
  MUX2_X1 U10829 ( .A(ram[1382]), .B(ram[1398]), .S(n4350), .Z(n1690) );
  MUX2_X1 U10830 ( .A(ram[1350]), .B(ram[1366]), .S(n4350), .Z(n1691) );
  MUX2_X1 U10831 ( .A(n1691), .B(n1690), .S(n4210), .Z(n1692) );
  MUX2_X1 U10832 ( .A(ram[1318]), .B(ram[1334]), .S(n4350), .Z(n1693) );
  MUX2_X1 U10833 ( .A(ram[1286]), .B(ram[1302]), .S(n4350), .Z(n1694) );
  MUX2_X1 U10834 ( .A(n1694), .B(n1693), .S(n4210), .Z(n1695) );
  MUX2_X1 U10835 ( .A(n1695), .B(n1692), .S(n4138), .Z(n1696) );
  MUX2_X1 U10836 ( .A(n1696), .B(n1689), .S(n4096), .Z(n1697) );
  MUX2_X1 U10837 ( .A(ram[1254]), .B(ram[1270]), .S(n4350), .Z(n1698) );
  MUX2_X1 U10838 ( .A(ram[1222]), .B(ram[1238]), .S(n4350), .Z(n1699) );
  MUX2_X1 U10839 ( .A(n1699), .B(n1698), .S(n4210), .Z(n1700) );
  MUX2_X1 U10840 ( .A(ram[1190]), .B(ram[1206]), .S(n4350), .Z(n1701) );
  MUX2_X1 U10841 ( .A(ram[1158]), .B(ram[1174]), .S(n4350), .Z(n1702) );
  MUX2_X1 U10842 ( .A(n1702), .B(n1701), .S(n4210), .Z(n1703) );
  MUX2_X1 U10843 ( .A(n1703), .B(n1700), .S(n4138), .Z(n1704) );
  MUX2_X1 U10844 ( .A(ram[1126]), .B(ram[1142]), .S(n4351), .Z(n1705) );
  MUX2_X1 U10845 ( .A(ram[1094]), .B(ram[1110]), .S(n4351), .Z(n1706) );
  MUX2_X1 U10846 ( .A(n1706), .B(n1705), .S(n4210), .Z(n1707) );
  MUX2_X1 U10847 ( .A(ram[1062]), .B(ram[1078]), .S(n4351), .Z(n1708) );
  MUX2_X1 U10848 ( .A(ram[1030]), .B(ram[1046]), .S(n4351), .Z(n1709) );
  MUX2_X1 U10849 ( .A(n1709), .B(n1708), .S(n4210), .Z(n1710) );
  MUX2_X1 U10850 ( .A(n1710), .B(n1707), .S(n4138), .Z(n1711) );
  MUX2_X1 U10851 ( .A(n1711), .B(n1704), .S(n4096), .Z(n1712) );
  MUX2_X1 U10852 ( .A(n1712), .B(n1697), .S(n4080), .Z(n1713) );
  MUX2_X1 U10853 ( .A(n1713), .B(n1682), .S(n4070), .Z(n1714) );
  MUX2_X1 U10854 ( .A(ram[998]), .B(ram[1014]), .S(n4351), .Z(n1715) );
  MUX2_X1 U10855 ( .A(ram[966]), .B(ram[982]), .S(n4351), .Z(n1716) );
  MUX2_X1 U10856 ( .A(n1716), .B(n1715), .S(n4210), .Z(n1717) );
  MUX2_X1 U10857 ( .A(ram[934]), .B(ram[950]), .S(n4351), .Z(n1718) );
  MUX2_X1 U10858 ( .A(ram[902]), .B(ram[918]), .S(n4351), .Z(n1719) );
  MUX2_X1 U10859 ( .A(n1719), .B(n1718), .S(n4210), .Z(n1720) );
  MUX2_X1 U10860 ( .A(n1720), .B(n1717), .S(n4138), .Z(n1721) );
  MUX2_X1 U10861 ( .A(ram[870]), .B(ram[886]), .S(n4351), .Z(n1722) );
  MUX2_X1 U10862 ( .A(ram[838]), .B(ram[854]), .S(n4351), .Z(n1723) );
  MUX2_X1 U10863 ( .A(n1723), .B(n1722), .S(n4210), .Z(n1724) );
  MUX2_X1 U10864 ( .A(ram[806]), .B(ram[822]), .S(n4351), .Z(n1725) );
  MUX2_X1 U10865 ( .A(ram[774]), .B(ram[790]), .S(n4351), .Z(n1726) );
  MUX2_X1 U10866 ( .A(n1726), .B(n1725), .S(n4210), .Z(n1727) );
  MUX2_X1 U10867 ( .A(n1727), .B(n1724), .S(n4138), .Z(n1728) );
  MUX2_X1 U10868 ( .A(n1728), .B(n1721), .S(n4096), .Z(n1729) );
  MUX2_X1 U10869 ( .A(ram[742]), .B(ram[758]), .S(n4352), .Z(n1730) );
  MUX2_X1 U10870 ( .A(ram[710]), .B(ram[726]), .S(n4352), .Z(n1731) );
  MUX2_X1 U10871 ( .A(n1731), .B(n1730), .S(n4211), .Z(n1732) );
  MUX2_X1 U10872 ( .A(ram[678]), .B(ram[694]), .S(n4352), .Z(n1733) );
  MUX2_X1 U10873 ( .A(ram[646]), .B(ram[662]), .S(n4352), .Z(n1734) );
  MUX2_X1 U10874 ( .A(n1734), .B(n1733), .S(n4211), .Z(n1735) );
  MUX2_X1 U10875 ( .A(n1735), .B(n1732), .S(n4138), .Z(n1736) );
  MUX2_X1 U10876 ( .A(ram[614]), .B(ram[630]), .S(n4352), .Z(n1737) );
  MUX2_X1 U10877 ( .A(ram[582]), .B(ram[598]), .S(n4352), .Z(n1738) );
  MUX2_X1 U10878 ( .A(n1738), .B(n1737), .S(n4211), .Z(n1739) );
  MUX2_X1 U10879 ( .A(ram[550]), .B(ram[566]), .S(n4352), .Z(n1740) );
  MUX2_X1 U10880 ( .A(ram[518]), .B(ram[534]), .S(n4352), .Z(n1741) );
  MUX2_X1 U10881 ( .A(n1741), .B(n1740), .S(n4211), .Z(n1742) );
  MUX2_X1 U10882 ( .A(n1742), .B(n1739), .S(n4138), .Z(n1743) );
  MUX2_X1 U10883 ( .A(n1743), .B(n1736), .S(n4096), .Z(n1744) );
  MUX2_X1 U10884 ( .A(n1744), .B(n1729), .S(n4080), .Z(n1745) );
  MUX2_X1 U10885 ( .A(ram[486]), .B(ram[502]), .S(n4352), .Z(n1746) );
  MUX2_X1 U10886 ( .A(ram[454]), .B(ram[470]), .S(n4352), .Z(n1747) );
  MUX2_X1 U10887 ( .A(n1747), .B(n1746), .S(n4211), .Z(n1748) );
  MUX2_X1 U10888 ( .A(ram[422]), .B(ram[438]), .S(n4352), .Z(n1749) );
  MUX2_X1 U10889 ( .A(ram[390]), .B(ram[406]), .S(n4352), .Z(n1750) );
  MUX2_X1 U10890 ( .A(n1750), .B(n1749), .S(n4211), .Z(n1751) );
  MUX2_X1 U10891 ( .A(n1751), .B(n1748), .S(n4138), .Z(n1752) );
  MUX2_X1 U10892 ( .A(ram[358]), .B(ram[374]), .S(n4353), .Z(n1753) );
  MUX2_X1 U10893 ( .A(ram[326]), .B(ram[342]), .S(n4353), .Z(n1754) );
  MUX2_X1 U10894 ( .A(n1754), .B(n1753), .S(n4211), .Z(n1755) );
  MUX2_X1 U10895 ( .A(ram[294]), .B(ram[310]), .S(n4353), .Z(n1756) );
  MUX2_X1 U10896 ( .A(ram[262]), .B(ram[278]), .S(n4353), .Z(n1757) );
  MUX2_X1 U10897 ( .A(n1757), .B(n1756), .S(n4211), .Z(n1758) );
  MUX2_X1 U10898 ( .A(n1758), .B(n1755), .S(n4138), .Z(n1759) );
  MUX2_X1 U10899 ( .A(n1759), .B(n1752), .S(n4096), .Z(n1760) );
  MUX2_X1 U10900 ( .A(ram[230]), .B(ram[246]), .S(n4353), .Z(n1761) );
  MUX2_X1 U10901 ( .A(ram[198]), .B(ram[214]), .S(n4353), .Z(n1762) );
  MUX2_X1 U10902 ( .A(n1762), .B(n1761), .S(n4211), .Z(n1763) );
  MUX2_X1 U10903 ( .A(ram[166]), .B(ram[182]), .S(n4353), .Z(n1764) );
  MUX2_X1 U10904 ( .A(ram[134]), .B(ram[150]), .S(n4353), .Z(n1765) );
  MUX2_X1 U10905 ( .A(n1765), .B(n1764), .S(n4211), .Z(n1766) );
  MUX2_X1 U10906 ( .A(n1766), .B(n1763), .S(n4138), .Z(n1767) );
  MUX2_X1 U10907 ( .A(ram[102]), .B(ram[118]), .S(n4353), .Z(n1768) );
  MUX2_X1 U10908 ( .A(ram[70]), .B(ram[86]), .S(n4353), .Z(n1769) );
  MUX2_X1 U10909 ( .A(n1769), .B(n1768), .S(n4211), .Z(n1770) );
  MUX2_X1 U10910 ( .A(ram[38]), .B(ram[54]), .S(n4353), .Z(n1771) );
  MUX2_X1 U10911 ( .A(ram[6]), .B(ram[22]), .S(n4353), .Z(n1772) );
  MUX2_X1 U10912 ( .A(n1772), .B(n1771), .S(n4211), .Z(n1773) );
  MUX2_X1 U10913 ( .A(n1773), .B(n1770), .S(n4138), .Z(n1774) );
  MUX2_X1 U10914 ( .A(n1774), .B(n1767), .S(n4096), .Z(n1775) );
  MUX2_X1 U10915 ( .A(n1775), .B(n1760), .S(n4080), .Z(n1776) );
  MUX2_X1 U10916 ( .A(n1776), .B(n1745), .S(n4070), .Z(n1777) );
  MUX2_X1 U10917 ( .A(n1777), .B(n1714), .S(n4066), .Z(n1778) );
  MUX2_X1 U10918 ( .A(n1778), .B(n1651), .S(mem_access_addr[9]), .Z(N295) );
  MUX2_X1 U10919 ( .A(ram[4071]), .B(ram[4087]), .S(n4354), .Z(n1779) );
  MUX2_X1 U10920 ( .A(ram[4039]), .B(ram[4055]), .S(n4354), .Z(n1780) );
  MUX2_X1 U10921 ( .A(n1780), .B(n1779), .S(n4212), .Z(n1781) );
  MUX2_X1 U10922 ( .A(ram[4007]), .B(ram[4023]), .S(n4354), .Z(n1782) );
  MUX2_X1 U10923 ( .A(ram[3975]), .B(ram[3991]), .S(n4354), .Z(n1783) );
  MUX2_X1 U10924 ( .A(n1783), .B(n1782), .S(n4212), .Z(n1784) );
  MUX2_X1 U10925 ( .A(n1784), .B(n1781), .S(n4139), .Z(n1785) );
  MUX2_X1 U10926 ( .A(ram[3943]), .B(ram[3959]), .S(n4354), .Z(n1786) );
  MUX2_X1 U10927 ( .A(ram[3911]), .B(ram[3927]), .S(n4354), .Z(n1787) );
  MUX2_X1 U10928 ( .A(n1787), .B(n1786), .S(n4212), .Z(n1788) );
  MUX2_X1 U10929 ( .A(ram[3879]), .B(ram[3895]), .S(n4354), .Z(n1789) );
  MUX2_X1 U10930 ( .A(ram[3847]), .B(ram[3863]), .S(n4354), .Z(n1790) );
  MUX2_X1 U10931 ( .A(n1790), .B(n1789), .S(n4212), .Z(n1791) );
  MUX2_X1 U10932 ( .A(n1791), .B(n1788), .S(n4139), .Z(n1792) );
  MUX2_X1 U10933 ( .A(n1792), .B(n1785), .S(n4097), .Z(n1793) );
  MUX2_X1 U10934 ( .A(ram[3815]), .B(ram[3831]), .S(n4354), .Z(n1794) );
  MUX2_X1 U10935 ( .A(ram[3783]), .B(ram[3799]), .S(n4354), .Z(n1795) );
  MUX2_X1 U10936 ( .A(n1795), .B(n1794), .S(n4212), .Z(n1796) );
  MUX2_X1 U10937 ( .A(ram[3751]), .B(ram[3767]), .S(n4354), .Z(n1797) );
  MUX2_X1 U10938 ( .A(ram[3719]), .B(ram[3735]), .S(n4354), .Z(n1798) );
  MUX2_X1 U10939 ( .A(n1798), .B(n1797), .S(n4212), .Z(n1799) );
  MUX2_X1 U10940 ( .A(n1799), .B(n1796), .S(n4139), .Z(n1800) );
  MUX2_X1 U10941 ( .A(ram[3687]), .B(ram[3703]), .S(n4355), .Z(n1801) );
  MUX2_X1 U10942 ( .A(ram[3655]), .B(ram[3671]), .S(n4355), .Z(n1802) );
  MUX2_X1 U10943 ( .A(n1802), .B(n1801), .S(n4212), .Z(n1803) );
  MUX2_X1 U10944 ( .A(ram[3623]), .B(ram[3639]), .S(n4355), .Z(n1804) );
  MUX2_X1 U10945 ( .A(ram[3591]), .B(ram[3607]), .S(n4355), .Z(n1805) );
  MUX2_X1 U10946 ( .A(n1805), .B(n1804), .S(n4212), .Z(n1806) );
  MUX2_X1 U10947 ( .A(n1806), .B(n1803), .S(n4139), .Z(n1807) );
  MUX2_X1 U10948 ( .A(n1807), .B(n1800), .S(n4097), .Z(n1808) );
  MUX2_X1 U10949 ( .A(n1808), .B(n1793), .S(n4081), .Z(n1809) );
  MUX2_X1 U10950 ( .A(ram[3559]), .B(ram[3575]), .S(n4355), .Z(n1810) );
  MUX2_X1 U10951 ( .A(ram[3527]), .B(ram[3543]), .S(n4355), .Z(n1811) );
  MUX2_X1 U10952 ( .A(n1811), .B(n1810), .S(n4212), .Z(n1812) );
  MUX2_X1 U10953 ( .A(ram[3495]), .B(ram[3511]), .S(n4355), .Z(n1813) );
  MUX2_X1 U10954 ( .A(ram[3463]), .B(ram[3479]), .S(n4355), .Z(n1814) );
  MUX2_X1 U10955 ( .A(n1814), .B(n1813), .S(n4212), .Z(n1815) );
  MUX2_X1 U10956 ( .A(n1815), .B(n1812), .S(n4139), .Z(n1816) );
  MUX2_X1 U10957 ( .A(ram[3431]), .B(ram[3447]), .S(n4355), .Z(n1817) );
  MUX2_X1 U10958 ( .A(ram[3399]), .B(ram[3415]), .S(n4355), .Z(n1818) );
  MUX2_X1 U10959 ( .A(n1818), .B(n1817), .S(n4212), .Z(n1819) );
  MUX2_X1 U10960 ( .A(ram[3367]), .B(ram[3383]), .S(n4355), .Z(n1820) );
  MUX2_X1 U10961 ( .A(ram[3335]), .B(ram[3351]), .S(n4355), .Z(n1821) );
  MUX2_X1 U10962 ( .A(n1821), .B(n1820), .S(n4212), .Z(n1822) );
  MUX2_X1 U10963 ( .A(n1822), .B(n1819), .S(n4139), .Z(n1823) );
  MUX2_X1 U10964 ( .A(n1823), .B(n1816), .S(n4097), .Z(n1824) );
  MUX2_X1 U10965 ( .A(ram[3303]), .B(ram[3319]), .S(n4356), .Z(n1825) );
  MUX2_X1 U10966 ( .A(ram[3271]), .B(ram[3287]), .S(n4356), .Z(n1826) );
  MUX2_X1 U10967 ( .A(n1826), .B(n1825), .S(n4213), .Z(n1827) );
  MUX2_X1 U10968 ( .A(ram[3239]), .B(ram[3255]), .S(n4356), .Z(n1828) );
  MUX2_X1 U10969 ( .A(ram[3207]), .B(ram[3223]), .S(n4356), .Z(n1829) );
  MUX2_X1 U10970 ( .A(n1829), .B(n1828), .S(n4213), .Z(n1830) );
  MUX2_X1 U10971 ( .A(n1830), .B(n1827), .S(n4139), .Z(n1831) );
  MUX2_X1 U10972 ( .A(ram[3175]), .B(ram[3191]), .S(n4356), .Z(n1832) );
  MUX2_X1 U10973 ( .A(ram[3143]), .B(ram[3159]), .S(n4356), .Z(n1833) );
  MUX2_X1 U10974 ( .A(n1833), .B(n1832), .S(n4213), .Z(n1834) );
  MUX2_X1 U10975 ( .A(ram[3111]), .B(ram[3127]), .S(n4356), .Z(n1835) );
  MUX2_X1 U10976 ( .A(ram[3079]), .B(ram[3095]), .S(n4356), .Z(n1836) );
  MUX2_X1 U10977 ( .A(n1836), .B(n1835), .S(n4213), .Z(n1837) );
  MUX2_X1 U10978 ( .A(n1837), .B(n1834), .S(n4139), .Z(n1838) );
  MUX2_X1 U10979 ( .A(n1838), .B(n1831), .S(n4097), .Z(n1839) );
  MUX2_X1 U10980 ( .A(n1839), .B(n1824), .S(n4081), .Z(n1840) );
  MUX2_X1 U10981 ( .A(n1840), .B(n1809), .S(n4071), .Z(n1841) );
  MUX2_X1 U10982 ( .A(ram[3047]), .B(ram[3063]), .S(n4356), .Z(n1842) );
  MUX2_X1 U10983 ( .A(ram[3015]), .B(ram[3031]), .S(n4356), .Z(n1843) );
  MUX2_X1 U10984 ( .A(n1843), .B(n1842), .S(n4213), .Z(n1844) );
  MUX2_X1 U10985 ( .A(ram[2983]), .B(ram[2999]), .S(n4356), .Z(n1845) );
  MUX2_X1 U10986 ( .A(ram[2951]), .B(ram[2967]), .S(n4356), .Z(n1846) );
  MUX2_X1 U10987 ( .A(n1846), .B(n1845), .S(n4213), .Z(n1847) );
  MUX2_X1 U10988 ( .A(n1847), .B(n1844), .S(n4139), .Z(n1848) );
  MUX2_X1 U10989 ( .A(ram[2919]), .B(ram[2935]), .S(n8757), .Z(n1849) );
  MUX2_X1 U10990 ( .A(ram[2887]), .B(ram[2903]), .S(n8757), .Z(n1850) );
  MUX2_X1 U10991 ( .A(n1850), .B(n1849), .S(n4213), .Z(n1851) );
  MUX2_X1 U10992 ( .A(ram[2855]), .B(ram[2871]), .S(n8757), .Z(n1852) );
  MUX2_X1 U10993 ( .A(ram[2823]), .B(ram[2839]), .S(n8757), .Z(n1853) );
  MUX2_X1 U10994 ( .A(n1853), .B(n1852), .S(n4213), .Z(n1854) );
  MUX2_X1 U10995 ( .A(n1854), .B(n1851), .S(n4139), .Z(n1855) );
  MUX2_X1 U10996 ( .A(n1855), .B(n1848), .S(n4097), .Z(n1856) );
  MUX2_X1 U10997 ( .A(ram[2791]), .B(ram[2807]), .S(n8757), .Z(n1857) );
  MUX2_X1 U10998 ( .A(ram[2759]), .B(ram[2775]), .S(n8757), .Z(n1858) );
  MUX2_X1 U10999 ( .A(n1858), .B(n1857), .S(n4213), .Z(n1859) );
  MUX2_X1 U11000 ( .A(ram[2727]), .B(ram[2743]), .S(n8757), .Z(n1860) );
  MUX2_X1 U11001 ( .A(ram[2695]), .B(ram[2711]), .S(n8757), .Z(n1861) );
  MUX2_X1 U11002 ( .A(n1861), .B(n1860), .S(n4213), .Z(n1862) );
  MUX2_X1 U11003 ( .A(n1862), .B(n1859), .S(n4139), .Z(n1863) );
  MUX2_X1 U11004 ( .A(ram[2663]), .B(ram[2679]), .S(n8757), .Z(n1864) );
  MUX2_X1 U11005 ( .A(ram[2631]), .B(ram[2647]), .S(n8757), .Z(n1865) );
  MUX2_X1 U11006 ( .A(n1865), .B(n1864), .S(n4213), .Z(n1866) );
  MUX2_X1 U11007 ( .A(ram[2599]), .B(ram[2615]), .S(n8757), .Z(n1867) );
  MUX2_X1 U11008 ( .A(ram[2567]), .B(ram[2583]), .S(n8757), .Z(n1868) );
  MUX2_X1 U11009 ( .A(n1868), .B(n1867), .S(n4213), .Z(n1869) );
  MUX2_X1 U11010 ( .A(n1869), .B(n1866), .S(n4139), .Z(n1870) );
  MUX2_X1 U11011 ( .A(n1870), .B(n1863), .S(n4097), .Z(n1871) );
  MUX2_X1 U11012 ( .A(n1871), .B(n1856), .S(n4081), .Z(n1872) );
  MUX2_X1 U11013 ( .A(ram[2535]), .B(ram[2551]), .S(n8758), .Z(n1873) );
  MUX2_X1 U11014 ( .A(ram[2503]), .B(ram[2519]), .S(n8758), .Z(n1874) );
  MUX2_X1 U11015 ( .A(n1874), .B(n1873), .S(n4214), .Z(n1875) );
  MUX2_X1 U11016 ( .A(ram[2471]), .B(ram[2487]), .S(n8758), .Z(n1876) );
  MUX2_X1 U11017 ( .A(ram[2439]), .B(ram[2455]), .S(n8758), .Z(n1877) );
  MUX2_X1 U11018 ( .A(n1877), .B(n1876), .S(n4214), .Z(n1878) );
  MUX2_X1 U11019 ( .A(n1878), .B(n1875), .S(n4140), .Z(n1879) );
  MUX2_X1 U11020 ( .A(ram[2407]), .B(ram[2423]), .S(n8758), .Z(n1880) );
  MUX2_X1 U11021 ( .A(ram[2375]), .B(ram[2391]), .S(n8758), .Z(n1881) );
  MUX2_X1 U11022 ( .A(n1881), .B(n1880), .S(n4214), .Z(n1882) );
  MUX2_X1 U11023 ( .A(ram[2343]), .B(ram[2359]), .S(n8758), .Z(n1883) );
  MUX2_X1 U11024 ( .A(ram[2311]), .B(ram[2327]), .S(n8758), .Z(n1884) );
  MUX2_X1 U11025 ( .A(n1884), .B(n1883), .S(n4214), .Z(n1885) );
  MUX2_X1 U11026 ( .A(n1885), .B(n1882), .S(n4140), .Z(n1886) );
  MUX2_X1 U11027 ( .A(n1886), .B(n1879), .S(n4097), .Z(n1887) );
  MUX2_X1 U11028 ( .A(ram[2279]), .B(ram[2295]), .S(n8758), .Z(n1888) );
  MUX2_X1 U11029 ( .A(ram[2247]), .B(ram[2263]), .S(n8758), .Z(n1889) );
  MUX2_X1 U11030 ( .A(n1889), .B(n1888), .S(n4214), .Z(n1890) );
  MUX2_X1 U11031 ( .A(ram[2215]), .B(ram[2231]), .S(n8758), .Z(n1891) );
  MUX2_X1 U11032 ( .A(ram[2183]), .B(ram[2199]), .S(n8758), .Z(n1892) );
  MUX2_X1 U11033 ( .A(n1892), .B(n1891), .S(n4214), .Z(n1893) );
  MUX2_X1 U11034 ( .A(n1893), .B(n1890), .S(n4140), .Z(n1894) );
  MUX2_X1 U11035 ( .A(ram[2151]), .B(ram[2167]), .S(n8759), .Z(n1895) );
  MUX2_X1 U11036 ( .A(ram[2119]), .B(ram[2135]), .S(n8759), .Z(n1896) );
  MUX2_X1 U11037 ( .A(n1896), .B(n1895), .S(n4214), .Z(n1897) );
  MUX2_X1 U11038 ( .A(ram[2087]), .B(ram[2103]), .S(n8759), .Z(n1898) );
  MUX2_X1 U11039 ( .A(ram[2055]), .B(ram[2071]), .S(n8759), .Z(n1899) );
  MUX2_X1 U11040 ( .A(n1899), .B(n1898), .S(n4214), .Z(n1900) );
  MUX2_X1 U11041 ( .A(n1900), .B(n1897), .S(n4140), .Z(n1901) );
  MUX2_X1 U11042 ( .A(n1901), .B(n1894), .S(n4097), .Z(n1902) );
  MUX2_X1 U11043 ( .A(n1902), .B(n1887), .S(n4081), .Z(n1903) );
  MUX2_X1 U11044 ( .A(n1903), .B(n1872), .S(n4071), .Z(n1904) );
  MUX2_X1 U11045 ( .A(n1904), .B(n1841), .S(n4066), .Z(n1905) );
  MUX2_X1 U11046 ( .A(ram[2023]), .B(ram[2039]), .S(n8759), .Z(n1906) );
  MUX2_X1 U11047 ( .A(ram[1991]), .B(ram[2007]), .S(n8759), .Z(n1907) );
  MUX2_X1 U11048 ( .A(n1907), .B(n1906), .S(n4214), .Z(n1908) );
  MUX2_X1 U11049 ( .A(ram[1959]), .B(ram[1975]), .S(n8759), .Z(n1909) );
  MUX2_X1 U11050 ( .A(ram[1927]), .B(ram[1943]), .S(n8759), .Z(n1910) );
  MUX2_X1 U11051 ( .A(n1910), .B(n1909), .S(n4214), .Z(n1911) );
  MUX2_X1 U11052 ( .A(n1911), .B(n1908), .S(n4140), .Z(n1912) );
  MUX2_X1 U11053 ( .A(ram[1895]), .B(ram[1911]), .S(n8759), .Z(n1913) );
  MUX2_X1 U11054 ( .A(ram[1863]), .B(ram[1879]), .S(n8759), .Z(n1914) );
  MUX2_X1 U11055 ( .A(n1914), .B(n1913), .S(n4214), .Z(n1915) );
  MUX2_X1 U11056 ( .A(ram[1831]), .B(ram[1847]), .S(n8759), .Z(n1916) );
  MUX2_X1 U11057 ( .A(ram[1799]), .B(ram[1815]), .S(n8759), .Z(n1917) );
  MUX2_X1 U11058 ( .A(n1917), .B(n1916), .S(n4214), .Z(n1918) );
  MUX2_X1 U11059 ( .A(n1918), .B(n1915), .S(n4140), .Z(n1919) );
  MUX2_X1 U11060 ( .A(n1919), .B(n1912), .S(n4097), .Z(n1920) );
  MUX2_X1 U11061 ( .A(ram[1767]), .B(ram[1783]), .S(n8760), .Z(n1921) );
  MUX2_X1 U11062 ( .A(ram[1735]), .B(ram[1751]), .S(n8760), .Z(n1922) );
  MUX2_X1 U11063 ( .A(n1922), .B(n1921), .S(n4215), .Z(n1923) );
  MUX2_X1 U11064 ( .A(ram[1703]), .B(ram[1719]), .S(n8760), .Z(n1924) );
  MUX2_X1 U11065 ( .A(ram[1671]), .B(ram[1687]), .S(n8760), .Z(n1925) );
  MUX2_X1 U11066 ( .A(n1925), .B(n1924), .S(n4215), .Z(n1926) );
  MUX2_X1 U11067 ( .A(n1926), .B(n1923), .S(n4140), .Z(n1927) );
  MUX2_X1 U11068 ( .A(ram[1639]), .B(ram[1655]), .S(n8760), .Z(n1928) );
  MUX2_X1 U11069 ( .A(ram[1607]), .B(ram[1623]), .S(n8760), .Z(n1929) );
  MUX2_X1 U11070 ( .A(n1929), .B(n1928), .S(n4215), .Z(n1930) );
  MUX2_X1 U11071 ( .A(ram[1575]), .B(ram[1591]), .S(n8760), .Z(n1931) );
  MUX2_X1 U11072 ( .A(ram[1543]), .B(ram[1559]), .S(n8760), .Z(n1932) );
  MUX2_X1 U11073 ( .A(n1932), .B(n1931), .S(n4215), .Z(n1933) );
  MUX2_X1 U11074 ( .A(n1933), .B(n1930), .S(n4140), .Z(n1934) );
  MUX2_X1 U11075 ( .A(n1934), .B(n1927), .S(n4097), .Z(n1935) );
  MUX2_X1 U11076 ( .A(n1935), .B(n1920), .S(n4081), .Z(n1936) );
  MUX2_X1 U11077 ( .A(ram[1511]), .B(ram[1527]), .S(n8760), .Z(n1937) );
  MUX2_X1 U11078 ( .A(ram[1479]), .B(ram[1495]), .S(n8760), .Z(n1938) );
  MUX2_X1 U11079 ( .A(n1938), .B(n1937), .S(n4215), .Z(n1939) );
  MUX2_X1 U11080 ( .A(ram[1447]), .B(ram[1463]), .S(n8760), .Z(n1940) );
  MUX2_X1 U11081 ( .A(ram[1415]), .B(ram[1431]), .S(n8760), .Z(n1941) );
  MUX2_X1 U11082 ( .A(n1941), .B(n1940), .S(n4215), .Z(n1942) );
  MUX2_X1 U11083 ( .A(n1942), .B(n1939), .S(n4140), .Z(n1943) );
  MUX2_X1 U11084 ( .A(ram[1383]), .B(ram[1399]), .S(n8761), .Z(n1944) );
  MUX2_X1 U11085 ( .A(ram[1351]), .B(ram[1367]), .S(n8761), .Z(n1945) );
  MUX2_X1 U11086 ( .A(n1945), .B(n1944), .S(n4215), .Z(n1946) );
  MUX2_X1 U11087 ( .A(ram[1319]), .B(ram[1335]), .S(n8761), .Z(n1947) );
  MUX2_X1 U11088 ( .A(ram[1287]), .B(ram[1303]), .S(n8761), .Z(n1948) );
  MUX2_X1 U11089 ( .A(n1948), .B(n1947), .S(n4215), .Z(n1949) );
  MUX2_X1 U11090 ( .A(n1949), .B(n1946), .S(n4140), .Z(n1950) );
  MUX2_X1 U11091 ( .A(n1950), .B(n1943), .S(n4097), .Z(n1951) );
  MUX2_X1 U11092 ( .A(ram[1255]), .B(ram[1271]), .S(n8761), .Z(n1952) );
  MUX2_X1 U11093 ( .A(ram[1223]), .B(ram[1239]), .S(n8761), .Z(n1953) );
  MUX2_X1 U11094 ( .A(n1953), .B(n1952), .S(n4215), .Z(n1954) );
  MUX2_X1 U11095 ( .A(ram[1191]), .B(ram[1207]), .S(n8761), .Z(n1955) );
  MUX2_X1 U11096 ( .A(ram[1159]), .B(ram[1175]), .S(n8761), .Z(n1956) );
  MUX2_X1 U11097 ( .A(n1956), .B(n1955), .S(n4215), .Z(n1957) );
  MUX2_X1 U11098 ( .A(n1957), .B(n1954), .S(n4140), .Z(n1958) );
  MUX2_X1 U11099 ( .A(ram[1127]), .B(ram[1143]), .S(n8761), .Z(n1959) );
  MUX2_X1 U11100 ( .A(ram[1095]), .B(ram[1111]), .S(n8761), .Z(n1960) );
  MUX2_X1 U11101 ( .A(n1960), .B(n1959), .S(n4215), .Z(n1961) );
  MUX2_X1 U11102 ( .A(ram[1063]), .B(ram[1079]), .S(n8761), .Z(n1962) );
  MUX2_X1 U11103 ( .A(ram[1031]), .B(ram[1047]), .S(n8761), .Z(n1963) );
  MUX2_X1 U11104 ( .A(n1963), .B(n1962), .S(n4215), .Z(n1964) );
  MUX2_X1 U11105 ( .A(n1964), .B(n1961), .S(n4140), .Z(n1965) );
  MUX2_X1 U11106 ( .A(n1965), .B(n1958), .S(n4097), .Z(n1966) );
  MUX2_X1 U11107 ( .A(n1966), .B(n1951), .S(n4081), .Z(n1967) );
  MUX2_X1 U11108 ( .A(n1967), .B(n1936), .S(n4071), .Z(n1968) );
  MUX2_X1 U11109 ( .A(ram[999]), .B(ram[1015]), .S(n8762), .Z(n1969) );
  MUX2_X1 U11110 ( .A(ram[967]), .B(ram[983]), .S(n8762), .Z(n1970) );
  MUX2_X1 U11111 ( .A(n1970), .B(n1969), .S(n4216), .Z(n1971) );
  MUX2_X1 U11112 ( .A(ram[935]), .B(ram[951]), .S(n8762), .Z(n1972) );
  MUX2_X1 U11113 ( .A(ram[903]), .B(ram[919]), .S(n8762), .Z(n1973) );
  MUX2_X1 U11114 ( .A(n1973), .B(n1972), .S(n4216), .Z(n1974) );
  MUX2_X1 U11115 ( .A(n1974), .B(n1971), .S(n4141), .Z(n1975) );
  MUX2_X1 U11116 ( .A(ram[871]), .B(ram[887]), .S(n8762), .Z(n1976) );
  MUX2_X1 U11117 ( .A(ram[839]), .B(ram[855]), .S(n8762), .Z(n1977) );
  MUX2_X1 U11118 ( .A(n1977), .B(n1976), .S(n4216), .Z(n1978) );
  MUX2_X1 U11119 ( .A(ram[807]), .B(ram[823]), .S(n8762), .Z(n1979) );
  MUX2_X1 U11120 ( .A(ram[775]), .B(ram[791]), .S(n8762), .Z(n1980) );
  MUX2_X1 U11121 ( .A(n1980), .B(n1979), .S(n4216), .Z(n1981) );
  MUX2_X1 U11122 ( .A(n1981), .B(n1978), .S(n4141), .Z(n1982) );
  MUX2_X1 U11123 ( .A(n1982), .B(n1975), .S(n4098), .Z(n1983) );
  MUX2_X1 U11124 ( .A(ram[743]), .B(ram[759]), .S(n8762), .Z(n1984) );
  MUX2_X1 U11125 ( .A(ram[711]), .B(ram[727]), .S(n8762), .Z(n1985) );
  MUX2_X1 U11126 ( .A(n1985), .B(n1984), .S(n4216), .Z(n1986) );
  MUX2_X1 U11127 ( .A(ram[679]), .B(ram[695]), .S(n8762), .Z(n1987) );
  MUX2_X1 U11128 ( .A(ram[647]), .B(ram[663]), .S(n8762), .Z(n1988) );
  MUX2_X1 U11129 ( .A(n1988), .B(n1987), .S(n4216), .Z(n1989) );
  MUX2_X1 U11130 ( .A(n1989), .B(n1986), .S(n4141), .Z(n1990) );
  MUX2_X1 U11131 ( .A(ram[615]), .B(ram[631]), .S(n8763), .Z(n1991) );
  MUX2_X1 U11132 ( .A(ram[583]), .B(ram[599]), .S(n8763), .Z(n1992) );
  MUX2_X1 U11133 ( .A(n1992), .B(n1991), .S(n4216), .Z(n1993) );
  MUX2_X1 U11134 ( .A(ram[551]), .B(ram[567]), .S(n8763), .Z(n1994) );
  MUX2_X1 U11135 ( .A(ram[519]), .B(ram[535]), .S(n8763), .Z(n1995) );
  MUX2_X1 U11136 ( .A(n1995), .B(n1994), .S(n4216), .Z(n1996) );
  MUX2_X1 U11137 ( .A(n1996), .B(n1993), .S(n4141), .Z(n1997) );
  MUX2_X1 U11138 ( .A(n1997), .B(n1990), .S(n4098), .Z(n1998) );
  MUX2_X1 U11139 ( .A(n1998), .B(n1983), .S(n4081), .Z(n1999) );
  MUX2_X1 U11140 ( .A(ram[487]), .B(ram[503]), .S(n8763), .Z(n20001) );
  MUX2_X1 U11141 ( .A(ram[455]), .B(ram[471]), .S(n8763), .Z(n2001) );
  MUX2_X1 U11142 ( .A(n2001), .B(n20001), .S(n4216), .Z(n2002) );
  MUX2_X1 U11143 ( .A(ram[423]), .B(ram[439]), .S(n8763), .Z(n2003) );
  MUX2_X1 U11144 ( .A(ram[391]), .B(ram[407]), .S(n8763), .Z(n2004) );
  MUX2_X1 U11145 ( .A(n2004), .B(n2003), .S(n4216), .Z(n2005) );
  MUX2_X1 U11146 ( .A(n2005), .B(n2002), .S(n4141), .Z(n2006) );
  MUX2_X1 U11147 ( .A(ram[359]), .B(ram[375]), .S(n8763), .Z(n2007) );
  MUX2_X1 U11148 ( .A(ram[327]), .B(ram[343]), .S(n8763), .Z(n2008) );
  MUX2_X1 U11149 ( .A(n2008), .B(n2007), .S(n4216), .Z(n2009) );
  MUX2_X1 U11150 ( .A(ram[295]), .B(ram[311]), .S(n8763), .Z(n2010) );
  MUX2_X1 U11151 ( .A(ram[263]), .B(ram[279]), .S(n8763), .Z(n2011) );
  MUX2_X1 U11152 ( .A(n2011), .B(n2010), .S(n4216), .Z(n2012) );
  MUX2_X1 U11153 ( .A(n2012), .B(n2009), .S(n4141), .Z(n2013) );
  MUX2_X1 U11154 ( .A(n2013), .B(n2006), .S(n4098), .Z(n2014) );
  MUX2_X1 U11155 ( .A(ram[231]), .B(ram[247]), .S(n8764), .Z(n2015) );
  MUX2_X1 U11156 ( .A(ram[199]), .B(ram[215]), .S(n8764), .Z(n2016) );
  MUX2_X1 U11157 ( .A(n2016), .B(n2015), .S(n4217), .Z(n2017) );
  MUX2_X1 U11158 ( .A(ram[167]), .B(ram[183]), .S(n8764), .Z(n2018) );
  MUX2_X1 U11159 ( .A(ram[135]), .B(ram[151]), .S(n8764), .Z(n2019) );
  MUX2_X1 U11160 ( .A(n2019), .B(n2018), .S(n4217), .Z(n2020) );
  MUX2_X1 U11161 ( .A(n2020), .B(n2017), .S(n4141), .Z(n2021) );
  MUX2_X1 U11162 ( .A(ram[103]), .B(ram[119]), .S(n8764), .Z(n2022) );
  MUX2_X1 U11163 ( .A(ram[71]), .B(ram[87]), .S(n8764), .Z(n2023) );
  MUX2_X1 U11164 ( .A(n2023), .B(n2022), .S(n4217), .Z(n2024) );
  MUX2_X1 U11165 ( .A(ram[39]), .B(ram[55]), .S(n8764), .Z(n2025) );
  MUX2_X1 U11166 ( .A(ram[7]), .B(ram[23]), .S(n8764), .Z(n2026) );
  MUX2_X1 U11167 ( .A(n2026), .B(n2025), .S(n4217), .Z(n2027) );
  MUX2_X1 U11168 ( .A(n2027), .B(n2024), .S(n4141), .Z(n2028) );
  MUX2_X1 U11169 ( .A(n2028), .B(n2021), .S(n4098), .Z(n2029) );
  MUX2_X1 U11170 ( .A(n2029), .B(n2014), .S(n4081), .Z(n2030) );
  MUX2_X1 U11171 ( .A(n2030), .B(n1999), .S(n4071), .Z(n2031) );
  MUX2_X1 U11172 ( .A(n2031), .B(n1968), .S(n4066), .Z(n2032) );
  MUX2_X1 U11173 ( .A(n2032), .B(n1905), .S(mem_access_addr[9]), .Z(N294) );
  MUX2_X1 U11174 ( .A(ram[4072]), .B(ram[4088]), .S(n8764), .Z(n2033) );
  MUX2_X1 U11175 ( .A(ram[4040]), .B(ram[4056]), .S(n8764), .Z(n2034) );
  MUX2_X1 U11176 ( .A(n2034), .B(n2033), .S(n4217), .Z(n2035) );
  MUX2_X1 U11177 ( .A(ram[4008]), .B(ram[4024]), .S(n8764), .Z(n2036) );
  MUX2_X1 U11178 ( .A(ram[3976]), .B(ram[3992]), .S(n8764), .Z(n2037) );
  MUX2_X1 U11179 ( .A(n2037), .B(n2036), .S(n4217), .Z(n2038) );
  MUX2_X1 U11180 ( .A(n2038), .B(n2035), .S(n4141), .Z(n2039) );
  MUX2_X1 U11181 ( .A(ram[3944]), .B(ram[3960]), .S(n8765), .Z(n2040) );
  MUX2_X1 U11182 ( .A(ram[3912]), .B(ram[3928]), .S(n8765), .Z(n2041) );
  MUX2_X1 U11183 ( .A(n2041), .B(n2040), .S(n4217), .Z(n2042) );
  MUX2_X1 U11184 ( .A(ram[3880]), .B(ram[3896]), .S(n8765), .Z(n2043) );
  MUX2_X1 U11185 ( .A(ram[3848]), .B(ram[3864]), .S(n8765), .Z(n2044) );
  MUX2_X1 U11186 ( .A(n2044), .B(n2043), .S(n4217), .Z(n2045) );
  MUX2_X1 U11187 ( .A(n2045), .B(n2042), .S(n4141), .Z(n2046) );
  MUX2_X1 U11188 ( .A(n2046), .B(n2039), .S(n4098), .Z(n2047) );
  MUX2_X1 U11189 ( .A(ram[3816]), .B(ram[3832]), .S(n8765), .Z(n2048) );
  MUX2_X1 U11190 ( .A(ram[3784]), .B(ram[3800]), .S(n8765), .Z(n2049) );
  MUX2_X1 U11191 ( .A(n2049), .B(n2048), .S(n4217), .Z(n2050) );
  MUX2_X1 U11192 ( .A(ram[3752]), .B(ram[3768]), .S(n8765), .Z(n2051) );
  MUX2_X1 U11193 ( .A(ram[3720]), .B(ram[3736]), .S(n8765), .Z(n2052) );
  MUX2_X1 U11194 ( .A(n2052), .B(n2051), .S(n4217), .Z(n2053) );
  MUX2_X1 U11195 ( .A(n2053), .B(n2050), .S(n4141), .Z(n2054) );
  MUX2_X1 U11196 ( .A(ram[3688]), .B(ram[3704]), .S(n8765), .Z(n2055) );
  MUX2_X1 U11197 ( .A(ram[3656]), .B(ram[3672]), .S(n8765), .Z(n2056) );
  MUX2_X1 U11198 ( .A(n2056), .B(n2055), .S(n4217), .Z(n2057) );
  MUX2_X1 U11199 ( .A(ram[3624]), .B(ram[3640]), .S(n8765), .Z(n2058) );
  MUX2_X1 U11200 ( .A(ram[3592]), .B(ram[3608]), .S(n8765), .Z(n2059) );
  MUX2_X1 U11201 ( .A(n2059), .B(n2058), .S(n4217), .Z(n2060) );
  MUX2_X1 U11202 ( .A(n2060), .B(n2057), .S(n4141), .Z(n2061) );
  MUX2_X1 U11203 ( .A(n2061), .B(n2054), .S(n4098), .Z(n2062) );
  MUX2_X1 U11204 ( .A(n2062), .B(n2047), .S(n4081), .Z(n2063) );
  MUX2_X1 U11205 ( .A(ram[3560]), .B(ram[3576]), .S(n8766), .Z(n2064) );
  MUX2_X1 U11206 ( .A(ram[3528]), .B(ram[3544]), .S(n8766), .Z(n2065) );
  MUX2_X1 U11207 ( .A(n2065), .B(n2064), .S(n4218), .Z(n2066) );
  MUX2_X1 U11208 ( .A(ram[3496]), .B(ram[3512]), .S(n8766), .Z(n2067) );
  MUX2_X1 U11209 ( .A(ram[3464]), .B(ram[3480]), .S(n8766), .Z(n2068) );
  MUX2_X1 U11210 ( .A(n2068), .B(n2067), .S(n4218), .Z(n2069) );
  MUX2_X1 U11211 ( .A(n2069), .B(n2066), .S(n4142), .Z(n2070) );
  MUX2_X1 U11212 ( .A(ram[3432]), .B(ram[3448]), .S(n8766), .Z(n2071) );
  MUX2_X1 U11213 ( .A(ram[3400]), .B(ram[3416]), .S(n8766), .Z(n2072) );
  MUX2_X1 U11214 ( .A(n2072), .B(n2071), .S(n4218), .Z(n2073) );
  MUX2_X1 U11215 ( .A(ram[3368]), .B(ram[3384]), .S(n8766), .Z(n2074) );
  MUX2_X1 U11216 ( .A(ram[3336]), .B(ram[3352]), .S(n8766), .Z(n2075) );
  MUX2_X1 U11217 ( .A(n2075), .B(n2074), .S(n4218), .Z(n2076) );
  MUX2_X1 U11218 ( .A(n2076), .B(n2073), .S(n4142), .Z(n2077) );
  MUX2_X1 U11219 ( .A(n2077), .B(n2070), .S(n4098), .Z(n2078) );
  MUX2_X1 U11220 ( .A(ram[3304]), .B(ram[3320]), .S(n8766), .Z(n2079) );
  MUX2_X1 U11221 ( .A(ram[3272]), .B(ram[3288]), .S(n8766), .Z(n2080) );
  MUX2_X1 U11222 ( .A(n2080), .B(n2079), .S(n4218), .Z(n2081) );
  MUX2_X1 U11223 ( .A(ram[3240]), .B(ram[3256]), .S(n8766), .Z(n2082) );
  MUX2_X1 U11224 ( .A(ram[3208]), .B(ram[3224]), .S(n8766), .Z(n2083) );
  MUX2_X1 U11225 ( .A(n2083), .B(n2082), .S(n4218), .Z(n2084) );
  MUX2_X1 U11226 ( .A(n2084), .B(n2081), .S(n4142), .Z(n2085) );
  MUX2_X1 U11227 ( .A(ram[3176]), .B(ram[3192]), .S(n8767), .Z(n2086) );
  MUX2_X1 U11228 ( .A(ram[3144]), .B(ram[3160]), .S(n8767), .Z(n2087) );
  MUX2_X1 U11229 ( .A(n2087), .B(n2086), .S(n4218), .Z(n2088) );
  MUX2_X1 U11230 ( .A(ram[3112]), .B(ram[3128]), .S(n8767), .Z(n2089) );
  MUX2_X1 U11231 ( .A(ram[3080]), .B(ram[3096]), .S(n8767), .Z(n2090) );
  MUX2_X1 U11232 ( .A(n2090), .B(n2089), .S(n4218), .Z(n2091) );
  MUX2_X1 U11233 ( .A(n2091), .B(n2088), .S(n4142), .Z(n2092) );
  MUX2_X1 U11234 ( .A(n2092), .B(n2085), .S(n4098), .Z(n2093) );
  MUX2_X1 U11235 ( .A(n2093), .B(n2078), .S(n4081), .Z(n2094) );
  MUX2_X1 U11236 ( .A(n2094), .B(n2063), .S(n4071), .Z(n2095) );
  MUX2_X1 U11237 ( .A(ram[3048]), .B(ram[3064]), .S(n8767), .Z(n2096) );
  MUX2_X1 U11238 ( .A(ram[3016]), .B(ram[3032]), .S(n8767), .Z(n2097) );
  MUX2_X1 U11239 ( .A(n2097), .B(n2096), .S(n4218), .Z(n2098) );
  MUX2_X1 U11240 ( .A(ram[2984]), .B(ram[3000]), .S(n8767), .Z(n2099) );
  MUX2_X1 U11241 ( .A(ram[2952]), .B(ram[2968]), .S(n8767), .Z(n21001) );
  MUX2_X1 U11242 ( .A(n21001), .B(n2099), .S(n4218), .Z(n2101) );
  MUX2_X1 U11243 ( .A(n2101), .B(n2098), .S(n4142), .Z(n2102) );
  MUX2_X1 U11244 ( .A(ram[2920]), .B(ram[2936]), .S(n8767), .Z(n2103) );
  MUX2_X1 U11245 ( .A(ram[2888]), .B(ram[2904]), .S(n8767), .Z(n2104) );
  MUX2_X1 U11246 ( .A(n2104), .B(n2103), .S(n4218), .Z(n2105) );
  MUX2_X1 U11247 ( .A(ram[2856]), .B(ram[2872]), .S(n8767), .Z(n2106) );
  MUX2_X1 U11248 ( .A(ram[2824]), .B(ram[2840]), .S(n8767), .Z(n2107) );
  MUX2_X1 U11249 ( .A(n2107), .B(n2106), .S(n4218), .Z(n2108) );
  MUX2_X1 U11250 ( .A(n2108), .B(n2105), .S(n4142), .Z(n2109) );
  MUX2_X1 U11251 ( .A(n2109), .B(n2102), .S(n4098), .Z(n2110) );
  MUX2_X1 U11252 ( .A(ram[2792]), .B(ram[2808]), .S(n8768), .Z(n2111) );
  MUX2_X1 U11253 ( .A(ram[2760]), .B(ram[2776]), .S(n8768), .Z(n2112) );
  MUX2_X1 U11254 ( .A(n2112), .B(n2111), .S(n4219), .Z(n2113) );
  MUX2_X1 U11255 ( .A(ram[2728]), .B(ram[2744]), .S(n8768), .Z(n2114) );
  MUX2_X1 U11256 ( .A(ram[2696]), .B(ram[2712]), .S(n8768), .Z(n2115) );
  MUX2_X1 U11257 ( .A(n2115), .B(n2114), .S(n4219), .Z(n2116) );
  MUX2_X1 U11258 ( .A(n2116), .B(n2113), .S(n4142), .Z(n2117) );
  MUX2_X1 U11259 ( .A(ram[2664]), .B(ram[2680]), .S(n8768), .Z(n2118) );
  MUX2_X1 U11260 ( .A(ram[2632]), .B(ram[2648]), .S(n8768), .Z(n2119) );
  MUX2_X1 U11261 ( .A(n2119), .B(n2118), .S(n4219), .Z(n2120) );
  MUX2_X1 U11262 ( .A(ram[2600]), .B(ram[2616]), .S(n8768), .Z(n2121) );
  MUX2_X1 U11263 ( .A(ram[2568]), .B(ram[2584]), .S(n8768), .Z(n2122) );
  MUX2_X1 U11264 ( .A(n2122), .B(n2121), .S(n4219), .Z(n2123) );
  MUX2_X1 U11265 ( .A(n2123), .B(n2120), .S(n4142), .Z(n2124) );
  MUX2_X1 U11266 ( .A(n2124), .B(n2117), .S(n4098), .Z(n2125) );
  MUX2_X1 U11267 ( .A(n2125), .B(n2110), .S(n4081), .Z(n2126) );
  MUX2_X1 U11268 ( .A(ram[2536]), .B(ram[2552]), .S(n8768), .Z(n2127) );
  MUX2_X1 U11269 ( .A(ram[2504]), .B(ram[2520]), .S(n8768), .Z(n2128) );
  MUX2_X1 U11270 ( .A(n2128), .B(n2127), .S(n4219), .Z(n2129) );
  MUX2_X1 U11271 ( .A(ram[2472]), .B(ram[2488]), .S(n8768), .Z(n2130) );
  MUX2_X1 U11272 ( .A(ram[2440]), .B(ram[2456]), .S(n8768), .Z(n2131) );
  MUX2_X1 U11273 ( .A(n2131), .B(n2130), .S(n4219), .Z(n2132) );
  MUX2_X1 U11274 ( .A(n2132), .B(n2129), .S(n4142), .Z(n2133) );
  MUX2_X1 U11275 ( .A(ram[2408]), .B(ram[2424]), .S(n8769), .Z(n2134) );
  MUX2_X1 U11276 ( .A(ram[2376]), .B(ram[2392]), .S(n8769), .Z(n2135) );
  MUX2_X1 U11277 ( .A(n2135), .B(n2134), .S(n4219), .Z(n2136) );
  MUX2_X1 U11278 ( .A(ram[2344]), .B(ram[2360]), .S(n8769), .Z(n2137) );
  MUX2_X1 U11279 ( .A(ram[2312]), .B(ram[2328]), .S(n8769), .Z(n2138) );
  MUX2_X1 U11280 ( .A(n2138), .B(n2137), .S(n4219), .Z(n2139) );
  MUX2_X1 U11281 ( .A(n2139), .B(n2136), .S(n4142), .Z(n2140) );
  MUX2_X1 U11282 ( .A(n2140), .B(n2133), .S(n4098), .Z(n2141) );
  MUX2_X1 U11283 ( .A(ram[2280]), .B(ram[2296]), .S(n8769), .Z(n2142) );
  MUX2_X1 U11284 ( .A(ram[2248]), .B(ram[2264]), .S(n8769), .Z(n2143) );
  MUX2_X1 U11285 ( .A(n2143), .B(n2142), .S(n4219), .Z(n2144) );
  MUX2_X1 U11286 ( .A(ram[2216]), .B(ram[2232]), .S(n8769), .Z(n2145) );
  MUX2_X1 U11287 ( .A(ram[2184]), .B(ram[2200]), .S(n8769), .Z(n2146) );
  MUX2_X1 U11288 ( .A(n2146), .B(n2145), .S(n4219), .Z(n2147) );
  MUX2_X1 U11289 ( .A(n2147), .B(n2144), .S(n4142), .Z(n2148) );
  MUX2_X1 U11290 ( .A(ram[2152]), .B(ram[2168]), .S(n8769), .Z(n2149) );
  MUX2_X1 U11291 ( .A(ram[2120]), .B(ram[2136]), .S(n8769), .Z(n2150) );
  MUX2_X1 U11292 ( .A(n2150), .B(n2149), .S(n4219), .Z(n2151) );
  MUX2_X1 U11293 ( .A(ram[2088]), .B(ram[2104]), .S(n8769), .Z(n2152) );
  MUX2_X1 U11294 ( .A(ram[2056]), .B(ram[2072]), .S(n8769), .Z(n2153) );
  MUX2_X1 U11295 ( .A(n2153), .B(n2152), .S(n4219), .Z(n2154) );
  MUX2_X1 U11296 ( .A(n2154), .B(n2151), .S(n4142), .Z(n2155) );
  MUX2_X1 U11297 ( .A(n2155), .B(n2148), .S(n4098), .Z(n2156) );
  MUX2_X1 U11298 ( .A(n2156), .B(n2141), .S(n4081), .Z(n2157) );
  MUX2_X1 U11299 ( .A(n2157), .B(n2126), .S(n4071), .Z(n2158) );
  MUX2_X1 U11300 ( .A(n2158), .B(n2095), .S(n4066), .Z(n2159) );
  MUX2_X1 U11301 ( .A(ram[2024]), .B(ram[2040]), .S(n8770), .Z(n2160) );
  MUX2_X1 U11302 ( .A(ram[1992]), .B(ram[2008]), .S(n8770), .Z(n2161) );
  MUX2_X1 U11303 ( .A(n2161), .B(n2160), .S(n4220), .Z(n2162) );
  MUX2_X1 U11304 ( .A(ram[1960]), .B(ram[1976]), .S(n8770), .Z(n2163) );
  MUX2_X1 U11305 ( .A(ram[1928]), .B(ram[1944]), .S(n8770), .Z(n2164) );
  MUX2_X1 U11306 ( .A(n2164), .B(n2163), .S(n4220), .Z(n2165) );
  MUX2_X1 U11307 ( .A(n2165), .B(n2162), .S(n4143), .Z(n2166) );
  MUX2_X1 U11308 ( .A(ram[1896]), .B(ram[1912]), .S(n8770), .Z(n2167) );
  MUX2_X1 U11309 ( .A(ram[1864]), .B(ram[1880]), .S(n8770), .Z(n2168) );
  MUX2_X1 U11310 ( .A(n2168), .B(n2167), .S(n4220), .Z(n2169) );
  MUX2_X1 U11311 ( .A(ram[1832]), .B(ram[1848]), .S(n8770), .Z(n2170) );
  MUX2_X1 U11312 ( .A(ram[1800]), .B(ram[1816]), .S(n8770), .Z(n2171) );
  MUX2_X1 U11313 ( .A(n2171), .B(n2170), .S(n4220), .Z(n2172) );
  MUX2_X1 U11314 ( .A(n2172), .B(n2169), .S(n4143), .Z(n2173) );
  MUX2_X1 U11315 ( .A(n2173), .B(n2166), .S(n4099), .Z(n2174) );
  MUX2_X1 U11316 ( .A(ram[1768]), .B(ram[1784]), .S(n8770), .Z(n2175) );
  MUX2_X1 U11317 ( .A(ram[1736]), .B(ram[1752]), .S(n8770), .Z(n2176) );
  MUX2_X1 U11318 ( .A(n2176), .B(n2175), .S(n4220), .Z(n2177) );
  MUX2_X1 U11319 ( .A(ram[1704]), .B(ram[1720]), .S(n8770), .Z(n2178) );
  MUX2_X1 U11320 ( .A(ram[1672]), .B(ram[1688]), .S(n8770), .Z(n2179) );
  MUX2_X1 U11321 ( .A(n2179), .B(n2178), .S(n4220), .Z(n2180) );
  MUX2_X1 U11322 ( .A(n2180), .B(n2177), .S(n4143), .Z(n2181) );
  MUX2_X1 U11323 ( .A(ram[1640]), .B(ram[1656]), .S(n8771), .Z(n2182) );
  MUX2_X1 U11324 ( .A(ram[1608]), .B(ram[1624]), .S(n8771), .Z(n2183) );
  MUX2_X1 U11325 ( .A(n2183), .B(n2182), .S(n4220), .Z(n2184) );
  MUX2_X1 U11326 ( .A(ram[1576]), .B(ram[1592]), .S(n8771), .Z(n2185) );
  MUX2_X1 U11327 ( .A(ram[1544]), .B(ram[1560]), .S(n8771), .Z(n2186) );
  MUX2_X1 U11328 ( .A(n2186), .B(n2185), .S(n4220), .Z(n2187) );
  MUX2_X1 U11329 ( .A(n2187), .B(n2184), .S(n4143), .Z(n2188) );
  MUX2_X1 U11330 ( .A(n2188), .B(n2181), .S(n4099), .Z(n2189) );
  MUX2_X1 U11331 ( .A(n2189), .B(n2174), .S(n4082), .Z(n2190) );
  MUX2_X1 U11332 ( .A(ram[1512]), .B(ram[1528]), .S(n8771), .Z(n2191) );
  MUX2_X1 U11333 ( .A(ram[1480]), .B(ram[1496]), .S(n8771), .Z(n2192) );
  MUX2_X1 U11334 ( .A(n2192), .B(n2191), .S(n4220), .Z(n2193) );
  MUX2_X1 U11335 ( .A(ram[1448]), .B(ram[1464]), .S(n8771), .Z(n2194) );
  MUX2_X1 U11336 ( .A(ram[1416]), .B(ram[1432]), .S(n8771), .Z(n2195) );
  MUX2_X1 U11337 ( .A(n2195), .B(n2194), .S(n4220), .Z(n2196) );
  MUX2_X1 U11338 ( .A(n2196), .B(n2193), .S(n4143), .Z(n2197) );
  MUX2_X1 U11339 ( .A(ram[1384]), .B(ram[1400]), .S(n8771), .Z(n2198) );
  MUX2_X1 U11340 ( .A(ram[1352]), .B(ram[1368]), .S(n8771), .Z(n2199) );
  MUX2_X1 U11341 ( .A(n2199), .B(n2198), .S(n4220), .Z(n22001) );
  MUX2_X1 U11342 ( .A(ram[1320]), .B(ram[1336]), .S(n8771), .Z(n2201) );
  MUX2_X1 U11343 ( .A(ram[1288]), .B(ram[1304]), .S(n8771), .Z(n2202) );
  MUX2_X1 U11344 ( .A(n2202), .B(n2201), .S(n4220), .Z(n2203) );
  MUX2_X1 U11345 ( .A(n2203), .B(n22001), .S(n4143), .Z(n2204) );
  MUX2_X1 U11346 ( .A(n2204), .B(n2197), .S(n4099), .Z(n2205) );
  MUX2_X1 U11347 ( .A(ram[1256]), .B(ram[1272]), .S(n8772), .Z(n2206) );
  MUX2_X1 U11348 ( .A(ram[1224]), .B(ram[1240]), .S(n8772), .Z(n2207) );
  MUX2_X1 U11349 ( .A(n2207), .B(n2206), .S(n4221), .Z(n2208) );
  MUX2_X1 U11350 ( .A(ram[1192]), .B(ram[1208]), .S(n8772), .Z(n2209) );
  MUX2_X1 U11351 ( .A(ram[1160]), .B(ram[1176]), .S(n8772), .Z(n2210) );
  MUX2_X1 U11352 ( .A(n2210), .B(n2209), .S(n4221), .Z(n2211) );
  MUX2_X1 U11353 ( .A(n2211), .B(n2208), .S(n4143), .Z(n2212) );
  MUX2_X1 U11354 ( .A(ram[1128]), .B(ram[1144]), .S(n8772), .Z(n2213) );
  MUX2_X1 U11355 ( .A(ram[1096]), .B(ram[1112]), .S(n8772), .Z(n2214) );
  MUX2_X1 U11356 ( .A(n2214), .B(n2213), .S(n4221), .Z(n2215) );
  MUX2_X1 U11357 ( .A(ram[1064]), .B(ram[1080]), .S(n8772), .Z(n2216) );
  MUX2_X1 U11358 ( .A(ram[1032]), .B(ram[1048]), .S(n8772), .Z(n2217) );
  MUX2_X1 U11359 ( .A(n2217), .B(n2216), .S(n4221), .Z(n2218) );
  MUX2_X1 U11360 ( .A(n2218), .B(n2215), .S(n4143), .Z(n2219) );
  MUX2_X1 U11361 ( .A(n2219), .B(n2212), .S(n4099), .Z(n2220) );
  MUX2_X1 U11362 ( .A(n2220), .B(n2205), .S(n4082), .Z(n2221) );
  MUX2_X1 U11363 ( .A(n2221), .B(n2190), .S(n4071), .Z(n2222) );
  MUX2_X1 U11364 ( .A(ram[1000]), .B(ram[1016]), .S(n8772), .Z(n2223) );
  MUX2_X1 U11365 ( .A(ram[968]), .B(ram[984]), .S(n8772), .Z(n2224) );
  MUX2_X1 U11366 ( .A(n2224), .B(n2223), .S(n4221), .Z(n2225) );
  MUX2_X1 U11367 ( .A(ram[936]), .B(ram[952]), .S(n8772), .Z(n2226) );
  MUX2_X1 U11368 ( .A(ram[904]), .B(ram[920]), .S(n8772), .Z(n2227) );
  MUX2_X1 U11369 ( .A(n2227), .B(n2226), .S(n4221), .Z(n2228) );
  MUX2_X1 U11370 ( .A(n2228), .B(n2225), .S(n4143), .Z(n2229) );
  MUX2_X1 U11371 ( .A(ram[872]), .B(ram[888]), .S(n8773), .Z(n2230) );
  MUX2_X1 U11372 ( .A(ram[840]), .B(ram[856]), .S(n8773), .Z(n2231) );
  MUX2_X1 U11373 ( .A(n2231), .B(n2230), .S(n4221), .Z(n2232) );
  MUX2_X1 U11374 ( .A(ram[808]), .B(ram[824]), .S(n8773), .Z(n2233) );
  MUX2_X1 U11375 ( .A(ram[776]), .B(ram[792]), .S(n8773), .Z(n2234) );
  MUX2_X1 U11376 ( .A(n2234), .B(n2233), .S(n4221), .Z(n2235) );
  MUX2_X1 U11377 ( .A(n2235), .B(n2232), .S(n4143), .Z(n2236) );
  MUX2_X1 U11378 ( .A(n2236), .B(n2229), .S(n4099), .Z(n2237) );
  MUX2_X1 U11379 ( .A(ram[744]), .B(ram[760]), .S(n8773), .Z(n2238) );
  MUX2_X1 U11380 ( .A(ram[712]), .B(ram[728]), .S(n8773), .Z(n2239) );
  MUX2_X1 U11381 ( .A(n2239), .B(n2238), .S(n4221), .Z(n2240) );
  MUX2_X1 U11382 ( .A(ram[680]), .B(ram[696]), .S(n8773), .Z(n2241) );
  MUX2_X1 U11383 ( .A(ram[648]), .B(ram[664]), .S(n8773), .Z(n2242) );
  MUX2_X1 U11384 ( .A(n2242), .B(n2241), .S(n4221), .Z(n2243) );
  MUX2_X1 U11385 ( .A(n2243), .B(n2240), .S(n4143), .Z(n2244) );
  MUX2_X1 U11386 ( .A(ram[616]), .B(ram[632]), .S(n8773), .Z(n2245) );
  MUX2_X1 U11387 ( .A(ram[584]), .B(ram[600]), .S(n8773), .Z(n2246) );
  MUX2_X1 U11388 ( .A(n2246), .B(n2245), .S(n4221), .Z(n2247) );
  MUX2_X1 U11389 ( .A(ram[552]), .B(ram[568]), .S(n8773), .Z(n2248) );
  MUX2_X1 U11390 ( .A(ram[520]), .B(ram[536]), .S(n8773), .Z(n2249) );
  MUX2_X1 U11391 ( .A(n2249), .B(n2248), .S(n4221), .Z(n2250) );
  MUX2_X1 U11392 ( .A(n2250), .B(n2247), .S(n4143), .Z(n2251) );
  MUX2_X1 U11393 ( .A(n2251), .B(n2244), .S(n4099), .Z(n2252) );
  MUX2_X1 U11394 ( .A(n2252), .B(n2237), .S(n4082), .Z(n2253) );
  MUX2_X1 U11395 ( .A(ram[488]), .B(ram[504]), .S(n8774), .Z(n2254) );
  MUX2_X1 U11396 ( .A(ram[456]), .B(ram[472]), .S(n8774), .Z(n2255) );
  MUX2_X1 U11397 ( .A(n2255), .B(n2254), .S(n4222), .Z(n2256) );
  MUX2_X1 U11398 ( .A(ram[424]), .B(ram[440]), .S(n8774), .Z(n2257) );
  MUX2_X1 U11399 ( .A(ram[392]), .B(ram[408]), .S(n8774), .Z(n2258) );
  MUX2_X1 U11400 ( .A(n2258), .B(n2257), .S(n4222), .Z(n2259) );
  MUX2_X1 U11401 ( .A(n2259), .B(n2256), .S(n4144), .Z(n2260) );
  MUX2_X1 U11402 ( .A(ram[360]), .B(ram[376]), .S(n8774), .Z(n2261) );
  MUX2_X1 U11403 ( .A(ram[328]), .B(ram[344]), .S(n8774), .Z(n2262) );
  MUX2_X1 U11404 ( .A(n2262), .B(n2261), .S(n4222), .Z(n2263) );
  MUX2_X1 U11405 ( .A(ram[296]), .B(ram[312]), .S(n8774), .Z(n2264) );
  MUX2_X1 U11406 ( .A(ram[264]), .B(ram[280]), .S(n8774), .Z(n2265) );
  MUX2_X1 U11407 ( .A(n2265), .B(n2264), .S(n4222), .Z(n2266) );
  MUX2_X1 U11408 ( .A(n2266), .B(n2263), .S(n4144), .Z(n2267) );
  MUX2_X1 U11409 ( .A(n2267), .B(n2260), .S(n4099), .Z(n2268) );
  MUX2_X1 U11410 ( .A(ram[232]), .B(ram[248]), .S(n8774), .Z(n2269) );
  MUX2_X1 U11411 ( .A(ram[200]), .B(ram[216]), .S(n8774), .Z(n2270) );
  MUX2_X1 U11412 ( .A(n2270), .B(n2269), .S(n4222), .Z(n2271) );
  MUX2_X1 U11413 ( .A(ram[168]), .B(ram[184]), .S(n8774), .Z(n2272) );
  MUX2_X1 U11414 ( .A(ram[136]), .B(ram[152]), .S(n8774), .Z(n2273) );
  MUX2_X1 U11415 ( .A(n2273), .B(n2272), .S(n4222), .Z(n2274) );
  MUX2_X1 U11416 ( .A(n2274), .B(n2271), .S(n4144), .Z(n2275) );
  MUX2_X1 U11417 ( .A(ram[104]), .B(ram[120]), .S(n8775), .Z(n2276) );
  MUX2_X1 U11418 ( .A(ram[72]), .B(ram[88]), .S(n8775), .Z(n2277) );
  MUX2_X1 U11419 ( .A(n2277), .B(n2276), .S(n4222), .Z(n2278) );
  MUX2_X1 U11420 ( .A(ram[40]), .B(ram[56]), .S(n8775), .Z(n2279) );
  MUX2_X1 U11421 ( .A(ram[8]), .B(ram[24]), .S(n8775), .Z(n2280) );
  MUX2_X1 U11422 ( .A(n2280), .B(n2279), .S(n4222), .Z(n2281) );
  MUX2_X1 U11423 ( .A(n2281), .B(n2278), .S(n4144), .Z(n2282) );
  MUX2_X1 U11424 ( .A(n2282), .B(n2275), .S(n4099), .Z(n2283) );
  MUX2_X1 U11425 ( .A(n2283), .B(n2268), .S(n4082), .Z(n2284) );
  MUX2_X1 U11426 ( .A(n2284), .B(n2253), .S(n4071), .Z(n2285) );
  MUX2_X1 U11427 ( .A(n2285), .B(n2222), .S(n4066), .Z(n2286) );
  MUX2_X1 U11428 ( .A(n2286), .B(n2159), .S(mem_access_addr[9]), .Z(N293) );
  MUX2_X1 U11429 ( .A(ram[4073]), .B(ram[4089]), .S(n8775), .Z(n2287) );
  MUX2_X1 U11430 ( .A(ram[4041]), .B(ram[4057]), .S(n8775), .Z(n2288) );
  MUX2_X1 U11431 ( .A(n2288), .B(n2287), .S(n4222), .Z(n2289) );
  MUX2_X1 U11432 ( .A(ram[4009]), .B(ram[4025]), .S(n8775), .Z(n2290) );
  MUX2_X1 U11433 ( .A(ram[3977]), .B(ram[3993]), .S(n8775), .Z(n2291) );
  MUX2_X1 U11434 ( .A(n2291), .B(n2290), .S(n4222), .Z(n2292) );
  MUX2_X1 U11435 ( .A(n2292), .B(n2289), .S(n4144), .Z(n2293) );
  MUX2_X1 U11436 ( .A(ram[3945]), .B(ram[3961]), .S(n8775), .Z(n2294) );
  MUX2_X1 U11437 ( .A(ram[3913]), .B(ram[3929]), .S(n8775), .Z(n2295) );
  MUX2_X1 U11438 ( .A(n2295), .B(n2294), .S(n4222), .Z(n2296) );
  MUX2_X1 U11439 ( .A(ram[3881]), .B(ram[3897]), .S(n8775), .Z(n2297) );
  MUX2_X1 U11440 ( .A(ram[3849]), .B(ram[3865]), .S(n8775), .Z(n2298) );
  MUX2_X1 U11441 ( .A(n2298), .B(n2297), .S(n4222), .Z(n2299) );
  MUX2_X1 U11442 ( .A(n2299), .B(n2296), .S(n4144), .Z(n23001) );
  MUX2_X1 U11443 ( .A(n23001), .B(n2293), .S(n4099), .Z(n2301) );
  MUX2_X1 U11444 ( .A(ram[3817]), .B(ram[3833]), .S(n8776), .Z(n2302) );
  MUX2_X1 U11445 ( .A(ram[3785]), .B(ram[3801]), .S(n8776), .Z(n2303) );
  MUX2_X1 U11446 ( .A(n2303), .B(n2302), .S(n4223), .Z(n2304) );
  MUX2_X1 U11447 ( .A(ram[3753]), .B(ram[3769]), .S(n8776), .Z(n2305) );
  MUX2_X1 U11448 ( .A(ram[3721]), .B(ram[3737]), .S(n8776), .Z(n2306) );
  MUX2_X1 U11449 ( .A(n2306), .B(n2305), .S(n4223), .Z(n2307) );
  MUX2_X1 U11450 ( .A(n2307), .B(n2304), .S(n4144), .Z(n2308) );
  MUX2_X1 U11451 ( .A(ram[3689]), .B(ram[3705]), .S(n8776), .Z(n2309) );
  MUX2_X1 U11452 ( .A(ram[3657]), .B(ram[3673]), .S(n8776), .Z(n2310) );
  MUX2_X1 U11453 ( .A(n2310), .B(n2309), .S(n4223), .Z(n2311) );
  MUX2_X1 U11454 ( .A(ram[3625]), .B(ram[3641]), .S(n8776), .Z(n2312) );
  MUX2_X1 U11455 ( .A(ram[3593]), .B(ram[3609]), .S(n8776), .Z(n2313) );
  MUX2_X1 U11456 ( .A(n2313), .B(n2312), .S(n4223), .Z(n2314) );
  MUX2_X1 U11457 ( .A(n2314), .B(n2311), .S(n4144), .Z(n2315) );
  MUX2_X1 U11458 ( .A(n2315), .B(n2308), .S(n4099), .Z(n2316) );
  MUX2_X1 U11459 ( .A(n2316), .B(n2301), .S(n4082), .Z(n2317) );
  MUX2_X1 U11460 ( .A(ram[3561]), .B(ram[3577]), .S(n8776), .Z(n2318) );
  MUX2_X1 U11461 ( .A(ram[3529]), .B(ram[3545]), .S(n8776), .Z(n2319) );
  MUX2_X1 U11462 ( .A(n2319), .B(n2318), .S(n4223), .Z(n2320) );
  MUX2_X1 U11463 ( .A(ram[3497]), .B(ram[3513]), .S(n8776), .Z(n2321) );
  MUX2_X1 U11464 ( .A(ram[3465]), .B(ram[3481]), .S(n8776), .Z(n2322) );
  MUX2_X1 U11465 ( .A(n2322), .B(n2321), .S(n4223), .Z(n2323) );
  MUX2_X1 U11466 ( .A(n2323), .B(n2320), .S(n4144), .Z(n2324) );
  MUX2_X1 U11467 ( .A(ram[3433]), .B(ram[3449]), .S(n8777), .Z(n2325) );
  MUX2_X1 U11468 ( .A(ram[3401]), .B(ram[3417]), .S(n8777), .Z(n2326) );
  MUX2_X1 U11469 ( .A(n2326), .B(n2325), .S(n4223), .Z(n2327) );
  MUX2_X1 U11470 ( .A(ram[3369]), .B(ram[3385]), .S(n8777), .Z(n2328) );
  MUX2_X1 U11471 ( .A(ram[3337]), .B(ram[3353]), .S(n8777), .Z(n2329) );
  MUX2_X1 U11472 ( .A(n2329), .B(n2328), .S(n4223), .Z(n2330) );
  MUX2_X1 U11473 ( .A(n2330), .B(n2327), .S(n4144), .Z(n2331) );
  MUX2_X1 U11474 ( .A(n2331), .B(n2324), .S(n4099), .Z(n2332) );
  MUX2_X1 U11475 ( .A(ram[3305]), .B(ram[3321]), .S(n8777), .Z(n2333) );
  MUX2_X1 U11476 ( .A(ram[3273]), .B(ram[3289]), .S(n8777), .Z(n2334) );
  MUX2_X1 U11477 ( .A(n2334), .B(n2333), .S(n4223), .Z(n2335) );
  MUX2_X1 U11478 ( .A(ram[3241]), .B(ram[3257]), .S(n8777), .Z(n2336) );
  MUX2_X1 U11479 ( .A(ram[3209]), .B(ram[3225]), .S(n8777), .Z(n2337) );
  MUX2_X1 U11480 ( .A(n2337), .B(n2336), .S(n4223), .Z(n2338) );
  MUX2_X1 U11481 ( .A(n2338), .B(n2335), .S(n4144), .Z(n2339) );
  MUX2_X1 U11482 ( .A(ram[3177]), .B(ram[3193]), .S(n8777), .Z(n2340) );
  MUX2_X1 U11483 ( .A(ram[3145]), .B(ram[3161]), .S(n8777), .Z(n2341) );
  MUX2_X1 U11484 ( .A(n2341), .B(n2340), .S(n4223), .Z(n2342) );
  MUX2_X1 U11485 ( .A(ram[3113]), .B(ram[3129]), .S(n8777), .Z(n2343) );
  MUX2_X1 U11486 ( .A(ram[3081]), .B(ram[3097]), .S(n8777), .Z(n2344) );
  MUX2_X1 U11487 ( .A(n2344), .B(n2343), .S(n4223), .Z(n2345) );
  MUX2_X1 U11488 ( .A(n2345), .B(n2342), .S(n4144), .Z(n2346) );
  MUX2_X1 U11489 ( .A(n2346), .B(n2339), .S(n4099), .Z(n2347) );
  MUX2_X1 U11490 ( .A(n2347), .B(n2332), .S(n4082), .Z(n2348) );
  MUX2_X1 U11491 ( .A(n2348), .B(n2317), .S(n4071), .Z(n2349) );
  MUX2_X1 U11492 ( .A(ram[3049]), .B(ram[3065]), .S(n8778), .Z(n2350) );
  MUX2_X1 U11493 ( .A(ram[3017]), .B(ram[3033]), .S(n8778), .Z(n2351) );
  MUX2_X1 U11494 ( .A(n2351), .B(n2350), .S(n4224), .Z(n2352) );
  MUX2_X1 U11495 ( .A(ram[2985]), .B(ram[3001]), .S(n8778), .Z(n2353) );
  MUX2_X1 U11496 ( .A(ram[2953]), .B(ram[2969]), .S(n8778), .Z(n2354) );
  MUX2_X1 U11497 ( .A(n2354), .B(n2353), .S(n4224), .Z(n2355) );
  MUX2_X1 U11498 ( .A(n2355), .B(n2352), .S(n4145), .Z(n2356) );
  MUX2_X1 U11499 ( .A(ram[2921]), .B(ram[2937]), .S(n8778), .Z(n2357) );
  MUX2_X1 U11500 ( .A(ram[2889]), .B(ram[2905]), .S(n8778), .Z(n2358) );
  MUX2_X1 U11501 ( .A(n2358), .B(n2357), .S(n4224), .Z(n2359) );
  MUX2_X1 U11502 ( .A(ram[2857]), .B(ram[2873]), .S(n8778), .Z(n2360) );
  MUX2_X1 U11503 ( .A(ram[2825]), .B(ram[2841]), .S(n8778), .Z(n2361) );
  MUX2_X1 U11504 ( .A(n2361), .B(n2360), .S(n4224), .Z(n2362) );
  MUX2_X1 U11505 ( .A(n2362), .B(n2359), .S(n4145), .Z(n2363) );
  MUX2_X1 U11506 ( .A(n2363), .B(n2356), .S(n4100), .Z(n2364) );
  MUX2_X1 U11507 ( .A(ram[2793]), .B(ram[2809]), .S(n8778), .Z(n2365) );
  MUX2_X1 U11508 ( .A(ram[2761]), .B(ram[2777]), .S(n8778), .Z(n2366) );
  MUX2_X1 U11509 ( .A(n2366), .B(n2365), .S(n4224), .Z(n2367) );
  MUX2_X1 U11510 ( .A(ram[2729]), .B(ram[2745]), .S(n8778), .Z(n2368) );
  MUX2_X1 U11511 ( .A(ram[2697]), .B(ram[2713]), .S(n8778), .Z(n2369) );
  MUX2_X1 U11512 ( .A(n2369), .B(n2368), .S(n4224), .Z(n2370) );
  MUX2_X1 U11513 ( .A(n2370), .B(n2367), .S(n4145), .Z(n2371) );
  MUX2_X1 U11514 ( .A(ram[2665]), .B(ram[2681]), .S(n8779), .Z(n2372) );
  MUX2_X1 U11515 ( .A(ram[2633]), .B(ram[2649]), .S(n8779), .Z(n2373) );
  MUX2_X1 U11516 ( .A(n2373), .B(n2372), .S(n4224), .Z(n2374) );
  MUX2_X1 U11517 ( .A(ram[2601]), .B(ram[2617]), .S(n8779), .Z(n2375) );
  MUX2_X1 U11518 ( .A(ram[2569]), .B(ram[2585]), .S(n8779), .Z(n2376) );
  MUX2_X1 U11519 ( .A(n2376), .B(n2375), .S(n4224), .Z(n2377) );
  MUX2_X1 U11520 ( .A(n2377), .B(n2374), .S(n4145), .Z(n2378) );
  MUX2_X1 U11521 ( .A(n2378), .B(n2371), .S(n4100), .Z(n2379) );
  MUX2_X1 U11522 ( .A(n2379), .B(n2364), .S(n4082), .Z(n2380) );
  MUX2_X1 U11523 ( .A(ram[2537]), .B(ram[2553]), .S(n8779), .Z(n2381) );
  MUX2_X1 U11524 ( .A(ram[2505]), .B(ram[2521]), .S(n8779), .Z(n2382) );
  MUX2_X1 U11525 ( .A(n2382), .B(n2381), .S(n4224), .Z(n2383) );
  MUX2_X1 U11526 ( .A(ram[2473]), .B(ram[2489]), .S(n8779), .Z(n2384) );
  MUX2_X1 U11527 ( .A(ram[2441]), .B(ram[2457]), .S(n8779), .Z(n2385) );
  MUX2_X1 U11528 ( .A(n2385), .B(n2384), .S(n4224), .Z(n2386) );
  MUX2_X1 U11529 ( .A(n2386), .B(n2383), .S(n4145), .Z(n2387) );
  MUX2_X1 U11530 ( .A(ram[2409]), .B(ram[2425]), .S(n8779), .Z(n2388) );
  MUX2_X1 U11531 ( .A(ram[2377]), .B(ram[2393]), .S(n8779), .Z(n2389) );
  MUX2_X1 U11532 ( .A(n2389), .B(n2388), .S(n4224), .Z(n2390) );
  MUX2_X1 U11533 ( .A(ram[2345]), .B(ram[2361]), .S(n8779), .Z(n2391) );
  MUX2_X1 U11534 ( .A(ram[2313]), .B(ram[2329]), .S(n8779), .Z(n2392) );
  MUX2_X1 U11535 ( .A(n2392), .B(n2391), .S(n4224), .Z(n2393) );
  MUX2_X1 U11536 ( .A(n2393), .B(n2390), .S(n4145), .Z(n2394) );
  MUX2_X1 U11537 ( .A(n2394), .B(n2387), .S(n4100), .Z(n2395) );
  MUX2_X1 U11538 ( .A(ram[2281]), .B(ram[2297]), .S(n8780), .Z(n2396) );
  MUX2_X1 U11539 ( .A(ram[2249]), .B(ram[2265]), .S(n8780), .Z(n2397) );
  MUX2_X1 U11540 ( .A(n2397), .B(n2396), .S(n4225), .Z(n2398) );
  MUX2_X1 U11541 ( .A(ram[2217]), .B(ram[2233]), .S(n8780), .Z(n2399) );
  MUX2_X1 U11542 ( .A(ram[2185]), .B(ram[2201]), .S(n8780), .Z(n24001) );
  MUX2_X1 U11543 ( .A(n24001), .B(n2399), .S(n4225), .Z(n2401) );
  MUX2_X1 U11544 ( .A(n2401), .B(n2398), .S(n4145), .Z(n2402) );
  MUX2_X1 U11545 ( .A(ram[2153]), .B(ram[2169]), .S(n8780), .Z(n2403) );
  MUX2_X1 U11546 ( .A(ram[2121]), .B(ram[2137]), .S(n8780), .Z(n2404) );
  MUX2_X1 U11547 ( .A(n2404), .B(n2403), .S(n4225), .Z(n2405) );
  MUX2_X1 U11548 ( .A(ram[2089]), .B(ram[2105]), .S(n8780), .Z(n2406) );
  MUX2_X1 U11549 ( .A(ram[2057]), .B(ram[2073]), .S(n8780), .Z(n2407) );
  MUX2_X1 U11550 ( .A(n2407), .B(n2406), .S(n4225), .Z(n2408) );
  MUX2_X1 U11551 ( .A(n2408), .B(n2405), .S(n4145), .Z(n2409) );
  MUX2_X1 U11552 ( .A(n2409), .B(n2402), .S(n4100), .Z(n2410) );
  MUX2_X1 U11553 ( .A(n2410), .B(n2395), .S(n4082), .Z(n2411) );
  MUX2_X1 U11554 ( .A(n2411), .B(n2380), .S(n4071), .Z(n2412) );
  MUX2_X1 U11555 ( .A(n2412), .B(n2349), .S(n4066), .Z(n2413) );
  MUX2_X1 U11556 ( .A(ram[2025]), .B(ram[2041]), .S(n8780), .Z(n2414) );
  MUX2_X1 U11557 ( .A(ram[1993]), .B(ram[2009]), .S(n8780), .Z(n2415) );
  MUX2_X1 U11558 ( .A(n2415), .B(n2414), .S(n4225), .Z(n2416) );
  MUX2_X1 U11559 ( .A(ram[1961]), .B(ram[1977]), .S(n8780), .Z(n2417) );
  MUX2_X1 U11560 ( .A(ram[1929]), .B(ram[1945]), .S(n8780), .Z(n2418) );
  MUX2_X1 U11561 ( .A(n2418), .B(n2417), .S(n4225), .Z(n2419) );
  MUX2_X1 U11562 ( .A(n2419), .B(n2416), .S(n4145), .Z(n2420) );
  MUX2_X1 U11563 ( .A(ram[1897]), .B(ram[1913]), .S(n8781), .Z(n2421) );
  MUX2_X1 U11564 ( .A(ram[1865]), .B(ram[1881]), .S(n8781), .Z(n2422) );
  MUX2_X1 U11565 ( .A(n2422), .B(n2421), .S(n4225), .Z(n2423) );
  MUX2_X1 U11566 ( .A(ram[1833]), .B(ram[1849]), .S(n8781), .Z(n2424) );
  MUX2_X1 U11567 ( .A(ram[1801]), .B(ram[1817]), .S(n8781), .Z(n2425) );
  MUX2_X1 U11568 ( .A(n2425), .B(n2424), .S(n4225), .Z(n2426) );
  MUX2_X1 U11569 ( .A(n2426), .B(n2423), .S(n4145), .Z(n2427) );
  MUX2_X1 U11570 ( .A(n2427), .B(n2420), .S(n4100), .Z(n2428) );
  MUX2_X1 U11571 ( .A(ram[1769]), .B(ram[1785]), .S(n8781), .Z(n2429) );
  MUX2_X1 U11572 ( .A(ram[1737]), .B(ram[1753]), .S(n8781), .Z(n2430) );
  MUX2_X1 U11573 ( .A(n2430), .B(n2429), .S(n4225), .Z(n2431) );
  MUX2_X1 U11574 ( .A(ram[1705]), .B(ram[1721]), .S(n8781), .Z(n2432) );
  MUX2_X1 U11575 ( .A(ram[1673]), .B(ram[1689]), .S(n8781), .Z(n2433) );
  MUX2_X1 U11576 ( .A(n2433), .B(n2432), .S(n4225), .Z(n2434) );
  MUX2_X1 U11577 ( .A(n2434), .B(n2431), .S(n4145), .Z(n2435) );
  MUX2_X1 U11578 ( .A(ram[1641]), .B(ram[1657]), .S(n8781), .Z(n2436) );
  MUX2_X1 U11579 ( .A(ram[1609]), .B(ram[1625]), .S(n8781), .Z(n2437) );
  MUX2_X1 U11580 ( .A(n2437), .B(n2436), .S(n4225), .Z(n2438) );
  MUX2_X1 U11581 ( .A(ram[1577]), .B(ram[1593]), .S(n8781), .Z(n2439) );
  MUX2_X1 U11582 ( .A(ram[1545]), .B(ram[1561]), .S(n8781), .Z(n2440) );
  MUX2_X1 U11583 ( .A(n2440), .B(n2439), .S(n4225), .Z(n2441) );
  MUX2_X1 U11584 ( .A(n2441), .B(n2438), .S(n4145), .Z(n2442) );
  MUX2_X1 U11585 ( .A(n2442), .B(n2435), .S(n4100), .Z(n2443) );
  MUX2_X1 U11586 ( .A(n2443), .B(n2428), .S(n4082), .Z(n2444) );
  MUX2_X1 U11587 ( .A(ram[1513]), .B(ram[1529]), .S(n8782), .Z(n2445) );
  MUX2_X1 U11588 ( .A(ram[1481]), .B(ram[1497]), .S(n8782), .Z(n2446) );
  MUX2_X1 U11589 ( .A(n2446), .B(n2445), .S(n4226), .Z(n2447) );
  MUX2_X1 U11590 ( .A(ram[1449]), .B(ram[1465]), .S(n8782), .Z(n2448) );
  MUX2_X1 U11591 ( .A(ram[1417]), .B(ram[1433]), .S(n8782), .Z(n2449) );
  MUX2_X1 U11592 ( .A(n2449), .B(n2448), .S(n4226), .Z(n2450) );
  MUX2_X1 U11593 ( .A(n2450), .B(n2447), .S(n4146), .Z(n2451) );
  MUX2_X1 U11594 ( .A(ram[1385]), .B(ram[1401]), .S(n8782), .Z(n2452) );
  MUX2_X1 U11595 ( .A(ram[1353]), .B(ram[1369]), .S(n8782), .Z(n2453) );
  MUX2_X1 U11596 ( .A(n2453), .B(n2452), .S(n4226), .Z(n2454) );
  MUX2_X1 U11597 ( .A(ram[1321]), .B(ram[1337]), .S(n8782), .Z(n2455) );
  MUX2_X1 U11598 ( .A(ram[1289]), .B(ram[1305]), .S(n8782), .Z(n2456) );
  MUX2_X1 U11599 ( .A(n2456), .B(n2455), .S(n4226), .Z(n2457) );
  MUX2_X1 U11600 ( .A(n2457), .B(n2454), .S(n4146), .Z(n2458) );
  MUX2_X1 U11601 ( .A(n2458), .B(n2451), .S(n4100), .Z(n2459) );
  MUX2_X1 U11602 ( .A(ram[1257]), .B(ram[1273]), .S(n8782), .Z(n2460) );
  MUX2_X1 U11603 ( .A(ram[1225]), .B(ram[1241]), .S(n8782), .Z(n2461) );
  MUX2_X1 U11604 ( .A(n2461), .B(n2460), .S(n4226), .Z(n2462) );
  MUX2_X1 U11605 ( .A(ram[1193]), .B(ram[1209]), .S(n8782), .Z(n2463) );
  MUX2_X1 U11606 ( .A(ram[1161]), .B(ram[1177]), .S(n8782), .Z(n2464) );
  MUX2_X1 U11607 ( .A(n2464), .B(n2463), .S(n4226), .Z(n2465) );
  MUX2_X1 U11608 ( .A(n2465), .B(n2462), .S(n4146), .Z(n2466) );
  MUX2_X1 U11609 ( .A(ram[1129]), .B(ram[1145]), .S(n8783), .Z(n2467) );
  MUX2_X1 U11610 ( .A(ram[1097]), .B(ram[1113]), .S(n8783), .Z(n2468) );
  MUX2_X1 U11611 ( .A(n2468), .B(n2467), .S(n4226), .Z(n2469) );
  MUX2_X1 U11612 ( .A(ram[1065]), .B(ram[1081]), .S(n8783), .Z(n2470) );
  MUX2_X1 U11613 ( .A(ram[1033]), .B(ram[1049]), .S(n8783), .Z(n2471) );
  MUX2_X1 U11614 ( .A(n2471), .B(n2470), .S(n4226), .Z(n2472) );
  MUX2_X1 U11615 ( .A(n2472), .B(n2469), .S(n4146), .Z(n2473) );
  MUX2_X1 U11616 ( .A(n2473), .B(n2466), .S(n4100), .Z(n2474) );
  MUX2_X1 U11617 ( .A(n2474), .B(n2459), .S(n4082), .Z(n2475) );
  MUX2_X1 U11618 ( .A(n2475), .B(n2444), .S(n4071), .Z(n2476) );
  MUX2_X1 U11619 ( .A(ram[1001]), .B(ram[1017]), .S(n8783), .Z(n2477) );
  MUX2_X1 U11620 ( .A(ram[969]), .B(ram[985]), .S(n8783), .Z(n2478) );
  MUX2_X1 U11621 ( .A(n2478), .B(n2477), .S(n4226), .Z(n2479) );
  MUX2_X1 U11622 ( .A(ram[937]), .B(ram[953]), .S(n8783), .Z(n2480) );
  MUX2_X1 U11623 ( .A(ram[905]), .B(ram[921]), .S(n8783), .Z(n2481) );
  MUX2_X1 U11624 ( .A(n2481), .B(n2480), .S(n4226), .Z(n2482) );
  MUX2_X1 U11625 ( .A(n2482), .B(n2479), .S(n4146), .Z(n2483) );
  MUX2_X1 U11626 ( .A(ram[873]), .B(ram[889]), .S(n8783), .Z(n2484) );
  MUX2_X1 U11627 ( .A(ram[841]), .B(ram[857]), .S(n8783), .Z(n2485) );
  MUX2_X1 U11628 ( .A(n2485), .B(n2484), .S(n4226), .Z(n2486) );
  MUX2_X1 U11629 ( .A(ram[809]), .B(ram[825]), .S(n8783), .Z(n2487) );
  MUX2_X1 U11630 ( .A(ram[777]), .B(ram[793]), .S(n8783), .Z(n2488) );
  MUX2_X1 U11631 ( .A(n2488), .B(n2487), .S(n4226), .Z(n2489) );
  MUX2_X1 U11632 ( .A(n2489), .B(n2486), .S(n4146), .Z(n2490) );
  MUX2_X1 U11633 ( .A(n2490), .B(n2483), .S(n4100), .Z(n2491) );
  MUX2_X1 U11634 ( .A(ram[745]), .B(ram[761]), .S(n8784), .Z(n2492) );
  MUX2_X1 U11635 ( .A(ram[713]), .B(ram[729]), .S(n8784), .Z(n2493) );
  MUX2_X1 U11636 ( .A(n2493), .B(n2492), .S(n4227), .Z(n2494) );
  MUX2_X1 U11637 ( .A(ram[681]), .B(ram[697]), .S(n8784), .Z(n2495) );
  MUX2_X1 U11638 ( .A(ram[649]), .B(ram[665]), .S(n8784), .Z(n2496) );
  MUX2_X1 U11639 ( .A(n2496), .B(n2495), .S(n4227), .Z(n2497) );
  MUX2_X1 U11640 ( .A(n2497), .B(n2494), .S(n4146), .Z(n2498) );
  MUX2_X1 U11641 ( .A(ram[617]), .B(ram[633]), .S(n8784), .Z(n2499) );
  MUX2_X1 U11642 ( .A(ram[585]), .B(ram[601]), .S(n8784), .Z(n25001) );
  MUX2_X1 U11643 ( .A(n25001), .B(n2499), .S(n4227), .Z(n2501) );
  MUX2_X1 U11644 ( .A(ram[553]), .B(ram[569]), .S(n8784), .Z(n2502) );
  MUX2_X1 U11645 ( .A(ram[521]), .B(ram[537]), .S(n8784), .Z(n2503) );
  MUX2_X1 U11646 ( .A(n2503), .B(n2502), .S(n4227), .Z(n2504) );
  MUX2_X1 U11647 ( .A(n2504), .B(n2501), .S(n4146), .Z(n2505) );
  MUX2_X1 U11648 ( .A(n2505), .B(n2498), .S(n4100), .Z(n2506) );
  MUX2_X1 U11649 ( .A(n2506), .B(n2491), .S(n4082), .Z(n2507) );
  MUX2_X1 U11650 ( .A(ram[489]), .B(ram[505]), .S(n8784), .Z(n2508) );
  MUX2_X1 U11651 ( .A(ram[457]), .B(ram[473]), .S(n8784), .Z(n2509) );
  MUX2_X1 U11652 ( .A(n2509), .B(n2508), .S(n4227), .Z(n2510) );
  MUX2_X1 U11653 ( .A(ram[425]), .B(ram[441]), .S(n8784), .Z(n2511) );
  MUX2_X1 U11654 ( .A(ram[393]), .B(ram[409]), .S(n8784), .Z(n2512) );
  MUX2_X1 U11655 ( .A(n2512), .B(n2511), .S(n4227), .Z(n2513) );
  MUX2_X1 U11656 ( .A(n2513), .B(n2510), .S(n4146), .Z(n2514) );
  MUX2_X1 U11657 ( .A(ram[361]), .B(ram[377]), .S(n8785), .Z(n2515) );
  MUX2_X1 U11658 ( .A(ram[329]), .B(ram[345]), .S(n8785), .Z(n2516) );
  MUX2_X1 U11659 ( .A(n2516), .B(n2515), .S(n4227), .Z(n2517) );
  MUX2_X1 U11660 ( .A(ram[297]), .B(ram[313]), .S(n8785), .Z(n2518) );
  MUX2_X1 U11661 ( .A(ram[265]), .B(ram[281]), .S(n8785), .Z(n2519) );
  MUX2_X1 U11662 ( .A(n2519), .B(n2518), .S(n4227), .Z(n2520) );
  MUX2_X1 U11663 ( .A(n2520), .B(n2517), .S(n4146), .Z(n2521) );
  MUX2_X1 U11664 ( .A(n2521), .B(n2514), .S(n4100), .Z(n2522) );
  MUX2_X1 U11665 ( .A(ram[233]), .B(ram[249]), .S(n8785), .Z(n2523) );
  MUX2_X1 U11666 ( .A(ram[201]), .B(ram[217]), .S(n8785), .Z(n2524) );
  MUX2_X1 U11667 ( .A(n2524), .B(n2523), .S(n4227), .Z(n2525) );
  MUX2_X1 U11668 ( .A(ram[169]), .B(ram[185]), .S(n8785), .Z(n2526) );
  MUX2_X1 U11669 ( .A(ram[137]), .B(ram[153]), .S(n8785), .Z(n2527) );
  MUX2_X1 U11670 ( .A(n2527), .B(n2526), .S(n4227), .Z(n2528) );
  MUX2_X1 U11671 ( .A(n2528), .B(n2525), .S(n4146), .Z(n2529) );
  MUX2_X1 U11672 ( .A(ram[105]), .B(ram[121]), .S(n8785), .Z(n2530) );
  MUX2_X1 U11673 ( .A(ram[73]), .B(ram[89]), .S(n8785), .Z(n2531) );
  MUX2_X1 U11674 ( .A(n2531), .B(n2530), .S(n4227), .Z(n2532) );
  MUX2_X1 U11675 ( .A(ram[41]), .B(ram[57]), .S(n8785), .Z(n2533) );
  MUX2_X1 U11676 ( .A(ram[9]), .B(ram[25]), .S(n8785), .Z(n2534) );
  MUX2_X1 U11677 ( .A(n2534), .B(n2533), .S(n4227), .Z(n2535) );
  MUX2_X1 U11678 ( .A(n2535), .B(n2532), .S(n4146), .Z(n2536) );
  MUX2_X1 U11679 ( .A(n2536), .B(n2529), .S(n4100), .Z(n2537) );
  MUX2_X1 U11680 ( .A(n2537), .B(n2522), .S(n4082), .Z(n2538) );
  MUX2_X1 U11681 ( .A(n2538), .B(n2507), .S(n4071), .Z(n2539) );
  MUX2_X1 U11682 ( .A(n2539), .B(n2476), .S(n4066), .Z(n2540) );
  MUX2_X1 U11683 ( .A(n2540), .B(n2413), .S(mem_access_addr[9]), .Z(N292) );
  MUX2_X1 U11684 ( .A(ram[4074]), .B(ram[4090]), .S(n8786), .Z(n2541) );
  MUX2_X1 U11685 ( .A(ram[4042]), .B(ram[4058]), .S(n8786), .Z(n2542) );
  MUX2_X1 U11686 ( .A(n2542), .B(n2541), .S(n4228), .Z(n2543) );
  MUX2_X1 U11687 ( .A(ram[4010]), .B(ram[4026]), .S(n8786), .Z(n2544) );
  MUX2_X1 U11688 ( .A(ram[3978]), .B(ram[3994]), .S(n8786), .Z(n2545) );
  MUX2_X1 U11689 ( .A(n2545), .B(n2544), .S(n4228), .Z(n2546) );
  MUX2_X1 U11690 ( .A(n2546), .B(n2543), .S(n4147), .Z(n2547) );
  MUX2_X1 U11691 ( .A(ram[3946]), .B(ram[3962]), .S(n8786), .Z(n2548) );
  MUX2_X1 U11692 ( .A(ram[3914]), .B(ram[3930]), .S(n8786), .Z(n2549) );
  MUX2_X1 U11693 ( .A(n2549), .B(n2548), .S(n4228), .Z(n2550) );
  MUX2_X1 U11694 ( .A(ram[3882]), .B(ram[3898]), .S(n8786), .Z(n2551) );
  MUX2_X1 U11695 ( .A(ram[3850]), .B(ram[3866]), .S(n8786), .Z(n2552) );
  MUX2_X1 U11696 ( .A(n2552), .B(n2551), .S(n4228), .Z(n2553) );
  MUX2_X1 U11697 ( .A(n2553), .B(n2550), .S(n4147), .Z(n2554) );
  MUX2_X1 U11698 ( .A(n2554), .B(n2547), .S(n4101), .Z(n2555) );
  MUX2_X1 U11699 ( .A(ram[3818]), .B(ram[3834]), .S(n8786), .Z(n2556) );
  MUX2_X1 U11700 ( .A(ram[3786]), .B(ram[3802]), .S(n8786), .Z(n2557) );
  MUX2_X1 U11701 ( .A(n2557), .B(n2556), .S(n4228), .Z(n2558) );
  MUX2_X1 U11702 ( .A(ram[3754]), .B(ram[3770]), .S(n8786), .Z(n2559) );
  MUX2_X1 U11703 ( .A(ram[3722]), .B(ram[3738]), .S(n8786), .Z(n2560) );
  MUX2_X1 U11704 ( .A(n2560), .B(n2559), .S(n4228), .Z(n2561) );
  MUX2_X1 U11705 ( .A(n2561), .B(n2558), .S(n4147), .Z(n2562) );
  MUX2_X1 U11706 ( .A(ram[3690]), .B(ram[3706]), .S(n8787), .Z(n2563) );
  MUX2_X1 U11707 ( .A(ram[3658]), .B(ram[3674]), .S(n8787), .Z(n2564) );
  MUX2_X1 U11708 ( .A(n2564), .B(n2563), .S(n4228), .Z(n2565) );
  MUX2_X1 U11709 ( .A(ram[3626]), .B(ram[3642]), .S(n8787), .Z(n2566) );
  MUX2_X1 U11710 ( .A(ram[3594]), .B(ram[3610]), .S(n8787), .Z(n2567) );
  MUX2_X1 U11711 ( .A(n2567), .B(n2566), .S(n4228), .Z(n2568) );
  MUX2_X1 U11712 ( .A(n2568), .B(n2565), .S(n4147), .Z(n2569) );
  MUX2_X1 U11713 ( .A(n2569), .B(n2562), .S(n4101), .Z(n2570) );
  MUX2_X1 U11714 ( .A(n2570), .B(n2555), .S(n4083), .Z(n2571) );
  MUX2_X1 U11715 ( .A(ram[3562]), .B(ram[3578]), .S(n8787), .Z(n2572) );
  MUX2_X1 U11716 ( .A(ram[3530]), .B(ram[3546]), .S(n8787), .Z(n2573) );
  MUX2_X1 U11717 ( .A(n2573), .B(n2572), .S(n4228), .Z(n2574) );
  MUX2_X1 U11718 ( .A(ram[3498]), .B(ram[3514]), .S(n8787), .Z(n2575) );
  MUX2_X1 U11719 ( .A(ram[3466]), .B(ram[3482]), .S(n8787), .Z(n2576) );
  MUX2_X1 U11720 ( .A(n2576), .B(n2575), .S(n4228), .Z(n2577) );
  MUX2_X1 U11721 ( .A(n2577), .B(n2574), .S(n4147), .Z(n2578) );
  MUX2_X1 U11722 ( .A(ram[3434]), .B(ram[3450]), .S(n8787), .Z(n2579) );
  MUX2_X1 U11723 ( .A(ram[3402]), .B(ram[3418]), .S(n8787), .Z(n2580) );
  MUX2_X1 U11724 ( .A(n2580), .B(n2579), .S(n4228), .Z(n2581) );
  MUX2_X1 U11725 ( .A(ram[3370]), .B(ram[3386]), .S(n8787), .Z(n2582) );
  MUX2_X1 U11726 ( .A(ram[3338]), .B(ram[3354]), .S(n8787), .Z(n2583) );
  MUX2_X1 U11727 ( .A(n2583), .B(n2582), .S(n4228), .Z(n2584) );
  MUX2_X1 U11728 ( .A(n2584), .B(n2581), .S(n4147), .Z(n2585) );
  MUX2_X1 U11729 ( .A(n2585), .B(n2578), .S(n4101), .Z(n2586) );
  MUX2_X1 U11730 ( .A(ram[3306]), .B(ram[3322]), .S(n8788), .Z(n2587) );
  MUX2_X1 U11731 ( .A(ram[3274]), .B(ram[3290]), .S(n8788), .Z(n2588) );
  MUX2_X1 U11732 ( .A(n2588), .B(n2587), .S(n4229), .Z(n2589) );
  MUX2_X1 U11733 ( .A(ram[3242]), .B(ram[3258]), .S(n8788), .Z(n2590) );
  MUX2_X1 U11734 ( .A(ram[3210]), .B(ram[3226]), .S(n8788), .Z(n2591) );
  MUX2_X1 U11735 ( .A(n2591), .B(n2590), .S(n4229), .Z(n2592) );
  MUX2_X1 U11736 ( .A(n2592), .B(n2589), .S(n4147), .Z(n2593) );
  MUX2_X1 U11737 ( .A(ram[3178]), .B(ram[3194]), .S(n8788), .Z(n2594) );
  MUX2_X1 U11738 ( .A(ram[3146]), .B(ram[3162]), .S(n8788), .Z(n2595) );
  MUX2_X1 U11739 ( .A(n2595), .B(n2594), .S(n4229), .Z(n2596) );
  MUX2_X1 U11740 ( .A(ram[3114]), .B(ram[3130]), .S(n8788), .Z(n2597) );
  MUX2_X1 U11741 ( .A(ram[3082]), .B(ram[3098]), .S(n8788), .Z(n2598) );
  MUX2_X1 U11742 ( .A(n2598), .B(n2597), .S(n4229), .Z(n2599) );
  MUX2_X1 U11743 ( .A(n2599), .B(n2596), .S(n4147), .Z(n26001) );
  MUX2_X1 U11744 ( .A(n26001), .B(n2593), .S(n4101), .Z(n2601) );
  MUX2_X1 U11745 ( .A(n2601), .B(n2586), .S(n4083), .Z(n2602) );
  MUX2_X1 U11746 ( .A(n2602), .B(n2571), .S(n4072), .Z(n2603) );
  MUX2_X1 U11747 ( .A(ram[3050]), .B(ram[3066]), .S(n8788), .Z(n2604) );
  MUX2_X1 U11748 ( .A(ram[3018]), .B(ram[3034]), .S(n8788), .Z(n2605) );
  MUX2_X1 U11749 ( .A(n2605), .B(n2604), .S(n4229), .Z(n2606) );
  MUX2_X1 U11750 ( .A(ram[2986]), .B(ram[3002]), .S(n8788), .Z(n2607) );
  MUX2_X1 U11751 ( .A(ram[2954]), .B(ram[2970]), .S(n8788), .Z(n2608) );
  MUX2_X1 U11752 ( .A(n2608), .B(n2607), .S(n4229), .Z(n2609) );
  MUX2_X1 U11753 ( .A(n2609), .B(n2606), .S(n4147), .Z(n2610) );
  MUX2_X1 U11754 ( .A(ram[2922]), .B(ram[2938]), .S(n8789), .Z(n2611) );
  MUX2_X1 U11755 ( .A(ram[2890]), .B(ram[2906]), .S(n8789), .Z(n2612) );
  MUX2_X1 U11756 ( .A(n2612), .B(n2611), .S(n4229), .Z(n2613) );
  MUX2_X1 U11757 ( .A(ram[2858]), .B(ram[2874]), .S(n8789), .Z(n2614) );
  MUX2_X1 U11758 ( .A(ram[2826]), .B(ram[2842]), .S(n8789), .Z(n2615) );
  MUX2_X1 U11759 ( .A(n2615), .B(n2614), .S(n4229), .Z(n2616) );
  MUX2_X1 U11760 ( .A(n2616), .B(n2613), .S(n4147), .Z(n2617) );
  MUX2_X1 U11761 ( .A(n2617), .B(n2610), .S(n4101), .Z(n2618) );
  MUX2_X1 U11762 ( .A(ram[2794]), .B(ram[2810]), .S(n8789), .Z(n2619) );
  MUX2_X1 U11763 ( .A(ram[2762]), .B(ram[2778]), .S(n8789), .Z(n2620) );
  MUX2_X1 U11764 ( .A(n2620), .B(n2619), .S(n4229), .Z(n2621) );
  MUX2_X1 U11765 ( .A(ram[2730]), .B(ram[2746]), .S(n8789), .Z(n2622) );
  MUX2_X1 U11766 ( .A(ram[2698]), .B(ram[2714]), .S(n8789), .Z(n2623) );
  MUX2_X1 U11767 ( .A(n2623), .B(n2622), .S(n4229), .Z(n2624) );
  MUX2_X1 U11768 ( .A(n2624), .B(n2621), .S(n4147), .Z(n2625) );
  MUX2_X1 U11769 ( .A(ram[2666]), .B(ram[2682]), .S(n8789), .Z(n2626) );
  MUX2_X1 U11770 ( .A(ram[2634]), .B(ram[2650]), .S(n8789), .Z(n2627) );
  MUX2_X1 U11771 ( .A(n2627), .B(n2626), .S(n4229), .Z(n2628) );
  MUX2_X1 U11772 ( .A(ram[2602]), .B(ram[2618]), .S(n8789), .Z(n2629) );
  MUX2_X1 U11773 ( .A(ram[2570]), .B(ram[2586]), .S(n8789), .Z(n2630) );
  MUX2_X1 U11774 ( .A(n2630), .B(n2629), .S(n4229), .Z(n2631) );
  MUX2_X1 U11775 ( .A(n2631), .B(n2628), .S(n4147), .Z(n2632) );
  MUX2_X1 U11776 ( .A(n2632), .B(n2625), .S(n4101), .Z(n2633) );
  MUX2_X1 U11777 ( .A(n2633), .B(n2618), .S(n4083), .Z(n2634) );
  MUX2_X1 U11778 ( .A(ram[2538]), .B(ram[2554]), .S(n8790), .Z(n2635) );
  MUX2_X1 U11779 ( .A(ram[2506]), .B(ram[2522]), .S(n8790), .Z(n2636) );
  MUX2_X1 U11780 ( .A(n2636), .B(n2635), .S(n4230), .Z(n2637) );
  MUX2_X1 U11781 ( .A(ram[2474]), .B(ram[2490]), .S(n8790), .Z(n2638) );
  MUX2_X1 U11782 ( .A(ram[2442]), .B(ram[2458]), .S(n8790), .Z(n2639) );
  MUX2_X1 U11783 ( .A(n2639), .B(n2638), .S(n4230), .Z(n2640) );
  MUX2_X1 U11784 ( .A(n2640), .B(n2637), .S(n4148), .Z(n2641) );
  MUX2_X1 U11785 ( .A(ram[2410]), .B(ram[2426]), .S(n8790), .Z(n2642) );
  MUX2_X1 U11786 ( .A(ram[2378]), .B(ram[2394]), .S(n8790), .Z(n2643) );
  MUX2_X1 U11787 ( .A(n2643), .B(n2642), .S(n4230), .Z(n2644) );
  MUX2_X1 U11788 ( .A(ram[2346]), .B(ram[2362]), .S(n8790), .Z(n2645) );
  MUX2_X1 U11789 ( .A(ram[2314]), .B(ram[2330]), .S(n8790), .Z(n2646) );
  MUX2_X1 U11790 ( .A(n2646), .B(n2645), .S(n4230), .Z(n2647) );
  MUX2_X1 U11791 ( .A(n2647), .B(n2644), .S(n4148), .Z(n2648) );
  MUX2_X1 U11792 ( .A(n2648), .B(n2641), .S(n4101), .Z(n2649) );
  MUX2_X1 U11793 ( .A(ram[2282]), .B(ram[2298]), .S(n8790), .Z(n2650) );
  MUX2_X1 U11794 ( .A(ram[2250]), .B(ram[2266]), .S(n8790), .Z(n2651) );
  MUX2_X1 U11795 ( .A(n2651), .B(n2650), .S(n4230), .Z(n2652) );
  MUX2_X1 U11796 ( .A(ram[2218]), .B(ram[2234]), .S(n8790), .Z(n2653) );
  MUX2_X1 U11797 ( .A(ram[2186]), .B(ram[2202]), .S(n8790), .Z(n2654) );
  MUX2_X1 U11798 ( .A(n2654), .B(n2653), .S(n4230), .Z(n2655) );
  MUX2_X1 U11799 ( .A(n2655), .B(n2652), .S(n4148), .Z(n2656) );
  MUX2_X1 U11800 ( .A(ram[2154]), .B(ram[2170]), .S(n8791), .Z(n2657) );
  MUX2_X1 U11801 ( .A(ram[2122]), .B(ram[2138]), .S(n8791), .Z(n2658) );
  MUX2_X1 U11802 ( .A(n2658), .B(n2657), .S(n4230), .Z(n2659) );
  MUX2_X1 U11803 ( .A(ram[2090]), .B(ram[2106]), .S(n8791), .Z(n2660) );
  MUX2_X1 U11804 ( .A(ram[2058]), .B(ram[2074]), .S(n8791), .Z(n2661) );
  MUX2_X1 U11805 ( .A(n2661), .B(n2660), .S(n4230), .Z(n2662) );
  MUX2_X1 U11806 ( .A(n2662), .B(n2659), .S(n4148), .Z(n2663) );
  MUX2_X1 U11807 ( .A(n2663), .B(n2656), .S(n4101), .Z(n2664) );
  MUX2_X1 U11808 ( .A(n2664), .B(n2649), .S(n4083), .Z(n2665) );
  MUX2_X1 U11809 ( .A(n2665), .B(n2634), .S(n4072), .Z(n2666) );
  MUX2_X1 U11810 ( .A(n2666), .B(n2603), .S(n4067), .Z(n2667) );
  MUX2_X1 U11811 ( .A(ram[2026]), .B(ram[2042]), .S(n8791), .Z(n2668) );
  MUX2_X1 U11812 ( .A(ram[1994]), .B(ram[2010]), .S(n8791), .Z(n2669) );
  MUX2_X1 U11813 ( .A(n2669), .B(n2668), .S(n4230), .Z(n2670) );
  MUX2_X1 U11814 ( .A(ram[1962]), .B(ram[1978]), .S(n8791), .Z(n2671) );
  MUX2_X1 U11815 ( .A(ram[1930]), .B(ram[1946]), .S(n8791), .Z(n2672) );
  MUX2_X1 U11816 ( .A(n2672), .B(n2671), .S(n4230), .Z(n2673) );
  MUX2_X1 U11817 ( .A(n2673), .B(n2670), .S(n4148), .Z(n2674) );
  MUX2_X1 U11818 ( .A(ram[1898]), .B(ram[1914]), .S(n8791), .Z(n2675) );
  MUX2_X1 U11819 ( .A(ram[1866]), .B(ram[1882]), .S(n8791), .Z(n2676) );
  MUX2_X1 U11820 ( .A(n2676), .B(n2675), .S(n4230), .Z(n2677) );
  MUX2_X1 U11821 ( .A(ram[1834]), .B(ram[1850]), .S(n8791), .Z(n2678) );
  MUX2_X1 U11822 ( .A(ram[1802]), .B(ram[1818]), .S(n8791), .Z(n2679) );
  MUX2_X1 U11823 ( .A(n2679), .B(n2678), .S(n4230), .Z(n2680) );
  MUX2_X1 U11824 ( .A(n2680), .B(n2677), .S(n4148), .Z(n2681) );
  MUX2_X1 U11825 ( .A(n2681), .B(n2674), .S(n4101), .Z(n2682) );
  MUX2_X1 U11826 ( .A(ram[1770]), .B(ram[1786]), .S(n8792), .Z(n2683) );
  MUX2_X1 U11827 ( .A(ram[1738]), .B(ram[1754]), .S(n8792), .Z(n2684) );
  MUX2_X1 U11828 ( .A(n2684), .B(n2683), .S(n4231), .Z(n2685) );
  MUX2_X1 U11829 ( .A(ram[1706]), .B(ram[1722]), .S(n8792), .Z(n2686) );
  MUX2_X1 U11830 ( .A(ram[1674]), .B(ram[1690]), .S(n8792), .Z(n2687) );
  MUX2_X1 U11831 ( .A(n2687), .B(n2686), .S(n4231), .Z(n2688) );
  MUX2_X1 U11832 ( .A(n2688), .B(n2685), .S(n4148), .Z(n2689) );
  MUX2_X1 U11833 ( .A(ram[1642]), .B(ram[1658]), .S(n8792), .Z(n2690) );
  MUX2_X1 U11834 ( .A(ram[1610]), .B(ram[1626]), .S(n8792), .Z(n2691) );
  MUX2_X1 U11835 ( .A(n2691), .B(n2690), .S(n4231), .Z(n2692) );
  MUX2_X1 U11836 ( .A(ram[1578]), .B(ram[1594]), .S(n8792), .Z(n2693) );
  MUX2_X1 U11837 ( .A(ram[1546]), .B(ram[1562]), .S(n8792), .Z(n2694) );
  MUX2_X1 U11838 ( .A(n2694), .B(n2693), .S(n4231), .Z(n2695) );
  MUX2_X1 U11839 ( .A(n2695), .B(n2692), .S(n4148), .Z(n2696) );
  MUX2_X1 U11840 ( .A(n2696), .B(n2689), .S(n4101), .Z(n2697) );
  MUX2_X1 U11841 ( .A(n2697), .B(n2682), .S(n4083), .Z(n2698) );
  MUX2_X1 U11842 ( .A(ram[1514]), .B(ram[1530]), .S(n8792), .Z(n2699) );
  MUX2_X1 U11843 ( .A(ram[1482]), .B(ram[1498]), .S(n8792), .Z(n27001) );
  MUX2_X1 U11844 ( .A(n27001), .B(n2699), .S(n4231), .Z(n2701) );
  MUX2_X1 U11845 ( .A(ram[1450]), .B(ram[1466]), .S(n8792), .Z(n2702) );
  MUX2_X1 U11846 ( .A(ram[1418]), .B(ram[1434]), .S(n8792), .Z(n2703) );
  MUX2_X1 U11847 ( .A(n2703), .B(n2702), .S(n4231), .Z(n2704) );
  MUX2_X1 U11848 ( .A(n2704), .B(n2701), .S(n4148), .Z(n2705) );
  MUX2_X1 U11849 ( .A(ram[1386]), .B(ram[1402]), .S(n8793), .Z(n2706) );
  MUX2_X1 U11850 ( .A(ram[1354]), .B(ram[1370]), .S(n8793), .Z(n2707) );
  MUX2_X1 U11851 ( .A(n2707), .B(n2706), .S(n4231), .Z(n2708) );
  MUX2_X1 U11852 ( .A(ram[1322]), .B(ram[1338]), .S(n8793), .Z(n2709) );
  MUX2_X1 U11853 ( .A(ram[1290]), .B(ram[1306]), .S(n8793), .Z(n2710) );
  MUX2_X1 U11854 ( .A(n2710), .B(n2709), .S(n4231), .Z(n2711) );
  MUX2_X1 U11855 ( .A(n2711), .B(n2708), .S(n4148), .Z(n2712) );
  MUX2_X1 U11856 ( .A(n2712), .B(n2705), .S(n4101), .Z(n2713) );
  MUX2_X1 U11857 ( .A(ram[1258]), .B(ram[1274]), .S(n8793), .Z(n2714) );
  MUX2_X1 U11858 ( .A(ram[1226]), .B(ram[1242]), .S(n8793), .Z(n2715) );
  MUX2_X1 U11859 ( .A(n2715), .B(n2714), .S(n4231), .Z(n2716) );
  MUX2_X1 U11860 ( .A(ram[1194]), .B(ram[1210]), .S(n8793), .Z(n2717) );
  MUX2_X1 U11861 ( .A(ram[1162]), .B(ram[1178]), .S(n8793), .Z(n2718) );
  MUX2_X1 U11862 ( .A(n2718), .B(n2717), .S(n4231), .Z(n2719) );
  MUX2_X1 U11863 ( .A(n2719), .B(n2716), .S(n4148), .Z(n2720) );
  MUX2_X1 U11864 ( .A(ram[1130]), .B(ram[1146]), .S(n8793), .Z(n2721) );
  MUX2_X1 U11865 ( .A(ram[1098]), .B(ram[1114]), .S(n8793), .Z(n2722) );
  MUX2_X1 U11866 ( .A(n2722), .B(n2721), .S(n4231), .Z(n2723) );
  MUX2_X1 U11867 ( .A(ram[1066]), .B(ram[1082]), .S(n8793), .Z(n2724) );
  MUX2_X1 U11868 ( .A(ram[1034]), .B(ram[1050]), .S(n8793), .Z(n2725) );
  MUX2_X1 U11869 ( .A(n2725), .B(n2724), .S(n4231), .Z(n2726) );
  MUX2_X1 U11870 ( .A(n2726), .B(n2723), .S(n4148), .Z(n2727) );
  MUX2_X1 U11871 ( .A(n2727), .B(n2720), .S(n4101), .Z(n2728) );
  MUX2_X1 U11872 ( .A(n2728), .B(n2713), .S(n4083), .Z(n2729) );
  MUX2_X1 U11873 ( .A(n2729), .B(n2698), .S(n4072), .Z(n2730) );
  MUX2_X1 U11874 ( .A(ram[1002]), .B(ram[1018]), .S(n8794), .Z(n2731) );
  MUX2_X1 U11875 ( .A(ram[970]), .B(ram[986]), .S(n8794), .Z(n2732) );
  MUX2_X1 U11876 ( .A(n2732), .B(n2731), .S(n4232), .Z(n2733) );
  MUX2_X1 U11877 ( .A(ram[938]), .B(ram[954]), .S(n8794), .Z(n2734) );
  MUX2_X1 U11878 ( .A(ram[906]), .B(ram[922]), .S(n8794), .Z(n2735) );
  MUX2_X1 U11879 ( .A(n2735), .B(n2734), .S(n4232), .Z(n2736) );
  MUX2_X1 U11880 ( .A(n2736), .B(n2733), .S(n4149), .Z(n2737) );
  MUX2_X1 U11881 ( .A(ram[874]), .B(ram[890]), .S(n8794), .Z(n2738) );
  MUX2_X1 U11882 ( .A(ram[842]), .B(ram[858]), .S(n8794), .Z(n2739) );
  MUX2_X1 U11883 ( .A(n2739), .B(n2738), .S(n4232), .Z(n2740) );
  MUX2_X1 U11884 ( .A(ram[810]), .B(ram[826]), .S(n8794), .Z(n2741) );
  MUX2_X1 U11885 ( .A(ram[778]), .B(ram[794]), .S(n8794), .Z(n2742) );
  MUX2_X1 U11886 ( .A(n2742), .B(n2741), .S(n4232), .Z(n2743) );
  MUX2_X1 U11887 ( .A(n2743), .B(n2740), .S(n4149), .Z(n2744) );
  MUX2_X1 U11888 ( .A(n2744), .B(n2737), .S(n4102), .Z(n2745) );
  MUX2_X1 U11889 ( .A(ram[746]), .B(ram[762]), .S(n8794), .Z(n2746) );
  MUX2_X1 U11890 ( .A(ram[714]), .B(ram[730]), .S(n8794), .Z(n2747) );
  MUX2_X1 U11891 ( .A(n2747), .B(n2746), .S(n4232), .Z(n2748) );
  MUX2_X1 U11892 ( .A(ram[682]), .B(ram[698]), .S(n8794), .Z(n2749) );
  MUX2_X1 U11893 ( .A(ram[650]), .B(ram[666]), .S(n8794), .Z(n2750) );
  MUX2_X1 U11894 ( .A(n2750), .B(n2749), .S(n4232), .Z(n2751) );
  MUX2_X1 U11895 ( .A(n2751), .B(n2748), .S(n4149), .Z(n2752) );
  MUX2_X1 U11896 ( .A(ram[618]), .B(ram[634]), .S(n8795), .Z(n2753) );
  MUX2_X1 U11897 ( .A(ram[586]), .B(ram[602]), .S(n8795), .Z(n2754) );
  MUX2_X1 U11898 ( .A(n2754), .B(n2753), .S(n4232), .Z(n2755) );
  MUX2_X1 U11899 ( .A(ram[554]), .B(ram[570]), .S(n8795), .Z(n2756) );
  MUX2_X1 U11900 ( .A(ram[522]), .B(ram[538]), .S(n8795), .Z(n2757) );
  MUX2_X1 U11901 ( .A(n2757), .B(n2756), .S(n4232), .Z(n2758) );
  MUX2_X1 U11902 ( .A(n2758), .B(n2755), .S(n4149), .Z(n2759) );
  MUX2_X1 U11903 ( .A(n2759), .B(n2752), .S(n4102), .Z(n2760) );
  MUX2_X1 U11904 ( .A(n2760), .B(n2745), .S(n4083), .Z(n2761) );
  MUX2_X1 U11905 ( .A(ram[490]), .B(ram[506]), .S(n8795), .Z(n2762) );
  MUX2_X1 U11906 ( .A(ram[458]), .B(ram[474]), .S(n8795), .Z(n2763) );
  MUX2_X1 U11907 ( .A(n2763), .B(n2762), .S(n4232), .Z(n2764) );
  MUX2_X1 U11908 ( .A(ram[426]), .B(ram[442]), .S(n8795), .Z(n2765) );
  MUX2_X1 U11909 ( .A(ram[394]), .B(ram[410]), .S(n8795), .Z(n2766) );
  MUX2_X1 U11910 ( .A(n2766), .B(n2765), .S(n4232), .Z(n2767) );
  MUX2_X1 U11911 ( .A(n2767), .B(n2764), .S(n4149), .Z(n2768) );
  MUX2_X1 U11912 ( .A(ram[362]), .B(ram[378]), .S(n8795), .Z(n2769) );
  MUX2_X1 U11913 ( .A(ram[330]), .B(ram[346]), .S(n8795), .Z(n2770) );
  MUX2_X1 U11914 ( .A(n2770), .B(n2769), .S(n4232), .Z(n2771) );
  MUX2_X1 U11915 ( .A(ram[298]), .B(ram[314]), .S(n8795), .Z(n2772) );
  MUX2_X1 U11916 ( .A(ram[266]), .B(ram[282]), .S(n8795), .Z(n2773) );
  MUX2_X1 U11917 ( .A(n2773), .B(n2772), .S(n4232), .Z(n2774) );
  MUX2_X1 U11918 ( .A(n2774), .B(n2771), .S(n4149), .Z(n2775) );
  MUX2_X1 U11919 ( .A(n2775), .B(n2768), .S(n4102), .Z(n2776) );
  MUX2_X1 U11920 ( .A(ram[234]), .B(ram[250]), .S(n8796), .Z(n2777) );
  MUX2_X1 U11921 ( .A(ram[202]), .B(ram[218]), .S(n8796), .Z(n2778) );
  MUX2_X1 U11922 ( .A(n2778), .B(n2777), .S(n4233), .Z(n2779) );
  MUX2_X1 U11923 ( .A(ram[170]), .B(ram[186]), .S(n8796), .Z(n2780) );
  MUX2_X1 U11924 ( .A(ram[138]), .B(ram[154]), .S(n8796), .Z(n2781) );
  MUX2_X1 U11925 ( .A(n2781), .B(n2780), .S(n4233), .Z(n2782) );
  MUX2_X1 U11926 ( .A(n2782), .B(n2779), .S(n4149), .Z(n2783) );
  MUX2_X1 U11927 ( .A(ram[106]), .B(ram[122]), .S(n8796), .Z(n2784) );
  MUX2_X1 U11928 ( .A(ram[74]), .B(ram[90]), .S(n8796), .Z(n2785) );
  MUX2_X1 U11929 ( .A(n2785), .B(n2784), .S(n4233), .Z(n2786) );
  MUX2_X1 U11930 ( .A(ram[42]), .B(ram[58]), .S(n8796), .Z(n2787) );
  MUX2_X1 U11931 ( .A(ram[10]), .B(ram[26]), .S(n8796), .Z(n2788) );
  MUX2_X1 U11932 ( .A(n2788), .B(n2787), .S(n4233), .Z(n2789) );
  MUX2_X1 U11933 ( .A(n2789), .B(n2786), .S(n4149), .Z(n2790) );
  MUX2_X1 U11934 ( .A(n2790), .B(n2783), .S(n4102), .Z(n2791) );
  MUX2_X1 U11935 ( .A(n2791), .B(n2776), .S(n4083), .Z(n2792) );
  MUX2_X1 U11936 ( .A(n2792), .B(n2761), .S(n4072), .Z(n2793) );
  MUX2_X1 U11937 ( .A(n2793), .B(n2730), .S(n4067), .Z(n2794) );
  MUX2_X1 U11938 ( .A(n2794), .B(n2667), .S(mem_access_addr[9]), .Z(N291) );
  MUX2_X1 U11939 ( .A(ram[4075]), .B(ram[4091]), .S(n8796), .Z(n2795) );
  MUX2_X1 U11940 ( .A(ram[4043]), .B(ram[4059]), .S(n8796), .Z(n2796) );
  MUX2_X1 U11941 ( .A(n2796), .B(n2795), .S(n4233), .Z(n2797) );
  MUX2_X1 U11942 ( .A(ram[4011]), .B(ram[4027]), .S(n8796), .Z(n2798) );
  MUX2_X1 U11943 ( .A(ram[3979]), .B(ram[3995]), .S(n8796), .Z(n2799) );
  MUX2_X1 U11944 ( .A(n2799), .B(n2798), .S(n4233), .Z(n2800) );
  MUX2_X1 U11945 ( .A(n2800), .B(n2797), .S(n4149), .Z(n2801) );
  MUX2_X1 U11946 ( .A(ram[3947]), .B(ram[3963]), .S(n8797), .Z(n2802) );
  MUX2_X1 U11947 ( .A(ram[3915]), .B(ram[3931]), .S(n8797), .Z(n2803) );
  MUX2_X1 U11948 ( .A(n2803), .B(n2802), .S(n4233), .Z(n2804) );
  MUX2_X1 U11949 ( .A(ram[3883]), .B(ram[3899]), .S(n8797), .Z(n2805) );
  MUX2_X1 U11950 ( .A(ram[3851]), .B(ram[3867]), .S(n8797), .Z(n2806) );
  MUX2_X1 U11951 ( .A(n2806), .B(n2805), .S(n4233), .Z(n2807) );
  MUX2_X1 U11952 ( .A(n2807), .B(n2804), .S(n4149), .Z(n2808) );
  MUX2_X1 U11953 ( .A(n2808), .B(n2801), .S(n4102), .Z(n2809) );
  MUX2_X1 U11954 ( .A(ram[3819]), .B(ram[3835]), .S(n8797), .Z(n2810) );
  MUX2_X1 U11955 ( .A(ram[3787]), .B(ram[3803]), .S(n8797), .Z(n2811) );
  MUX2_X1 U11956 ( .A(n2811), .B(n2810), .S(n4233), .Z(n2812) );
  MUX2_X1 U11957 ( .A(ram[3755]), .B(ram[3771]), .S(n8797), .Z(n2813) );
  MUX2_X1 U11958 ( .A(ram[3723]), .B(ram[3739]), .S(n8797), .Z(n2814) );
  MUX2_X1 U11959 ( .A(n2814), .B(n2813), .S(n4233), .Z(n2815) );
  MUX2_X1 U11960 ( .A(n2815), .B(n2812), .S(n4149), .Z(n2816) );
  MUX2_X1 U11961 ( .A(ram[3691]), .B(ram[3707]), .S(n8797), .Z(n2817) );
  MUX2_X1 U11962 ( .A(ram[3659]), .B(ram[3675]), .S(n8797), .Z(n2818) );
  MUX2_X1 U11963 ( .A(n2818), .B(n2817), .S(n4233), .Z(n2819) );
  MUX2_X1 U11964 ( .A(ram[3627]), .B(ram[3643]), .S(n8797), .Z(n2820) );
  MUX2_X1 U11965 ( .A(ram[3595]), .B(ram[3611]), .S(n8797), .Z(n2821) );
  MUX2_X1 U11966 ( .A(n2821), .B(n2820), .S(n4233), .Z(n2822) );
  MUX2_X1 U11967 ( .A(n2822), .B(n2819), .S(n4149), .Z(n2823) );
  MUX2_X1 U11968 ( .A(n2823), .B(n2816), .S(n4102), .Z(n2824) );
  MUX2_X1 U11969 ( .A(n2824), .B(n2809), .S(n4083), .Z(n2825) );
  MUX2_X1 U11970 ( .A(ram[3563]), .B(ram[3579]), .S(n8798), .Z(n2826) );
  MUX2_X1 U11971 ( .A(ram[3531]), .B(ram[3547]), .S(n8798), .Z(n2827) );
  MUX2_X1 U11972 ( .A(n2827), .B(n2826), .S(n4234), .Z(n2828) );
  MUX2_X1 U11973 ( .A(ram[3499]), .B(ram[3515]), .S(n8798), .Z(n2829) );
  MUX2_X1 U11974 ( .A(ram[3467]), .B(ram[3483]), .S(n8798), .Z(n2830) );
  MUX2_X1 U11975 ( .A(n2830), .B(n2829), .S(n4234), .Z(n2831) );
  MUX2_X1 U11976 ( .A(n2831), .B(n2828), .S(n4150), .Z(n2832) );
  MUX2_X1 U11977 ( .A(ram[3435]), .B(ram[3451]), .S(n8798), .Z(n2833) );
  MUX2_X1 U11978 ( .A(ram[3403]), .B(ram[3419]), .S(n8798), .Z(n2834) );
  MUX2_X1 U11979 ( .A(n2834), .B(n2833), .S(n4234), .Z(n2835) );
  MUX2_X1 U11980 ( .A(ram[3371]), .B(ram[3387]), .S(n8798), .Z(n2836) );
  MUX2_X1 U11981 ( .A(ram[3339]), .B(ram[3355]), .S(n8798), .Z(n2837) );
  MUX2_X1 U11982 ( .A(n2837), .B(n2836), .S(n4234), .Z(n2838) );
  MUX2_X1 U11983 ( .A(n2838), .B(n2835), .S(n4150), .Z(n2839) );
  MUX2_X1 U11984 ( .A(n2839), .B(n2832), .S(n4102), .Z(n2840) );
  MUX2_X1 U11985 ( .A(ram[3307]), .B(ram[3323]), .S(n8798), .Z(n2841) );
  MUX2_X1 U11986 ( .A(ram[3275]), .B(ram[3291]), .S(n8798), .Z(n2842) );
  MUX2_X1 U11987 ( .A(n2842), .B(n2841), .S(n4234), .Z(n2843) );
  MUX2_X1 U11988 ( .A(ram[3243]), .B(ram[3259]), .S(n8798), .Z(n2844) );
  MUX2_X1 U11989 ( .A(ram[3211]), .B(ram[3227]), .S(n8798), .Z(n2845) );
  MUX2_X1 U11990 ( .A(n2845), .B(n2844), .S(n4234), .Z(n2846) );
  MUX2_X1 U11991 ( .A(n2846), .B(n2843), .S(n4150), .Z(n2847) );
  MUX2_X1 U11992 ( .A(ram[3179]), .B(ram[3195]), .S(n8799), .Z(n2848) );
  MUX2_X1 U11993 ( .A(ram[3147]), .B(ram[3163]), .S(n8799), .Z(n2849) );
  MUX2_X1 U11994 ( .A(n2849), .B(n2848), .S(n4234), .Z(n2850) );
  MUX2_X1 U11995 ( .A(ram[3115]), .B(ram[3131]), .S(n8799), .Z(n2851) );
  MUX2_X1 U11996 ( .A(ram[3083]), .B(ram[3099]), .S(n8799), .Z(n2852) );
  MUX2_X1 U11997 ( .A(n2852), .B(n2851), .S(n4234), .Z(n2853) );
  MUX2_X1 U11998 ( .A(n2853), .B(n2850), .S(n4150), .Z(n2854) );
  MUX2_X1 U11999 ( .A(n2854), .B(n2847), .S(n4102), .Z(n2855) );
  MUX2_X1 U12000 ( .A(n2855), .B(n2840), .S(n4083), .Z(n2856) );
  MUX2_X1 U12001 ( .A(n2856), .B(n2825), .S(n4072), .Z(n2857) );
  MUX2_X1 U12002 ( .A(ram[3051]), .B(ram[3067]), .S(n8799), .Z(n2858) );
  MUX2_X1 U12003 ( .A(ram[3019]), .B(ram[3035]), .S(n8799), .Z(n2859) );
  MUX2_X1 U12004 ( .A(n2859), .B(n2858), .S(n4234), .Z(n28601) );
  MUX2_X1 U12005 ( .A(ram[2987]), .B(ram[3003]), .S(n8799), .Z(n2861) );
  MUX2_X1 U12006 ( .A(ram[2955]), .B(ram[2971]), .S(n8799), .Z(n2862) );
  MUX2_X1 U12007 ( .A(n2862), .B(n2861), .S(n4234), .Z(n2863) );
  MUX2_X1 U12008 ( .A(n2863), .B(n28601), .S(n4150), .Z(n2864) );
  MUX2_X1 U12009 ( .A(ram[2923]), .B(ram[2939]), .S(n8799), .Z(n2865) );
  MUX2_X1 U12010 ( .A(ram[2891]), .B(ram[2907]), .S(n8799), .Z(n2866) );
  MUX2_X1 U12011 ( .A(n2866), .B(n2865), .S(n4234), .Z(n2867) );
  MUX2_X1 U12012 ( .A(ram[2859]), .B(ram[2875]), .S(n8799), .Z(n2868) );
  MUX2_X1 U12013 ( .A(ram[2827]), .B(ram[2843]), .S(n8799), .Z(n2869) );
  MUX2_X1 U12014 ( .A(n2869), .B(n2868), .S(n4234), .Z(n28701) );
  MUX2_X1 U12015 ( .A(n28701), .B(n2867), .S(n4150), .Z(n2871) );
  MUX2_X1 U12016 ( .A(n2871), .B(n2864), .S(n4102), .Z(n2872) );
  MUX2_X1 U12017 ( .A(ram[2795]), .B(ram[2811]), .S(n8800), .Z(n2873) );
  MUX2_X1 U12018 ( .A(ram[2763]), .B(ram[2779]), .S(n8800), .Z(n2874) );
  MUX2_X1 U12019 ( .A(n2874), .B(n2873), .S(n4235), .Z(n2875) );
  MUX2_X1 U12020 ( .A(ram[2731]), .B(ram[2747]), .S(n8800), .Z(n2876) );
  MUX2_X1 U12021 ( .A(ram[2699]), .B(ram[2715]), .S(n8800), .Z(n2877) );
  MUX2_X1 U12022 ( .A(n2877), .B(n2876), .S(n4235), .Z(n2878) );
  MUX2_X1 U12023 ( .A(n2878), .B(n2875), .S(n4150), .Z(n2879) );
  MUX2_X1 U12024 ( .A(ram[2667]), .B(ram[2683]), .S(n8800), .Z(n28801) );
  MUX2_X1 U12025 ( .A(ram[2635]), .B(ram[2651]), .S(n8800), .Z(n2881) );
  MUX2_X1 U12026 ( .A(n2881), .B(n28801), .S(n4235), .Z(n2882) );
  MUX2_X1 U12027 ( .A(ram[2603]), .B(ram[2619]), .S(n8800), .Z(n2883) );
  MUX2_X1 U12028 ( .A(ram[2571]), .B(ram[2587]), .S(n8800), .Z(n2884) );
  MUX2_X1 U12029 ( .A(n2884), .B(n2883), .S(n4235), .Z(n2885) );
  MUX2_X1 U12030 ( .A(n2885), .B(n2882), .S(n4150), .Z(n2886) );
  MUX2_X1 U12031 ( .A(n2886), .B(n2879), .S(n4102), .Z(n2887) );
  MUX2_X1 U12032 ( .A(n2887), .B(n2872), .S(n4083), .Z(n2888) );
  MUX2_X1 U12033 ( .A(ram[2539]), .B(ram[2555]), .S(n8800), .Z(n2889) );
  MUX2_X1 U12034 ( .A(ram[2507]), .B(ram[2523]), .S(n8800), .Z(n28901) );
  MUX2_X1 U12035 ( .A(n28901), .B(n2889), .S(n4235), .Z(n2891) );
  MUX2_X1 U12036 ( .A(ram[2475]), .B(ram[2491]), .S(n8800), .Z(n2892) );
  MUX2_X1 U12037 ( .A(ram[2443]), .B(ram[2459]), .S(n8800), .Z(n2893) );
  MUX2_X1 U12038 ( .A(n2893), .B(n2892), .S(n4235), .Z(n2894) );
  MUX2_X1 U12039 ( .A(n2894), .B(n2891), .S(n4150), .Z(n2895) );
  MUX2_X1 U12040 ( .A(ram[2411]), .B(ram[2427]), .S(n8801), .Z(n2896) );
  MUX2_X1 U12041 ( .A(ram[2379]), .B(ram[2395]), .S(n8801), .Z(n2897) );
  MUX2_X1 U12042 ( .A(n2897), .B(n2896), .S(n4235), .Z(n2898) );
  MUX2_X1 U12043 ( .A(ram[2347]), .B(ram[2363]), .S(n8801), .Z(n2899) );
  MUX2_X1 U12044 ( .A(ram[2315]), .B(ram[2331]), .S(n8801), .Z(n29001) );
  MUX2_X1 U12045 ( .A(n29001), .B(n2899), .S(n4235), .Z(n2901) );
  MUX2_X1 U12046 ( .A(n2901), .B(n2898), .S(n4150), .Z(n2902) );
  MUX2_X1 U12047 ( .A(n2902), .B(n2895), .S(n4102), .Z(n2903) );
  MUX2_X1 U12048 ( .A(ram[2283]), .B(ram[2299]), .S(n8801), .Z(n2904) );
  MUX2_X1 U12049 ( .A(ram[2251]), .B(ram[2267]), .S(n8801), .Z(n2905) );
  MUX2_X1 U12050 ( .A(n2905), .B(n2904), .S(n4235), .Z(n2906) );
  MUX2_X1 U12051 ( .A(ram[2219]), .B(ram[2235]), .S(n8801), .Z(n2907) );
  MUX2_X1 U12052 ( .A(ram[2187]), .B(ram[2203]), .S(n8801), .Z(n2908) );
  MUX2_X1 U12053 ( .A(n2908), .B(n2907), .S(n4235), .Z(n2909) );
  MUX2_X1 U12054 ( .A(n2909), .B(n2906), .S(n4150), .Z(n29101) );
  MUX2_X1 U12055 ( .A(ram[2155]), .B(ram[2171]), .S(n8801), .Z(n2911) );
  MUX2_X1 U12056 ( .A(ram[2123]), .B(ram[2139]), .S(n8801), .Z(n2912) );
  MUX2_X1 U12057 ( .A(n2912), .B(n2911), .S(n4235), .Z(n2913) );
  MUX2_X1 U12058 ( .A(ram[2091]), .B(ram[2107]), .S(n8801), .Z(n2914) );
  MUX2_X1 U12059 ( .A(ram[2059]), .B(ram[2075]), .S(n8801), .Z(n2915) );
  MUX2_X1 U12060 ( .A(n2915), .B(n2914), .S(n4235), .Z(n2916) );
  MUX2_X1 U12061 ( .A(n2916), .B(n2913), .S(n4150), .Z(n2917) );
  MUX2_X1 U12062 ( .A(n2917), .B(n29101), .S(n4102), .Z(n2918) );
  MUX2_X1 U12063 ( .A(n2918), .B(n2903), .S(n4083), .Z(n2919) );
  MUX2_X1 U12064 ( .A(n2919), .B(n2888), .S(n4072), .Z(n29201) );
  MUX2_X1 U12065 ( .A(n29201), .B(n2857), .S(n4067), .Z(n2921) );
  MUX2_X1 U12066 ( .A(ram[2027]), .B(ram[2043]), .S(n8802), .Z(n2922) );
  MUX2_X1 U12067 ( .A(ram[1995]), .B(ram[2011]), .S(n8802), .Z(n2923) );
  MUX2_X1 U12068 ( .A(n2923), .B(n2922), .S(n4236), .Z(n2924) );
  MUX2_X1 U12069 ( .A(ram[1963]), .B(ram[1979]), .S(n8802), .Z(n2925) );
  MUX2_X1 U12070 ( .A(ram[1931]), .B(ram[1947]), .S(n8802), .Z(n2926) );
  MUX2_X1 U12071 ( .A(n2926), .B(n2925), .S(n4236), .Z(n2927) );
  MUX2_X1 U12072 ( .A(n2927), .B(n2924), .S(n4151), .Z(n2928) );
  MUX2_X1 U12073 ( .A(ram[1899]), .B(ram[1915]), .S(n8802), .Z(n2929) );
  MUX2_X1 U12074 ( .A(ram[1867]), .B(ram[1883]), .S(n8802), .Z(n29301) );
  MUX2_X1 U12075 ( .A(n29301), .B(n2929), .S(n4236), .Z(n2931) );
  MUX2_X1 U12076 ( .A(ram[1835]), .B(ram[1851]), .S(n8802), .Z(n2932) );
  MUX2_X1 U12077 ( .A(ram[1803]), .B(ram[1819]), .S(n8802), .Z(n2933) );
  MUX2_X1 U12078 ( .A(n2933), .B(n2932), .S(n4236), .Z(n2934) );
  MUX2_X1 U12079 ( .A(n2934), .B(n2931), .S(n4151), .Z(n2935) );
  MUX2_X1 U12080 ( .A(n2935), .B(n2928), .S(n4103), .Z(n2936) );
  MUX2_X1 U12081 ( .A(ram[1771]), .B(ram[1787]), .S(n8802), .Z(n2937) );
  MUX2_X1 U12082 ( .A(ram[1739]), .B(ram[1755]), .S(n8802), .Z(n2938) );
  MUX2_X1 U12083 ( .A(n2938), .B(n2937), .S(n4236), .Z(n2939) );
  MUX2_X1 U12084 ( .A(ram[1707]), .B(ram[1723]), .S(n8802), .Z(n29401) );
  MUX2_X1 U12085 ( .A(ram[1675]), .B(ram[1691]), .S(n8802), .Z(n2941) );
  MUX2_X1 U12086 ( .A(n2941), .B(n29401), .S(n4236), .Z(n2942) );
  MUX2_X1 U12087 ( .A(n2942), .B(n2939), .S(n4151), .Z(n2943) );
  MUX2_X1 U12088 ( .A(ram[1643]), .B(ram[1659]), .S(n8803), .Z(n2944) );
  MUX2_X1 U12089 ( .A(ram[1611]), .B(ram[1627]), .S(n8803), .Z(n2945) );
  MUX2_X1 U12090 ( .A(n2945), .B(n2944), .S(n4236), .Z(n2946) );
  MUX2_X1 U12091 ( .A(ram[1579]), .B(ram[1595]), .S(n8803), .Z(n2947) );
  MUX2_X1 U12092 ( .A(ram[1547]), .B(ram[1563]), .S(n8803), .Z(n2948) );
  MUX2_X1 U12093 ( .A(n2948), .B(n2947), .S(n4236), .Z(n2949) );
  MUX2_X1 U12094 ( .A(n2949), .B(n2946), .S(n4151), .Z(n29501) );
  MUX2_X1 U12095 ( .A(n29501), .B(n2943), .S(n4103), .Z(n2951) );
  MUX2_X1 U12096 ( .A(n2951), .B(n2936), .S(n4084), .Z(n2952) );
  MUX2_X1 U12097 ( .A(ram[1515]), .B(ram[1531]), .S(n8803), .Z(n2953) );
  MUX2_X1 U12098 ( .A(ram[1483]), .B(ram[1499]), .S(n8803), .Z(n2954) );
  MUX2_X1 U12099 ( .A(n2954), .B(n2953), .S(n4236), .Z(n2955) );
  MUX2_X1 U12100 ( .A(ram[1451]), .B(ram[1467]), .S(n8803), .Z(n2956) );
  MUX2_X1 U12101 ( .A(ram[1419]), .B(ram[1435]), .S(n8803), .Z(n2957) );
  MUX2_X1 U12102 ( .A(n2957), .B(n2956), .S(n4236), .Z(n2958) );
  MUX2_X1 U12103 ( .A(n2958), .B(n2955), .S(n4151), .Z(n2959) );
  MUX2_X1 U12104 ( .A(ram[1387]), .B(ram[1403]), .S(n8803), .Z(n29601) );
  MUX2_X1 U12105 ( .A(ram[1355]), .B(ram[1371]), .S(n8803), .Z(n2961) );
  MUX2_X1 U12106 ( .A(n2961), .B(n29601), .S(n4236), .Z(n2962) );
  MUX2_X1 U12107 ( .A(ram[1323]), .B(ram[1339]), .S(n8803), .Z(n2963) );
  MUX2_X1 U12108 ( .A(ram[1291]), .B(ram[1307]), .S(n8803), .Z(n2964) );
  MUX2_X1 U12109 ( .A(n2964), .B(n2963), .S(n4236), .Z(n2965) );
  MUX2_X1 U12110 ( .A(n2965), .B(n2962), .S(n4151), .Z(n2966) );
  MUX2_X1 U12111 ( .A(n2966), .B(n2959), .S(n4103), .Z(n2967) );
  MUX2_X1 U12112 ( .A(ram[1259]), .B(ram[1275]), .S(n8804), .Z(n2968) );
  MUX2_X1 U12113 ( .A(ram[1227]), .B(ram[1243]), .S(n8804), .Z(n2969) );
  MUX2_X1 U12114 ( .A(n2969), .B(n2968), .S(n4237), .Z(n29701) );
  MUX2_X1 U12115 ( .A(ram[1195]), .B(ram[1211]), .S(n8804), .Z(n2971) );
  MUX2_X1 U12116 ( .A(ram[1163]), .B(ram[1179]), .S(n8804), .Z(n2972) );
  MUX2_X1 U12117 ( .A(n2972), .B(n2971), .S(n4237), .Z(n2973) );
  MUX2_X1 U12118 ( .A(n2973), .B(n29701), .S(n4151), .Z(n2974) );
  MUX2_X1 U12119 ( .A(ram[1131]), .B(ram[1147]), .S(n8804), .Z(n2975) );
  MUX2_X1 U12120 ( .A(ram[1099]), .B(ram[1115]), .S(n8804), .Z(n2976) );
  MUX2_X1 U12121 ( .A(n2976), .B(n2975), .S(n4237), .Z(n2977) );
  MUX2_X1 U12122 ( .A(ram[1067]), .B(ram[1083]), .S(n8804), .Z(n2978) );
  MUX2_X1 U12123 ( .A(ram[1035]), .B(ram[1051]), .S(n8804), .Z(n2979) );
  MUX2_X1 U12124 ( .A(n2979), .B(n2978), .S(n4237), .Z(n29801) );
  MUX2_X1 U12125 ( .A(n29801), .B(n2977), .S(n4151), .Z(n2981) );
  MUX2_X1 U12126 ( .A(n2981), .B(n2974), .S(n4103), .Z(n2982) );
  MUX2_X1 U12127 ( .A(n2982), .B(n2967), .S(n4084), .Z(n2983) );
  MUX2_X1 U12128 ( .A(n2983), .B(n2952), .S(n4072), .Z(n2984) );
  MUX2_X1 U12129 ( .A(ram[1003]), .B(ram[1019]), .S(n8804), .Z(n2985) );
  MUX2_X1 U12130 ( .A(ram[971]), .B(ram[987]), .S(n8804), .Z(n2986) );
  MUX2_X1 U12131 ( .A(n2986), .B(n2985), .S(n4237), .Z(n2987) );
  MUX2_X1 U12132 ( .A(ram[939]), .B(ram[955]), .S(n8804), .Z(n2988) );
  MUX2_X1 U12133 ( .A(ram[907]), .B(ram[923]), .S(n8804), .Z(n2989) );
  MUX2_X1 U12134 ( .A(n2989), .B(n2988), .S(n4237), .Z(n29901) );
  MUX2_X1 U12135 ( .A(n29901), .B(n2987), .S(n4151), .Z(n2991) );
  MUX2_X1 U12136 ( .A(ram[875]), .B(ram[891]), .S(n8805), .Z(n2992) );
  MUX2_X1 U12137 ( .A(ram[843]), .B(ram[859]), .S(n8805), .Z(n2993) );
  MUX2_X1 U12138 ( .A(n2993), .B(n2992), .S(n4237), .Z(n2994) );
  MUX2_X1 U12139 ( .A(ram[811]), .B(ram[827]), .S(n8805), .Z(n2995) );
  MUX2_X1 U12140 ( .A(ram[779]), .B(ram[795]), .S(n8805), .Z(n2996) );
  MUX2_X1 U12141 ( .A(n2996), .B(n2995), .S(n4237), .Z(n2997) );
  MUX2_X1 U12142 ( .A(n2997), .B(n2994), .S(n4151), .Z(n2998) );
  MUX2_X1 U12143 ( .A(n2998), .B(n2991), .S(n4103), .Z(n2999) );
  MUX2_X1 U12144 ( .A(ram[747]), .B(ram[763]), .S(n8805), .Z(n30001) );
  MUX2_X1 U12145 ( .A(ram[715]), .B(ram[731]), .S(n8805), .Z(n3001) );
  MUX2_X1 U12146 ( .A(n3001), .B(n30001), .S(n4237), .Z(n3002) );
  MUX2_X1 U12147 ( .A(ram[683]), .B(ram[699]), .S(n8805), .Z(n3003) );
  MUX2_X1 U12148 ( .A(ram[651]), .B(ram[667]), .S(n8805), .Z(n3004) );
  MUX2_X1 U12149 ( .A(n3004), .B(n3003), .S(n4237), .Z(n3005) );
  MUX2_X1 U12150 ( .A(n3005), .B(n3002), .S(n4151), .Z(n3006) );
  MUX2_X1 U12151 ( .A(ram[619]), .B(ram[635]), .S(n8805), .Z(n3007) );
  MUX2_X1 U12152 ( .A(ram[587]), .B(ram[603]), .S(n8805), .Z(n3008) );
  MUX2_X1 U12153 ( .A(n3008), .B(n3007), .S(n4237), .Z(n3009) );
  MUX2_X1 U12154 ( .A(ram[555]), .B(ram[571]), .S(n8805), .Z(n30101) );
  MUX2_X1 U12155 ( .A(ram[523]), .B(ram[539]), .S(n8805), .Z(n3011) );
  MUX2_X1 U12156 ( .A(n3011), .B(n30101), .S(n4237), .Z(n3012) );
  MUX2_X1 U12157 ( .A(n3012), .B(n3009), .S(n4151), .Z(n3013) );
  MUX2_X1 U12158 ( .A(n3013), .B(n3006), .S(n4103), .Z(n3014) );
  MUX2_X1 U12159 ( .A(n3014), .B(n2999), .S(n4084), .Z(n3015) );
  MUX2_X1 U12160 ( .A(ram[491]), .B(ram[507]), .S(n8806), .Z(n3016) );
  MUX2_X1 U12161 ( .A(ram[459]), .B(ram[475]), .S(n8806), .Z(n3017) );
  MUX2_X1 U12162 ( .A(n3017), .B(n3016), .S(n4238), .Z(n3018) );
  MUX2_X1 U12163 ( .A(ram[427]), .B(ram[443]), .S(n8806), .Z(n3019) );
  MUX2_X1 U12164 ( .A(ram[395]), .B(ram[411]), .S(n8806), .Z(n3020) );
  MUX2_X1 U12165 ( .A(n3020), .B(n3019), .S(n4238), .Z(n3021) );
  MUX2_X1 U12166 ( .A(n3021), .B(n3018), .S(n4152), .Z(n3022) );
  MUX2_X1 U12167 ( .A(ram[363]), .B(ram[379]), .S(n8806), .Z(n3023) );
  MUX2_X1 U12168 ( .A(ram[331]), .B(ram[347]), .S(n8806), .Z(n3024) );
  MUX2_X1 U12169 ( .A(n3024), .B(n3023), .S(n4238), .Z(n3025) );
  MUX2_X1 U12170 ( .A(ram[299]), .B(ram[315]), .S(n8806), .Z(n3026) );
  MUX2_X1 U12171 ( .A(ram[267]), .B(ram[283]), .S(n8806), .Z(n3027) );
  MUX2_X1 U12172 ( .A(n3027), .B(n3026), .S(n4238), .Z(n3028) );
  MUX2_X1 U12173 ( .A(n3028), .B(n3025), .S(n4152), .Z(n3029) );
  MUX2_X1 U12174 ( .A(n3029), .B(n3022), .S(n4103), .Z(n3030) );
  MUX2_X1 U12175 ( .A(ram[235]), .B(ram[251]), .S(n8806), .Z(n3031) );
  MUX2_X1 U12176 ( .A(ram[203]), .B(ram[219]), .S(n8806), .Z(n3032) );
  MUX2_X1 U12177 ( .A(n3032), .B(n3031), .S(n4238), .Z(n3033) );
  MUX2_X1 U12178 ( .A(ram[171]), .B(ram[187]), .S(n8806), .Z(n3034) );
  MUX2_X1 U12179 ( .A(ram[139]), .B(ram[155]), .S(n8806), .Z(n3035) );
  MUX2_X1 U12180 ( .A(n3035), .B(n3034), .S(n4238), .Z(n3036) );
  MUX2_X1 U12181 ( .A(n3036), .B(n3033), .S(n4152), .Z(n3037) );
  MUX2_X1 U12182 ( .A(ram[107]), .B(ram[123]), .S(n8807), .Z(n3038) );
  MUX2_X1 U12183 ( .A(ram[75]), .B(ram[91]), .S(n8807), .Z(n3039) );
  MUX2_X1 U12184 ( .A(n3039), .B(n3038), .S(n4238), .Z(n3040) );
  MUX2_X1 U12185 ( .A(ram[43]), .B(ram[59]), .S(n8807), .Z(n3041) );
  MUX2_X1 U12186 ( .A(ram[11]), .B(ram[27]), .S(n8807), .Z(n3042) );
  MUX2_X1 U12187 ( .A(n3042), .B(n3041), .S(n4238), .Z(n3043) );
  MUX2_X1 U12188 ( .A(n3043), .B(n3040), .S(n4152), .Z(n3044) );
  MUX2_X1 U12189 ( .A(n3044), .B(n3037), .S(n4103), .Z(n3045) );
  MUX2_X1 U12190 ( .A(n3045), .B(n3030), .S(n4084), .Z(n3046) );
  MUX2_X1 U12191 ( .A(n3046), .B(n3015), .S(n4072), .Z(n3047) );
  MUX2_X1 U12192 ( .A(n3047), .B(n2984), .S(n4067), .Z(n3048) );
  MUX2_X1 U12193 ( .A(n3048), .B(n2921), .S(mem_access_addr[9]), .Z(N290) );
  MUX2_X1 U12194 ( .A(ram[4076]), .B(ram[4092]), .S(n8807), .Z(n3049) );
  MUX2_X1 U12195 ( .A(ram[4044]), .B(ram[4060]), .S(n8807), .Z(n3050) );
  MUX2_X1 U12196 ( .A(n3050), .B(n3049), .S(n4238), .Z(n3051) );
  MUX2_X1 U12197 ( .A(ram[4012]), .B(ram[4028]), .S(n8807), .Z(n3052) );
  MUX2_X1 U12198 ( .A(ram[3980]), .B(ram[3996]), .S(n8807), .Z(n3053) );
  MUX2_X1 U12199 ( .A(n3053), .B(n3052), .S(n4238), .Z(n3054) );
  MUX2_X1 U12200 ( .A(n3054), .B(n3051), .S(n4152), .Z(n3055) );
  MUX2_X1 U12201 ( .A(ram[3948]), .B(ram[3964]), .S(n8807), .Z(n3056) );
  MUX2_X1 U12202 ( .A(ram[3916]), .B(ram[3932]), .S(n8807), .Z(n3057) );
  MUX2_X1 U12203 ( .A(n3057), .B(n3056), .S(n4238), .Z(n3058) );
  MUX2_X1 U12204 ( .A(ram[3884]), .B(ram[3900]), .S(n8807), .Z(n3059) );
  MUX2_X1 U12205 ( .A(ram[3852]), .B(ram[3868]), .S(n8807), .Z(n3060) );
  MUX2_X1 U12206 ( .A(n3060), .B(n3059), .S(n4238), .Z(n3061) );
  MUX2_X1 U12207 ( .A(n3061), .B(n3058), .S(n4152), .Z(n3062) );
  MUX2_X1 U12208 ( .A(n3062), .B(n3055), .S(n4103), .Z(n3063) );
  MUX2_X1 U12209 ( .A(ram[3820]), .B(ram[3836]), .S(n8808), .Z(n3064) );
  MUX2_X1 U12210 ( .A(ram[3788]), .B(ram[3804]), .S(n8808), .Z(n3065) );
  MUX2_X1 U12211 ( .A(n3065), .B(n3064), .S(n4239), .Z(n3066) );
  MUX2_X1 U12212 ( .A(ram[3756]), .B(ram[3772]), .S(n8808), .Z(n3067) );
  MUX2_X1 U12213 ( .A(ram[3724]), .B(ram[3740]), .S(n8808), .Z(n3068) );
  MUX2_X1 U12214 ( .A(n3068), .B(n3067), .S(n4239), .Z(n3069) );
  MUX2_X1 U12215 ( .A(n3069), .B(n3066), .S(n4152), .Z(n3070) );
  MUX2_X1 U12216 ( .A(ram[3692]), .B(ram[3708]), .S(n8808), .Z(n3071) );
  MUX2_X1 U12217 ( .A(ram[3660]), .B(ram[3676]), .S(n8808), .Z(n3072) );
  MUX2_X1 U12218 ( .A(n3072), .B(n3071), .S(n4239), .Z(n3073) );
  MUX2_X1 U12219 ( .A(ram[3628]), .B(ram[3644]), .S(n8808), .Z(n3074) );
  MUX2_X1 U12220 ( .A(ram[3596]), .B(ram[3612]), .S(n8808), .Z(n3075) );
  MUX2_X1 U12221 ( .A(n3075), .B(n3074), .S(n4239), .Z(n3076) );
  MUX2_X1 U12222 ( .A(n3076), .B(n3073), .S(n4152), .Z(n3077) );
  MUX2_X1 U12223 ( .A(n3077), .B(n3070), .S(n4103), .Z(n3078) );
  MUX2_X1 U12224 ( .A(n3078), .B(n3063), .S(n4084), .Z(n3079) );
  MUX2_X1 U12225 ( .A(ram[3564]), .B(ram[3580]), .S(n8808), .Z(n3080) );
  MUX2_X1 U12226 ( .A(ram[3532]), .B(ram[3548]), .S(n8808), .Z(n3081) );
  MUX2_X1 U12227 ( .A(n3081), .B(n3080), .S(n4239), .Z(n3082) );
  MUX2_X1 U12228 ( .A(ram[3500]), .B(ram[3516]), .S(n8808), .Z(n3083) );
  MUX2_X1 U12229 ( .A(ram[3468]), .B(ram[3484]), .S(n8808), .Z(n3084) );
  MUX2_X1 U12230 ( .A(n3084), .B(n3083), .S(n4239), .Z(n3085) );
  MUX2_X1 U12231 ( .A(n3085), .B(n3082), .S(n4152), .Z(n3086) );
  MUX2_X1 U12232 ( .A(ram[3436]), .B(ram[3452]), .S(n8809), .Z(n3087) );
  MUX2_X1 U12233 ( .A(ram[3404]), .B(ram[3420]), .S(n8809), .Z(n3088) );
  MUX2_X1 U12234 ( .A(n3088), .B(n3087), .S(n4239), .Z(n3089) );
  MUX2_X1 U12235 ( .A(ram[3372]), .B(ram[3388]), .S(n8809), .Z(n3090) );
  MUX2_X1 U12236 ( .A(ram[3340]), .B(ram[3356]), .S(n8809), .Z(n3091) );
  MUX2_X1 U12237 ( .A(n3091), .B(n3090), .S(n4239), .Z(n3092) );
  MUX2_X1 U12238 ( .A(n3092), .B(n3089), .S(n4152), .Z(n3093) );
  MUX2_X1 U12239 ( .A(n3093), .B(n3086), .S(n4103), .Z(n3094) );
  MUX2_X1 U12240 ( .A(ram[3308]), .B(ram[3324]), .S(n8809), .Z(n3095) );
  MUX2_X1 U12241 ( .A(ram[3276]), .B(ram[3292]), .S(n8809), .Z(n3096) );
  MUX2_X1 U12242 ( .A(n3096), .B(n3095), .S(n4239), .Z(n3097) );
  MUX2_X1 U12243 ( .A(ram[3244]), .B(ram[3260]), .S(n8809), .Z(n3098) );
  MUX2_X1 U12244 ( .A(ram[3212]), .B(ram[3228]), .S(n8809), .Z(n3099) );
  MUX2_X1 U12245 ( .A(n3099), .B(n3098), .S(n4239), .Z(n3100) );
  MUX2_X1 U12246 ( .A(n3100), .B(n3097), .S(n4152), .Z(n3101) );
  MUX2_X1 U12247 ( .A(ram[3180]), .B(ram[3196]), .S(n8809), .Z(n3102) );
  MUX2_X1 U12248 ( .A(ram[3148]), .B(ram[3164]), .S(n8809), .Z(n3103) );
  MUX2_X1 U12249 ( .A(n3103), .B(n3102), .S(n4239), .Z(n3104) );
  MUX2_X1 U12250 ( .A(ram[3116]), .B(ram[3132]), .S(n8809), .Z(n3105) );
  MUX2_X1 U12251 ( .A(ram[3084]), .B(ram[3100]), .S(n8809), .Z(n3106) );
  MUX2_X1 U12252 ( .A(n3106), .B(n3105), .S(n4239), .Z(n3107) );
  MUX2_X1 U12253 ( .A(n3107), .B(n3104), .S(n4152), .Z(n3108) );
  MUX2_X1 U12254 ( .A(n3108), .B(n3101), .S(n4103), .Z(n3109) );
  MUX2_X1 U12255 ( .A(n3109), .B(n3094), .S(n4084), .Z(n3110) );
  MUX2_X1 U12256 ( .A(n3110), .B(n3079), .S(n4072), .Z(n3111) );
  MUX2_X1 U12257 ( .A(ram[3052]), .B(ram[3068]), .S(n8810), .Z(n3112) );
  MUX2_X1 U12258 ( .A(ram[3020]), .B(ram[3036]), .S(n8810), .Z(n3113) );
  MUX2_X1 U12259 ( .A(n3113), .B(n3112), .S(n4240), .Z(n3114) );
  MUX2_X1 U12260 ( .A(ram[2988]), .B(ram[3004]), .S(n8810), .Z(n3115) );
  MUX2_X1 U12261 ( .A(ram[2956]), .B(ram[2972]), .S(n8810), .Z(n3116) );
  MUX2_X1 U12262 ( .A(n3116), .B(n3115), .S(n4240), .Z(n3117) );
  MUX2_X1 U12263 ( .A(n3117), .B(n3114), .S(n4153), .Z(n3118) );
  MUX2_X1 U12264 ( .A(ram[2924]), .B(ram[2940]), .S(n8810), .Z(n3119) );
  MUX2_X1 U12265 ( .A(ram[2892]), .B(ram[2908]), .S(n8810), .Z(n3120) );
  MUX2_X1 U12266 ( .A(n3120), .B(n3119), .S(n4240), .Z(n3121) );
  MUX2_X1 U12267 ( .A(ram[2860]), .B(ram[2876]), .S(n8810), .Z(n3122) );
  MUX2_X1 U12268 ( .A(ram[2828]), .B(ram[2844]), .S(n8810), .Z(n3123) );
  MUX2_X1 U12269 ( .A(n3123), .B(n3122), .S(n4240), .Z(n3124) );
  MUX2_X1 U12270 ( .A(n3124), .B(n3121), .S(n4153), .Z(n3125) );
  MUX2_X1 U12271 ( .A(n3125), .B(n3118), .S(n4104), .Z(n3126) );
  MUX2_X1 U12272 ( .A(ram[2796]), .B(ram[2812]), .S(n8810), .Z(n3127) );
  MUX2_X1 U12273 ( .A(ram[2764]), .B(ram[2780]), .S(n8810), .Z(n3128) );
  MUX2_X1 U12274 ( .A(n3128), .B(n3127), .S(n4240), .Z(n3129) );
  MUX2_X1 U12275 ( .A(ram[2732]), .B(ram[2748]), .S(n8810), .Z(n3130) );
  MUX2_X1 U12276 ( .A(ram[2700]), .B(ram[2716]), .S(n8810), .Z(n3131) );
  MUX2_X1 U12277 ( .A(n3131), .B(n3130), .S(n4240), .Z(n3132) );
  MUX2_X1 U12278 ( .A(n3132), .B(n3129), .S(n4153), .Z(n3133) );
  MUX2_X1 U12279 ( .A(ram[2668]), .B(ram[2684]), .S(n8811), .Z(n3134) );
  MUX2_X1 U12280 ( .A(ram[2636]), .B(ram[2652]), .S(n8811), .Z(n3135) );
  MUX2_X1 U12281 ( .A(n3135), .B(n3134), .S(n4240), .Z(n3136) );
  MUX2_X1 U12282 ( .A(ram[2604]), .B(ram[2620]), .S(n8811), .Z(n3137) );
  MUX2_X1 U12283 ( .A(ram[2572]), .B(ram[2588]), .S(n8811), .Z(n3138) );
  MUX2_X1 U12284 ( .A(n3138), .B(n3137), .S(n4240), .Z(n3139) );
  MUX2_X1 U12285 ( .A(n3139), .B(n3136), .S(n4153), .Z(n3140) );
  MUX2_X1 U12286 ( .A(n3140), .B(n3133), .S(n4104), .Z(n3141) );
  MUX2_X1 U12287 ( .A(n3141), .B(n3126), .S(n4084), .Z(n3142) );
  MUX2_X1 U12288 ( .A(ram[2540]), .B(ram[2556]), .S(n8811), .Z(n3143) );
  MUX2_X1 U12289 ( .A(ram[2508]), .B(ram[2524]), .S(n8811), .Z(n3144) );
  MUX2_X1 U12290 ( .A(n3144), .B(n3143), .S(n4240), .Z(n3145) );
  MUX2_X1 U12291 ( .A(ram[2476]), .B(ram[2492]), .S(n8811), .Z(n3146) );
  MUX2_X1 U12292 ( .A(ram[2444]), .B(ram[2460]), .S(n8811), .Z(n3147) );
  MUX2_X1 U12293 ( .A(n3147), .B(n3146), .S(n4240), .Z(n3148) );
  MUX2_X1 U12294 ( .A(n3148), .B(n3145), .S(n4153), .Z(n3149) );
  MUX2_X1 U12295 ( .A(ram[2412]), .B(ram[2428]), .S(n8811), .Z(n3150) );
  MUX2_X1 U12296 ( .A(ram[2380]), .B(ram[2396]), .S(n8811), .Z(n3151) );
  MUX2_X1 U12297 ( .A(n3151), .B(n3150), .S(n4240), .Z(n3152) );
  MUX2_X1 U12298 ( .A(ram[2348]), .B(ram[2364]), .S(n8811), .Z(n3153) );
  MUX2_X1 U12299 ( .A(ram[2316]), .B(ram[2332]), .S(n8811), .Z(n3154) );
  MUX2_X1 U12300 ( .A(n3154), .B(n3153), .S(n4240), .Z(n3155) );
  MUX2_X1 U12301 ( .A(n3155), .B(n3152), .S(n4153), .Z(n3156) );
  MUX2_X1 U12302 ( .A(n3156), .B(n3149), .S(n4104), .Z(n3157) );
  MUX2_X1 U12303 ( .A(ram[2284]), .B(ram[2300]), .S(n8812), .Z(n3158) );
  MUX2_X1 U12304 ( .A(ram[2252]), .B(ram[2268]), .S(n8812), .Z(n3159) );
  MUX2_X1 U12305 ( .A(n3159), .B(n3158), .S(n4241), .Z(n3160) );
  MUX2_X1 U12306 ( .A(ram[2220]), .B(ram[2236]), .S(n8812), .Z(n3161) );
  MUX2_X1 U12307 ( .A(ram[2188]), .B(ram[2204]), .S(n8812), .Z(n3162) );
  MUX2_X1 U12308 ( .A(n3162), .B(n3161), .S(n4241), .Z(n3163) );
  MUX2_X1 U12309 ( .A(n3163), .B(n3160), .S(n4153), .Z(n3164) );
  MUX2_X1 U12310 ( .A(ram[2156]), .B(ram[2172]), .S(n8812), .Z(n3165) );
  MUX2_X1 U12311 ( .A(ram[2124]), .B(ram[2140]), .S(n8812), .Z(n3166) );
  MUX2_X1 U12312 ( .A(n3166), .B(n3165), .S(n4241), .Z(n3167) );
  MUX2_X1 U12313 ( .A(ram[2092]), .B(ram[2108]), .S(n8812), .Z(n3168) );
  MUX2_X1 U12314 ( .A(ram[2060]), .B(ram[2076]), .S(n8812), .Z(n3169) );
  MUX2_X1 U12315 ( .A(n3169), .B(n3168), .S(n4241), .Z(n3170) );
  MUX2_X1 U12316 ( .A(n3170), .B(n3167), .S(n4153), .Z(n3171) );
  MUX2_X1 U12317 ( .A(n3171), .B(n3164), .S(n4104), .Z(n3172) );
  MUX2_X1 U12318 ( .A(n3172), .B(n3157), .S(n4084), .Z(n3173) );
  MUX2_X1 U12319 ( .A(n3173), .B(n3142), .S(n4072), .Z(n3174) );
  MUX2_X1 U12320 ( .A(n3174), .B(n3111), .S(n4067), .Z(n3175) );
  MUX2_X1 U12321 ( .A(ram[2028]), .B(ram[2044]), .S(n8812), .Z(n3176) );
  MUX2_X1 U12322 ( .A(ram[1996]), .B(ram[2012]), .S(n8812), .Z(n3177) );
  MUX2_X1 U12323 ( .A(n3177), .B(n3176), .S(n4241), .Z(n3178) );
  MUX2_X1 U12324 ( .A(ram[1964]), .B(ram[1980]), .S(n8812), .Z(n3179) );
  MUX2_X1 U12325 ( .A(ram[1932]), .B(ram[1948]), .S(n8812), .Z(n3180) );
  MUX2_X1 U12326 ( .A(n3180), .B(n3179), .S(n4241), .Z(n3181) );
  MUX2_X1 U12327 ( .A(n3181), .B(n3178), .S(n4153), .Z(n3182) );
  MUX2_X1 U12328 ( .A(ram[1900]), .B(ram[1916]), .S(n8813), .Z(n3183) );
  MUX2_X1 U12329 ( .A(ram[1868]), .B(ram[1884]), .S(n8813), .Z(n3184) );
  MUX2_X1 U12330 ( .A(n3184), .B(n3183), .S(n4241), .Z(n3185) );
  MUX2_X1 U12331 ( .A(ram[1836]), .B(ram[1852]), .S(n8813), .Z(n3186) );
  MUX2_X1 U12332 ( .A(ram[1804]), .B(ram[1820]), .S(n8813), .Z(n3187) );
  MUX2_X1 U12333 ( .A(n3187), .B(n3186), .S(n4241), .Z(n3188) );
  MUX2_X1 U12334 ( .A(n3188), .B(n3185), .S(n4153), .Z(n3189) );
  MUX2_X1 U12335 ( .A(n3189), .B(n3182), .S(n4104), .Z(n3190) );
  MUX2_X1 U12336 ( .A(ram[1772]), .B(ram[1788]), .S(n8813), .Z(n3191) );
  MUX2_X1 U12337 ( .A(ram[1740]), .B(ram[1756]), .S(n8813), .Z(n3192) );
  MUX2_X1 U12338 ( .A(n3192), .B(n3191), .S(n4241), .Z(n3193) );
  MUX2_X1 U12339 ( .A(ram[1708]), .B(ram[1724]), .S(n8813), .Z(n3194) );
  MUX2_X1 U12340 ( .A(ram[1676]), .B(ram[1692]), .S(n8813), .Z(n3195) );
  MUX2_X1 U12341 ( .A(n3195), .B(n3194), .S(n4241), .Z(n3196) );
  MUX2_X1 U12342 ( .A(n3196), .B(n3193), .S(n4153), .Z(n3197) );
  MUX2_X1 U12343 ( .A(ram[1644]), .B(ram[1660]), .S(n8813), .Z(n3198) );
  MUX2_X1 U12344 ( .A(ram[1612]), .B(ram[1628]), .S(n8813), .Z(n3199) );
  MUX2_X1 U12345 ( .A(n3199), .B(n3198), .S(n4241), .Z(n3200) );
  MUX2_X1 U12346 ( .A(ram[1580]), .B(ram[1596]), .S(n8813), .Z(n3201) );
  MUX2_X1 U12347 ( .A(ram[1548]), .B(ram[1564]), .S(n8813), .Z(n3202) );
  MUX2_X1 U12348 ( .A(n3202), .B(n3201), .S(n4241), .Z(n3203) );
  MUX2_X1 U12349 ( .A(n3203), .B(n3200), .S(n4153), .Z(n3204) );
  MUX2_X1 U12350 ( .A(n3204), .B(n3197), .S(n4104), .Z(n3205) );
  MUX2_X1 U12351 ( .A(n3205), .B(n3190), .S(n4084), .Z(n3206) );
  MUX2_X1 U12352 ( .A(ram[1516]), .B(ram[1532]), .S(n8814), .Z(n3207) );
  MUX2_X1 U12353 ( .A(ram[1484]), .B(ram[1500]), .S(n8814), .Z(n3208) );
  MUX2_X1 U12354 ( .A(n3208), .B(n3207), .S(n4242), .Z(n3209) );
  MUX2_X1 U12355 ( .A(ram[1452]), .B(ram[1468]), .S(n8814), .Z(n3210) );
  MUX2_X1 U12356 ( .A(ram[1420]), .B(ram[1436]), .S(n8814), .Z(n3211) );
  MUX2_X1 U12357 ( .A(n3211), .B(n3210), .S(n4242), .Z(n3212) );
  MUX2_X1 U12358 ( .A(n3212), .B(n3209), .S(n4154), .Z(n3213) );
  MUX2_X1 U12359 ( .A(ram[1388]), .B(ram[1404]), .S(n8814), .Z(n3214) );
  MUX2_X1 U12360 ( .A(ram[1356]), .B(ram[1372]), .S(n8814), .Z(n3215) );
  MUX2_X1 U12361 ( .A(n3215), .B(n3214), .S(n4242), .Z(n3216) );
  MUX2_X1 U12362 ( .A(ram[1324]), .B(ram[1340]), .S(n8814), .Z(n3217) );
  MUX2_X1 U12363 ( .A(ram[1292]), .B(ram[1308]), .S(n8814), .Z(n3218) );
  MUX2_X1 U12364 ( .A(n3218), .B(n3217), .S(n4242), .Z(n3219) );
  MUX2_X1 U12365 ( .A(n3219), .B(n3216), .S(n4154), .Z(n3220) );
  MUX2_X1 U12366 ( .A(n3220), .B(n3213), .S(n4104), .Z(n3221) );
  MUX2_X1 U12367 ( .A(ram[1260]), .B(ram[1276]), .S(n8814), .Z(n3222) );
  MUX2_X1 U12368 ( .A(ram[1228]), .B(ram[1244]), .S(n8814), .Z(n3223) );
  MUX2_X1 U12369 ( .A(n3223), .B(n3222), .S(n4242), .Z(n3224) );
  MUX2_X1 U12370 ( .A(ram[1196]), .B(ram[1212]), .S(n8814), .Z(n3225) );
  MUX2_X1 U12371 ( .A(ram[1164]), .B(ram[1180]), .S(n8814), .Z(n3226) );
  MUX2_X1 U12372 ( .A(n3226), .B(n3225), .S(n4242), .Z(n3227) );
  MUX2_X1 U12373 ( .A(n3227), .B(n3224), .S(n4154), .Z(n3228) );
  MUX2_X1 U12374 ( .A(ram[1132]), .B(ram[1148]), .S(n8815), .Z(n3229) );
  MUX2_X1 U12375 ( .A(ram[1100]), .B(ram[1116]), .S(n8815), .Z(n3230) );
  MUX2_X1 U12376 ( .A(n3230), .B(n3229), .S(n4242), .Z(n3231) );
  MUX2_X1 U12377 ( .A(ram[1068]), .B(ram[1084]), .S(n8815), .Z(n3232) );
  MUX2_X1 U12378 ( .A(ram[1036]), .B(ram[1052]), .S(n8815), .Z(n3233) );
  MUX2_X1 U12379 ( .A(n3233), .B(n3232), .S(n4242), .Z(n3234) );
  MUX2_X1 U12380 ( .A(n3234), .B(n3231), .S(n4154), .Z(n3235) );
  MUX2_X1 U12381 ( .A(n3235), .B(n3228), .S(n4104), .Z(n3236) );
  MUX2_X1 U12382 ( .A(n3236), .B(n3221), .S(n4084), .Z(n3237) );
  MUX2_X1 U12383 ( .A(n3237), .B(n3206), .S(n4072), .Z(n3238) );
  MUX2_X1 U12384 ( .A(ram[1004]), .B(ram[1020]), .S(n8815), .Z(n3239) );
  MUX2_X1 U12385 ( .A(ram[972]), .B(ram[988]), .S(n8815), .Z(n3240) );
  MUX2_X1 U12386 ( .A(n3240), .B(n3239), .S(n4242), .Z(n3241) );
  MUX2_X1 U12387 ( .A(ram[940]), .B(ram[956]), .S(n8815), .Z(n3242) );
  MUX2_X1 U12388 ( .A(ram[908]), .B(ram[924]), .S(n8815), .Z(n3243) );
  MUX2_X1 U12389 ( .A(n3243), .B(n3242), .S(n4242), .Z(n3244) );
  MUX2_X1 U12390 ( .A(n3244), .B(n3241), .S(n4154), .Z(n3245) );
  MUX2_X1 U12391 ( .A(ram[876]), .B(ram[892]), .S(n8815), .Z(n3246) );
  MUX2_X1 U12392 ( .A(ram[844]), .B(ram[860]), .S(n8815), .Z(n3247) );
  MUX2_X1 U12393 ( .A(n3247), .B(n3246), .S(n4242), .Z(n3248) );
  MUX2_X1 U12394 ( .A(ram[812]), .B(ram[828]), .S(n8815), .Z(n3249) );
  MUX2_X1 U12395 ( .A(ram[780]), .B(ram[796]), .S(n8815), .Z(n3250) );
  MUX2_X1 U12396 ( .A(n3250), .B(n3249), .S(n4242), .Z(n3251) );
  MUX2_X1 U12397 ( .A(n3251), .B(n3248), .S(n4154), .Z(n3252) );
  MUX2_X1 U12398 ( .A(n3252), .B(n3245), .S(n4104), .Z(n3253) );
  MUX2_X1 U12399 ( .A(ram[748]), .B(ram[764]), .S(n8816), .Z(n3254) );
  MUX2_X1 U12400 ( .A(ram[716]), .B(ram[732]), .S(n8816), .Z(n3255) );
  MUX2_X1 U12401 ( .A(n3255), .B(n3254), .S(n4243), .Z(n3256) );
  MUX2_X1 U12402 ( .A(ram[684]), .B(ram[700]), .S(n8816), .Z(n3257) );
  MUX2_X1 U12403 ( .A(ram[652]), .B(ram[668]), .S(n8816), .Z(n3258) );
  MUX2_X1 U12404 ( .A(n3258), .B(n3257), .S(n4243), .Z(n3259) );
  MUX2_X1 U12405 ( .A(n3259), .B(n3256), .S(n4154), .Z(n3260) );
  MUX2_X1 U12406 ( .A(ram[620]), .B(ram[636]), .S(n8816), .Z(n3261) );
  MUX2_X1 U12407 ( .A(ram[588]), .B(ram[604]), .S(n8816), .Z(n3262) );
  MUX2_X1 U12408 ( .A(n3262), .B(n3261), .S(n4243), .Z(n3263) );
  MUX2_X1 U12409 ( .A(ram[556]), .B(ram[572]), .S(n8816), .Z(n3264) );
  MUX2_X1 U12410 ( .A(ram[524]), .B(ram[540]), .S(n8816), .Z(n3265) );
  MUX2_X1 U12411 ( .A(n3265), .B(n3264), .S(n4243), .Z(n3266) );
  MUX2_X1 U12412 ( .A(n3266), .B(n3263), .S(n4154), .Z(n3267) );
  MUX2_X1 U12413 ( .A(n3267), .B(n3260), .S(n4104), .Z(n3268) );
  MUX2_X1 U12414 ( .A(n3268), .B(n3253), .S(n4084), .Z(n3269) );
  MUX2_X1 U12415 ( .A(ram[492]), .B(ram[508]), .S(n8816), .Z(n3270) );
  MUX2_X1 U12416 ( .A(ram[460]), .B(ram[476]), .S(n8816), .Z(n3271) );
  MUX2_X1 U12417 ( .A(n3271), .B(n3270), .S(n4243), .Z(n3272) );
  MUX2_X1 U12418 ( .A(ram[428]), .B(ram[444]), .S(n8816), .Z(n3273) );
  MUX2_X1 U12419 ( .A(ram[396]), .B(ram[412]), .S(n8816), .Z(n3274) );
  MUX2_X1 U12420 ( .A(n3274), .B(n3273), .S(n4243), .Z(n3275) );
  MUX2_X1 U12421 ( .A(n3275), .B(n3272), .S(n4154), .Z(n3276) );
  MUX2_X1 U12422 ( .A(ram[364]), .B(ram[380]), .S(n8817), .Z(n3277) );
  MUX2_X1 U12423 ( .A(ram[332]), .B(ram[348]), .S(n8817), .Z(n3278) );
  MUX2_X1 U12424 ( .A(n3278), .B(n3277), .S(n4243), .Z(n3279) );
  MUX2_X1 U12425 ( .A(ram[300]), .B(ram[316]), .S(n8817), .Z(n3280) );
  MUX2_X1 U12426 ( .A(ram[268]), .B(ram[284]), .S(n8817), .Z(n3281) );
  MUX2_X1 U12427 ( .A(n3281), .B(n3280), .S(n4243), .Z(n3282) );
  MUX2_X1 U12428 ( .A(n3282), .B(n3279), .S(n4154), .Z(n3283) );
  MUX2_X1 U12429 ( .A(n3283), .B(n3276), .S(n4104), .Z(n3284) );
  MUX2_X1 U12430 ( .A(ram[236]), .B(ram[252]), .S(n8817), .Z(n3285) );
  MUX2_X1 U12431 ( .A(ram[204]), .B(ram[220]), .S(n8817), .Z(n3286) );
  MUX2_X1 U12432 ( .A(n3286), .B(n3285), .S(n4243), .Z(n3287) );
  MUX2_X1 U12433 ( .A(ram[172]), .B(ram[188]), .S(n8817), .Z(n3288) );
  MUX2_X1 U12434 ( .A(ram[140]), .B(ram[156]), .S(n8817), .Z(n3289) );
  MUX2_X1 U12435 ( .A(n3289), .B(n3288), .S(n4243), .Z(n3290) );
  MUX2_X1 U12436 ( .A(n3290), .B(n3287), .S(n4154), .Z(n3291) );
  MUX2_X1 U12437 ( .A(ram[108]), .B(ram[124]), .S(n8817), .Z(n3292) );
  MUX2_X1 U12438 ( .A(ram[76]), .B(ram[92]), .S(n8817), .Z(n3293) );
  MUX2_X1 U12439 ( .A(n3293), .B(n3292), .S(n4243), .Z(n3294) );
  MUX2_X1 U12440 ( .A(ram[44]), .B(ram[60]), .S(n8817), .Z(n3295) );
  MUX2_X1 U12441 ( .A(ram[12]), .B(ram[28]), .S(n8817), .Z(n3296) );
  MUX2_X1 U12442 ( .A(n3296), .B(n3295), .S(n4243), .Z(n3297) );
  MUX2_X1 U12443 ( .A(n3297), .B(n3294), .S(n4154), .Z(n3298) );
  MUX2_X1 U12444 ( .A(n3298), .B(n3291), .S(n4104), .Z(n3299) );
  MUX2_X1 U12445 ( .A(n3299), .B(n3284), .S(n4084), .Z(n3300) );
  MUX2_X1 U12446 ( .A(n3300), .B(n3269), .S(n4072), .Z(n3301) );
  MUX2_X1 U12447 ( .A(n3301), .B(n3238), .S(n4067), .Z(n3302) );
  MUX2_X1 U12448 ( .A(n3302), .B(n3175), .S(mem_access_addr[9]), .Z(N289) );
  MUX2_X1 U12449 ( .A(ram[4077]), .B(ram[4093]), .S(n8818), .Z(n3303) );
  MUX2_X1 U12450 ( .A(ram[4045]), .B(ram[4061]), .S(n8818), .Z(n3304) );
  MUX2_X1 U12451 ( .A(n3304), .B(n3303), .S(n4244), .Z(n3305) );
  MUX2_X1 U12452 ( .A(ram[4013]), .B(ram[4029]), .S(n8818), .Z(n3306) );
  MUX2_X1 U12453 ( .A(ram[3981]), .B(ram[3997]), .S(n8818), .Z(n3307) );
  MUX2_X1 U12454 ( .A(n3307), .B(n3306), .S(n4244), .Z(n3308) );
  MUX2_X1 U12455 ( .A(n3308), .B(n3305), .S(n4155), .Z(n3309) );
  MUX2_X1 U12456 ( .A(ram[3949]), .B(ram[3965]), .S(n8818), .Z(n3310) );
  MUX2_X1 U12457 ( .A(ram[3917]), .B(ram[3933]), .S(n8818), .Z(n3311) );
  MUX2_X1 U12458 ( .A(n3311), .B(n3310), .S(n4244), .Z(n3312) );
  MUX2_X1 U12459 ( .A(ram[3885]), .B(ram[3901]), .S(n8818), .Z(n3313) );
  MUX2_X1 U12460 ( .A(ram[3853]), .B(ram[3869]), .S(n8818), .Z(n3314) );
  MUX2_X1 U12461 ( .A(n3314), .B(n3313), .S(n4244), .Z(n3315) );
  MUX2_X1 U12462 ( .A(n3315), .B(n3312), .S(n4155), .Z(n3316) );
  MUX2_X1 U12463 ( .A(n3316), .B(n3309), .S(n4105), .Z(n3317) );
  MUX2_X1 U12464 ( .A(ram[3821]), .B(ram[3837]), .S(n8818), .Z(n3318) );
  MUX2_X1 U12465 ( .A(ram[3789]), .B(ram[3805]), .S(n8818), .Z(n3319) );
  MUX2_X1 U12466 ( .A(n3319), .B(n3318), .S(n4244), .Z(n3320) );
  MUX2_X1 U12467 ( .A(ram[3757]), .B(ram[3773]), .S(n8818), .Z(n3321) );
  MUX2_X1 U12468 ( .A(ram[3725]), .B(ram[3741]), .S(n8818), .Z(n3322) );
  MUX2_X1 U12469 ( .A(n3322), .B(n3321), .S(n4244), .Z(n3323) );
  MUX2_X1 U12470 ( .A(n3323), .B(n3320), .S(n4155), .Z(n3324) );
  MUX2_X1 U12471 ( .A(ram[3693]), .B(ram[3709]), .S(n8819), .Z(n3325) );
  MUX2_X1 U12472 ( .A(ram[3661]), .B(ram[3677]), .S(n8819), .Z(n3326) );
  MUX2_X1 U12473 ( .A(n3326), .B(n3325), .S(n4244), .Z(n3327) );
  MUX2_X1 U12474 ( .A(ram[3629]), .B(ram[3645]), .S(n8819), .Z(n3328) );
  MUX2_X1 U12475 ( .A(ram[3597]), .B(ram[3613]), .S(n8819), .Z(n3329) );
  MUX2_X1 U12476 ( .A(n3329), .B(n3328), .S(n4244), .Z(n3330) );
  MUX2_X1 U12477 ( .A(n3330), .B(n3327), .S(n4155), .Z(n3331) );
  MUX2_X1 U12478 ( .A(n3331), .B(n3324), .S(n4105), .Z(n3332) );
  MUX2_X1 U12479 ( .A(n3332), .B(n3317), .S(n4085), .Z(n3333) );
  MUX2_X1 U12480 ( .A(ram[3565]), .B(ram[3581]), .S(n8819), .Z(n3334) );
  MUX2_X1 U12481 ( .A(ram[3533]), .B(ram[3549]), .S(n8819), .Z(n3335) );
  MUX2_X1 U12482 ( .A(n3335), .B(n3334), .S(n4244), .Z(n3336) );
  MUX2_X1 U12483 ( .A(ram[3501]), .B(ram[3517]), .S(n8819), .Z(n3337) );
  MUX2_X1 U12484 ( .A(ram[3469]), .B(ram[3485]), .S(n8819), .Z(n3338) );
  MUX2_X1 U12485 ( .A(n3338), .B(n3337), .S(n4244), .Z(n3339) );
  MUX2_X1 U12486 ( .A(n3339), .B(n3336), .S(n4155), .Z(n3340) );
  MUX2_X1 U12487 ( .A(ram[3437]), .B(ram[3453]), .S(n8819), .Z(n3341) );
  MUX2_X1 U12488 ( .A(ram[3405]), .B(ram[3421]), .S(n8819), .Z(n3342) );
  MUX2_X1 U12489 ( .A(n3342), .B(n3341), .S(n4244), .Z(n3343) );
  MUX2_X1 U12490 ( .A(ram[3373]), .B(ram[3389]), .S(n8819), .Z(n3344) );
  MUX2_X1 U12491 ( .A(ram[3341]), .B(ram[3357]), .S(n8819), .Z(n3345) );
  MUX2_X1 U12492 ( .A(n3345), .B(n3344), .S(n4244), .Z(n3346) );
  MUX2_X1 U12493 ( .A(n3346), .B(n3343), .S(n4155), .Z(n3347) );
  MUX2_X1 U12494 ( .A(n3347), .B(n3340), .S(n4105), .Z(n3348) );
  MUX2_X1 U12495 ( .A(ram[3309]), .B(ram[3325]), .S(n8820), .Z(n3349) );
  MUX2_X1 U12496 ( .A(ram[3277]), .B(ram[3293]), .S(n8820), .Z(n3350) );
  MUX2_X1 U12497 ( .A(n3350), .B(n3349), .S(n4245), .Z(n3351) );
  MUX2_X1 U12498 ( .A(ram[3245]), .B(ram[3261]), .S(n8820), .Z(n3352) );
  MUX2_X1 U12499 ( .A(ram[3213]), .B(ram[3229]), .S(n8820), .Z(n3353) );
  MUX2_X1 U12500 ( .A(n3353), .B(n3352), .S(n4245), .Z(n3354) );
  MUX2_X1 U12501 ( .A(n3354), .B(n3351), .S(n4155), .Z(n3355) );
  MUX2_X1 U12502 ( .A(ram[3181]), .B(ram[3197]), .S(n8820), .Z(n3356) );
  MUX2_X1 U12503 ( .A(ram[3149]), .B(ram[3165]), .S(n8820), .Z(n3357) );
  MUX2_X1 U12504 ( .A(n3357), .B(n3356), .S(n4245), .Z(n3358) );
  MUX2_X1 U12505 ( .A(ram[3117]), .B(ram[3133]), .S(n8820), .Z(n3359) );
  MUX2_X1 U12506 ( .A(ram[3085]), .B(ram[3101]), .S(n8820), .Z(n3360) );
  MUX2_X1 U12507 ( .A(n3360), .B(n3359), .S(n4245), .Z(n3361) );
  MUX2_X1 U12508 ( .A(n3361), .B(n3358), .S(n4155), .Z(n3362) );
  MUX2_X1 U12509 ( .A(n3362), .B(n3355), .S(n4105), .Z(n3363) );
  MUX2_X1 U12510 ( .A(n3363), .B(n3348), .S(n4085), .Z(n3364) );
  MUX2_X1 U12511 ( .A(n3364), .B(n3333), .S(n4073), .Z(n3365) );
  MUX2_X1 U12512 ( .A(ram[3053]), .B(ram[3069]), .S(n8820), .Z(n3366) );
  MUX2_X1 U12513 ( .A(ram[3021]), .B(ram[3037]), .S(n8820), .Z(n3367) );
  MUX2_X1 U12514 ( .A(n3367), .B(n3366), .S(n4245), .Z(n3368) );
  MUX2_X1 U12515 ( .A(ram[2989]), .B(ram[3005]), .S(n8820), .Z(n3369) );
  MUX2_X1 U12516 ( .A(ram[2957]), .B(ram[2973]), .S(n8820), .Z(n3370) );
  MUX2_X1 U12517 ( .A(n3370), .B(n3369), .S(n4245), .Z(n3371) );
  MUX2_X1 U12518 ( .A(n3371), .B(n3368), .S(n4155), .Z(n3372) );
  MUX2_X1 U12519 ( .A(ram[2925]), .B(ram[2941]), .S(n8821), .Z(n3373) );
  MUX2_X1 U12520 ( .A(ram[2893]), .B(ram[2909]), .S(n8821), .Z(n3374) );
  MUX2_X1 U12521 ( .A(n3374), .B(n3373), .S(n4245), .Z(n3375) );
  MUX2_X1 U12522 ( .A(ram[2861]), .B(ram[2877]), .S(n8821), .Z(n3376) );
  MUX2_X1 U12523 ( .A(ram[2829]), .B(ram[2845]), .S(n8821), .Z(n3377) );
  MUX2_X1 U12524 ( .A(n3377), .B(n3376), .S(n4245), .Z(n3378) );
  MUX2_X1 U12525 ( .A(n3378), .B(n3375), .S(n4155), .Z(n3379) );
  MUX2_X1 U12526 ( .A(n3379), .B(n3372), .S(n4105), .Z(n3380) );
  MUX2_X1 U12527 ( .A(ram[2797]), .B(ram[2813]), .S(n8821), .Z(n3381) );
  MUX2_X1 U12528 ( .A(ram[2765]), .B(ram[2781]), .S(n8821), .Z(n3382) );
  MUX2_X1 U12529 ( .A(n3382), .B(n3381), .S(n4245), .Z(n3383) );
  MUX2_X1 U12530 ( .A(ram[2733]), .B(ram[2749]), .S(n8821), .Z(n3384) );
  MUX2_X1 U12531 ( .A(ram[2701]), .B(ram[2717]), .S(n8821), .Z(n3385) );
  MUX2_X1 U12532 ( .A(n3385), .B(n3384), .S(n4245), .Z(n3386) );
  MUX2_X1 U12533 ( .A(n3386), .B(n3383), .S(n4155), .Z(n3387) );
  MUX2_X1 U12534 ( .A(ram[2669]), .B(ram[2685]), .S(n8821), .Z(n3388) );
  MUX2_X1 U12535 ( .A(ram[2637]), .B(ram[2653]), .S(n8821), .Z(n3389) );
  MUX2_X1 U12536 ( .A(n3389), .B(n3388), .S(n4245), .Z(n3390) );
  MUX2_X1 U12537 ( .A(ram[2605]), .B(ram[2621]), .S(n8821), .Z(n3391) );
  MUX2_X1 U12538 ( .A(ram[2573]), .B(ram[2589]), .S(n8821), .Z(n3392) );
  MUX2_X1 U12539 ( .A(n3392), .B(n3391), .S(n4245), .Z(n3393) );
  MUX2_X1 U12540 ( .A(n3393), .B(n3390), .S(n4155), .Z(n3394) );
  MUX2_X1 U12541 ( .A(n3394), .B(n3387), .S(n4105), .Z(n3395) );
  MUX2_X1 U12542 ( .A(n3395), .B(n3380), .S(n4085), .Z(n3396) );
  MUX2_X1 U12543 ( .A(ram[2541]), .B(ram[2557]), .S(n8822), .Z(n3397) );
  MUX2_X1 U12544 ( .A(ram[2509]), .B(ram[2525]), .S(n8822), .Z(n3398) );
  MUX2_X1 U12545 ( .A(n3398), .B(n3397), .S(n4246), .Z(n3399) );
  MUX2_X1 U12546 ( .A(ram[2477]), .B(ram[2493]), .S(n8822), .Z(n3400) );
  MUX2_X1 U12547 ( .A(ram[2445]), .B(ram[2461]), .S(n8822), .Z(n3401) );
  MUX2_X1 U12548 ( .A(n3401), .B(n3400), .S(n4246), .Z(n3402) );
  MUX2_X1 U12549 ( .A(n3402), .B(n3399), .S(n4156), .Z(n3403) );
  MUX2_X1 U12550 ( .A(ram[2413]), .B(ram[2429]), .S(n8822), .Z(n3404) );
  MUX2_X1 U12551 ( .A(ram[2381]), .B(ram[2397]), .S(n8822), .Z(n3405) );
  MUX2_X1 U12552 ( .A(n3405), .B(n3404), .S(n4246), .Z(n3406) );
  MUX2_X1 U12553 ( .A(ram[2349]), .B(ram[2365]), .S(n8822), .Z(n3407) );
  MUX2_X1 U12554 ( .A(ram[2317]), .B(ram[2333]), .S(n8822), .Z(n3408) );
  MUX2_X1 U12555 ( .A(n3408), .B(n3407), .S(n4246), .Z(n3409) );
  MUX2_X1 U12556 ( .A(n3409), .B(n3406), .S(n4156), .Z(n3410) );
  MUX2_X1 U12557 ( .A(n3410), .B(n3403), .S(n4105), .Z(n3411) );
  MUX2_X1 U12558 ( .A(ram[2285]), .B(ram[2301]), .S(n8822), .Z(n3412) );
  MUX2_X1 U12559 ( .A(ram[2253]), .B(ram[2269]), .S(n8822), .Z(n3413) );
  MUX2_X1 U12560 ( .A(n3413), .B(n3412), .S(n4246), .Z(n3414) );
  MUX2_X1 U12561 ( .A(ram[2221]), .B(ram[2237]), .S(n8822), .Z(n3415) );
  MUX2_X1 U12562 ( .A(ram[2189]), .B(ram[2205]), .S(n8822), .Z(n3416) );
  MUX2_X1 U12563 ( .A(n3416), .B(n3415), .S(n4246), .Z(n3417) );
  MUX2_X1 U12564 ( .A(n3417), .B(n3414), .S(n4156), .Z(n3418) );
  MUX2_X1 U12565 ( .A(ram[2157]), .B(ram[2173]), .S(n8823), .Z(n3419) );
  MUX2_X1 U12566 ( .A(ram[2125]), .B(ram[2141]), .S(n8823), .Z(n3420) );
  MUX2_X1 U12567 ( .A(n3420), .B(n3419), .S(n4246), .Z(n3421) );
  MUX2_X1 U12568 ( .A(ram[2093]), .B(ram[2109]), .S(n8823), .Z(n3422) );
  MUX2_X1 U12569 ( .A(ram[2061]), .B(ram[2077]), .S(n8823), .Z(n3423) );
  MUX2_X1 U12570 ( .A(n3423), .B(n3422), .S(n4246), .Z(n3424) );
  MUX2_X1 U12571 ( .A(n3424), .B(n3421), .S(n4156), .Z(n3425) );
  MUX2_X1 U12572 ( .A(n3425), .B(n3418), .S(n4105), .Z(n3426) );
  MUX2_X1 U12573 ( .A(n3426), .B(n3411), .S(n4085), .Z(n3427) );
  MUX2_X1 U12574 ( .A(n3427), .B(n3396), .S(n4073), .Z(n3428) );
  MUX2_X1 U12575 ( .A(n3428), .B(n3365), .S(n4067), .Z(n3429) );
  MUX2_X1 U12576 ( .A(ram[2029]), .B(ram[2045]), .S(n8823), .Z(n3430) );
  MUX2_X1 U12577 ( .A(ram[1997]), .B(ram[2013]), .S(n8823), .Z(n3431) );
  MUX2_X1 U12578 ( .A(n3431), .B(n3430), .S(n4246), .Z(n3432) );
  MUX2_X1 U12579 ( .A(ram[1965]), .B(ram[1981]), .S(n8823), .Z(n3433) );
  MUX2_X1 U12580 ( .A(ram[1933]), .B(ram[1949]), .S(n8823), .Z(n3434) );
  MUX2_X1 U12581 ( .A(n3434), .B(n3433), .S(n4246), .Z(n3435) );
  MUX2_X1 U12582 ( .A(n3435), .B(n3432), .S(n4156), .Z(n3436) );
  MUX2_X1 U12583 ( .A(ram[1901]), .B(ram[1917]), .S(n8823), .Z(n3437) );
  MUX2_X1 U12584 ( .A(ram[1869]), .B(ram[1885]), .S(n8823), .Z(n3438) );
  MUX2_X1 U12585 ( .A(n3438), .B(n3437), .S(n4246), .Z(n3439) );
  MUX2_X1 U12586 ( .A(ram[1837]), .B(ram[1853]), .S(n8823), .Z(n3440) );
  MUX2_X1 U12587 ( .A(ram[1805]), .B(ram[1821]), .S(n8823), .Z(n3441) );
  MUX2_X1 U12588 ( .A(n3441), .B(n3440), .S(n4246), .Z(n3442) );
  MUX2_X1 U12589 ( .A(n3442), .B(n3439), .S(n4156), .Z(n3443) );
  MUX2_X1 U12590 ( .A(n3443), .B(n3436), .S(n4105), .Z(n3444) );
  MUX2_X1 U12591 ( .A(ram[1773]), .B(ram[1789]), .S(n8824), .Z(n3445) );
  MUX2_X1 U12592 ( .A(ram[1741]), .B(ram[1757]), .S(n8824), .Z(n3446) );
  MUX2_X1 U12593 ( .A(n3446), .B(n3445), .S(n4247), .Z(n3447) );
  MUX2_X1 U12594 ( .A(ram[1709]), .B(ram[1725]), .S(n8824), .Z(n3448) );
  MUX2_X1 U12595 ( .A(ram[1677]), .B(ram[1693]), .S(n8824), .Z(n3449) );
  MUX2_X1 U12596 ( .A(n3449), .B(n3448), .S(n4247), .Z(n3450) );
  MUX2_X1 U12597 ( .A(n3450), .B(n3447), .S(n4156), .Z(n3451) );
  MUX2_X1 U12598 ( .A(ram[1645]), .B(ram[1661]), .S(n8824), .Z(n3452) );
  MUX2_X1 U12599 ( .A(ram[1613]), .B(ram[1629]), .S(n8824), .Z(n3453) );
  MUX2_X1 U12600 ( .A(n3453), .B(n3452), .S(n4247), .Z(n3454) );
  MUX2_X1 U12601 ( .A(ram[1581]), .B(ram[1597]), .S(n8824), .Z(n3455) );
  MUX2_X1 U12602 ( .A(ram[1549]), .B(ram[1565]), .S(n8824), .Z(n3456) );
  MUX2_X1 U12603 ( .A(n3456), .B(n3455), .S(n4247), .Z(n3457) );
  MUX2_X1 U12604 ( .A(n3457), .B(n3454), .S(n4156), .Z(n3458) );
  MUX2_X1 U12605 ( .A(n3458), .B(n3451), .S(n4105), .Z(n3459) );
  MUX2_X1 U12606 ( .A(n3459), .B(n3444), .S(n4085), .Z(n3460) );
  MUX2_X1 U12607 ( .A(ram[1517]), .B(ram[1533]), .S(n8824), .Z(n3461) );
  MUX2_X1 U12608 ( .A(ram[1485]), .B(ram[1501]), .S(n8824), .Z(n3462) );
  MUX2_X1 U12609 ( .A(n3462), .B(n3461), .S(n4247), .Z(n3463) );
  MUX2_X1 U12610 ( .A(ram[1453]), .B(ram[1469]), .S(n8824), .Z(n3464) );
  MUX2_X1 U12611 ( .A(ram[1421]), .B(ram[1437]), .S(n8824), .Z(n3465) );
  MUX2_X1 U12612 ( .A(n3465), .B(n3464), .S(n4247), .Z(n3466) );
  MUX2_X1 U12613 ( .A(n3466), .B(n3463), .S(n4156), .Z(n3467) );
  MUX2_X1 U12614 ( .A(ram[1389]), .B(ram[1405]), .S(n8825), .Z(n3468) );
  MUX2_X1 U12615 ( .A(ram[1357]), .B(ram[1373]), .S(n8825), .Z(n3469) );
  MUX2_X1 U12616 ( .A(n3469), .B(n3468), .S(n4247), .Z(n3470) );
  MUX2_X1 U12617 ( .A(ram[1325]), .B(ram[1341]), .S(n8825), .Z(n3471) );
  MUX2_X1 U12618 ( .A(ram[1293]), .B(ram[1309]), .S(n8825), .Z(n3472) );
  MUX2_X1 U12619 ( .A(n3472), .B(n3471), .S(n4247), .Z(n3473) );
  MUX2_X1 U12620 ( .A(n3473), .B(n3470), .S(n4156), .Z(n3474) );
  MUX2_X1 U12621 ( .A(n3474), .B(n3467), .S(n4105), .Z(n3475) );
  MUX2_X1 U12622 ( .A(ram[1261]), .B(ram[1277]), .S(n8825), .Z(n3476) );
  MUX2_X1 U12623 ( .A(ram[1229]), .B(ram[1245]), .S(n8825), .Z(n3477) );
  MUX2_X1 U12624 ( .A(n3477), .B(n3476), .S(n4247), .Z(n3478) );
  MUX2_X1 U12625 ( .A(ram[1197]), .B(ram[1213]), .S(n8825), .Z(n3479) );
  MUX2_X1 U12626 ( .A(ram[1165]), .B(ram[1181]), .S(n8825), .Z(n3480) );
  MUX2_X1 U12627 ( .A(n3480), .B(n3479), .S(n4247), .Z(n3481) );
  MUX2_X1 U12628 ( .A(n3481), .B(n3478), .S(n4156), .Z(n3482) );
  MUX2_X1 U12629 ( .A(ram[1133]), .B(ram[1149]), .S(n8825), .Z(n3483) );
  MUX2_X1 U12630 ( .A(ram[1101]), .B(ram[1117]), .S(n8825), .Z(n3484) );
  MUX2_X1 U12631 ( .A(n3484), .B(n3483), .S(n4247), .Z(n3485) );
  MUX2_X1 U12632 ( .A(ram[1069]), .B(ram[1085]), .S(n8825), .Z(n3486) );
  MUX2_X1 U12633 ( .A(ram[1037]), .B(ram[1053]), .S(n8825), .Z(n3487) );
  MUX2_X1 U12634 ( .A(n3487), .B(n3486), .S(n4247), .Z(n3488) );
  MUX2_X1 U12635 ( .A(n3488), .B(n3485), .S(n4156), .Z(n3489) );
  MUX2_X1 U12636 ( .A(n3489), .B(n3482), .S(n4105), .Z(n3490) );
  MUX2_X1 U12637 ( .A(n3490), .B(n3475), .S(n4085), .Z(n3491) );
  MUX2_X1 U12638 ( .A(n3491), .B(n3460), .S(n4073), .Z(n3492) );
  MUX2_X1 U12639 ( .A(ram[1005]), .B(ram[1021]), .S(n8826), .Z(n3493) );
  MUX2_X1 U12640 ( .A(ram[973]), .B(ram[989]), .S(n8826), .Z(n3494) );
  MUX2_X1 U12641 ( .A(n3494), .B(n3493), .S(n4248), .Z(n3495) );
  MUX2_X1 U12642 ( .A(ram[941]), .B(ram[957]), .S(n8826), .Z(n3496) );
  MUX2_X1 U12643 ( .A(ram[909]), .B(ram[925]), .S(n8826), .Z(n3497) );
  MUX2_X1 U12644 ( .A(n3497), .B(n3496), .S(n4248), .Z(n3498) );
  MUX2_X1 U12645 ( .A(n3498), .B(n3495), .S(n4157), .Z(n3499) );
  MUX2_X1 U12646 ( .A(ram[877]), .B(ram[893]), .S(n8826), .Z(n3500) );
  MUX2_X1 U12647 ( .A(ram[845]), .B(ram[861]), .S(n8826), .Z(n3501) );
  MUX2_X1 U12648 ( .A(n3501), .B(n3500), .S(n4248), .Z(n3502) );
  MUX2_X1 U12649 ( .A(ram[813]), .B(ram[829]), .S(n8826), .Z(n3503) );
  MUX2_X1 U12650 ( .A(ram[781]), .B(ram[797]), .S(n8826), .Z(n3504) );
  MUX2_X1 U12651 ( .A(n3504), .B(n3503), .S(n4248), .Z(n3505) );
  MUX2_X1 U12652 ( .A(n3505), .B(n3502), .S(n4157), .Z(n3506) );
  MUX2_X1 U12653 ( .A(n3506), .B(n3499), .S(n4106), .Z(n3507) );
  MUX2_X1 U12654 ( .A(ram[749]), .B(ram[765]), .S(n8826), .Z(n3508) );
  MUX2_X1 U12655 ( .A(ram[717]), .B(ram[733]), .S(n8826), .Z(n3509) );
  MUX2_X1 U12656 ( .A(n3509), .B(n3508), .S(n4248), .Z(n3510) );
  MUX2_X1 U12657 ( .A(ram[685]), .B(ram[701]), .S(n8826), .Z(n3511) );
  MUX2_X1 U12658 ( .A(ram[653]), .B(ram[669]), .S(n8826), .Z(n3512) );
  MUX2_X1 U12659 ( .A(n3512), .B(n3511), .S(n4248), .Z(n3513) );
  MUX2_X1 U12660 ( .A(n3513), .B(n3510), .S(n4157), .Z(n3514) );
  MUX2_X1 U12661 ( .A(ram[621]), .B(ram[637]), .S(n8827), .Z(n3515) );
  MUX2_X1 U12662 ( .A(ram[589]), .B(ram[605]), .S(n8827), .Z(n3516) );
  MUX2_X1 U12663 ( .A(n3516), .B(n3515), .S(n4248), .Z(n3517) );
  MUX2_X1 U12664 ( .A(ram[557]), .B(ram[573]), .S(n8827), .Z(n3518) );
  MUX2_X1 U12665 ( .A(ram[525]), .B(ram[541]), .S(n8827), .Z(n3519) );
  MUX2_X1 U12666 ( .A(n3519), .B(n3518), .S(n4248), .Z(n3520) );
  MUX2_X1 U12667 ( .A(n3520), .B(n3517), .S(n4157), .Z(n3521) );
  MUX2_X1 U12668 ( .A(n3521), .B(n3514), .S(n4106), .Z(n3522) );
  MUX2_X1 U12669 ( .A(n3522), .B(n3507), .S(n4085), .Z(n3523) );
  MUX2_X1 U12670 ( .A(ram[493]), .B(ram[509]), .S(n8827), .Z(n3524) );
  MUX2_X1 U12671 ( .A(ram[461]), .B(ram[477]), .S(n8827), .Z(n3525) );
  MUX2_X1 U12672 ( .A(n3525), .B(n3524), .S(n4248), .Z(n3526) );
  MUX2_X1 U12673 ( .A(ram[429]), .B(ram[445]), .S(n8827), .Z(n3527) );
  MUX2_X1 U12674 ( .A(ram[397]), .B(ram[413]), .S(n8827), .Z(n3528) );
  MUX2_X1 U12675 ( .A(n3528), .B(n3527), .S(n4248), .Z(n3529) );
  MUX2_X1 U12676 ( .A(n3529), .B(n3526), .S(n4157), .Z(n3530) );
  MUX2_X1 U12677 ( .A(ram[365]), .B(ram[381]), .S(n8827), .Z(n3531) );
  MUX2_X1 U12678 ( .A(ram[333]), .B(ram[349]), .S(n8827), .Z(n3532) );
  MUX2_X1 U12679 ( .A(n3532), .B(n3531), .S(n4248), .Z(n3533) );
  MUX2_X1 U12680 ( .A(ram[301]), .B(ram[317]), .S(n8827), .Z(n3534) );
  MUX2_X1 U12681 ( .A(ram[269]), .B(ram[285]), .S(n8827), .Z(n3535) );
  MUX2_X1 U12682 ( .A(n3535), .B(n3534), .S(n4248), .Z(n3536) );
  MUX2_X1 U12683 ( .A(n3536), .B(n3533), .S(n4157), .Z(n3537) );
  MUX2_X1 U12684 ( .A(n3537), .B(n3530), .S(n4106), .Z(n3538) );
  MUX2_X1 U12685 ( .A(ram[237]), .B(ram[253]), .S(n8828), .Z(n3539) );
  MUX2_X1 U12686 ( .A(ram[205]), .B(ram[221]), .S(n8828), .Z(n3540) );
  MUX2_X1 U12687 ( .A(n3540), .B(n3539), .S(n4249), .Z(n3541) );
  MUX2_X1 U12688 ( .A(ram[173]), .B(ram[189]), .S(n8828), .Z(n3542) );
  MUX2_X1 U12689 ( .A(ram[141]), .B(ram[157]), .S(n8828), .Z(n3543) );
  MUX2_X1 U12690 ( .A(n3543), .B(n3542), .S(n4249), .Z(n3544) );
  MUX2_X1 U12691 ( .A(n3544), .B(n3541), .S(n4157), .Z(n3545) );
  MUX2_X1 U12692 ( .A(ram[109]), .B(ram[125]), .S(n8828), .Z(n3546) );
  MUX2_X1 U12693 ( .A(ram[77]), .B(ram[93]), .S(n8828), .Z(n3547) );
  MUX2_X1 U12694 ( .A(n3547), .B(n3546), .S(n4249), .Z(n3548) );
  MUX2_X1 U12695 ( .A(ram[45]), .B(ram[61]), .S(n8828), .Z(n3549) );
  MUX2_X1 U12696 ( .A(ram[13]), .B(ram[29]), .S(n8828), .Z(n3550) );
  MUX2_X1 U12697 ( .A(n3550), .B(n3549), .S(n4249), .Z(n3551) );
  MUX2_X1 U12698 ( .A(n3551), .B(n3548), .S(n4157), .Z(n3552) );
  MUX2_X1 U12699 ( .A(n3552), .B(n3545), .S(n4106), .Z(n3553) );
  MUX2_X1 U12700 ( .A(n3553), .B(n3538), .S(n4085), .Z(n3554) );
  MUX2_X1 U12701 ( .A(n3554), .B(n3523), .S(n4073), .Z(n3555) );
  MUX2_X1 U12702 ( .A(n3555), .B(n3492), .S(n4067), .Z(n3556) );
  MUX2_X1 U12703 ( .A(n3556), .B(n3429), .S(mem_access_addr[9]), .Z(N288) );
  MUX2_X1 U12704 ( .A(ram[4078]), .B(ram[4094]), .S(n8828), .Z(n3557) );
  MUX2_X1 U12705 ( .A(ram[4046]), .B(ram[4062]), .S(n8828), .Z(n3558) );
  MUX2_X1 U12706 ( .A(n3558), .B(n3557), .S(n4249), .Z(n3559) );
  MUX2_X1 U12707 ( .A(ram[4014]), .B(ram[4030]), .S(n8828), .Z(n3560) );
  MUX2_X1 U12708 ( .A(ram[3982]), .B(ram[3998]), .S(n8828), .Z(n3561) );
  MUX2_X1 U12709 ( .A(n3561), .B(n3560), .S(n4249), .Z(n3562) );
  MUX2_X1 U12710 ( .A(n3562), .B(n3559), .S(n4157), .Z(n3563) );
  MUX2_X1 U12711 ( .A(ram[3950]), .B(ram[3966]), .S(n8829), .Z(n3564) );
  MUX2_X1 U12712 ( .A(ram[3918]), .B(ram[3934]), .S(n8829), .Z(n3565) );
  MUX2_X1 U12713 ( .A(n3565), .B(n3564), .S(n4249), .Z(n3566) );
  MUX2_X1 U12714 ( .A(ram[3886]), .B(ram[3902]), .S(n8829), .Z(n3567) );
  MUX2_X1 U12715 ( .A(ram[3854]), .B(ram[3870]), .S(n8829), .Z(n3568) );
  MUX2_X1 U12716 ( .A(n3568), .B(n3567), .S(n4249), .Z(n3569) );
  MUX2_X1 U12717 ( .A(n3569), .B(n3566), .S(n4157), .Z(n3570) );
  MUX2_X1 U12718 ( .A(n3570), .B(n3563), .S(n4106), .Z(n3571) );
  MUX2_X1 U12719 ( .A(ram[3822]), .B(ram[3838]), .S(n8829), .Z(n3572) );
  MUX2_X1 U12720 ( .A(ram[3790]), .B(ram[3806]), .S(n8829), .Z(n3573) );
  MUX2_X1 U12721 ( .A(n3573), .B(n3572), .S(n4249), .Z(n3574) );
  MUX2_X1 U12722 ( .A(ram[3758]), .B(ram[3774]), .S(n8829), .Z(n3575) );
  MUX2_X1 U12723 ( .A(ram[3726]), .B(ram[3742]), .S(n8829), .Z(n3576) );
  MUX2_X1 U12724 ( .A(n3576), .B(n3575), .S(n4249), .Z(n3577) );
  MUX2_X1 U12725 ( .A(n3577), .B(n3574), .S(n4157), .Z(n3578) );
  MUX2_X1 U12726 ( .A(ram[3694]), .B(ram[3710]), .S(n8829), .Z(n3579) );
  MUX2_X1 U12727 ( .A(ram[3662]), .B(ram[3678]), .S(n8829), .Z(n3580) );
  MUX2_X1 U12728 ( .A(n3580), .B(n3579), .S(n4249), .Z(n3581) );
  MUX2_X1 U12729 ( .A(ram[3630]), .B(ram[3646]), .S(n8829), .Z(n3582) );
  MUX2_X1 U12730 ( .A(ram[3598]), .B(ram[3614]), .S(n8829), .Z(n3583) );
  MUX2_X1 U12731 ( .A(n3583), .B(n3582), .S(n4249), .Z(n3584) );
  MUX2_X1 U12732 ( .A(n3584), .B(n3581), .S(n4157), .Z(n3585) );
  MUX2_X1 U12733 ( .A(n3585), .B(n3578), .S(n4106), .Z(n3586) );
  MUX2_X1 U12734 ( .A(n3586), .B(n3571), .S(n4085), .Z(n3587) );
  MUX2_X1 U12735 ( .A(ram[3566]), .B(ram[3582]), .S(n8830), .Z(n3588) );
  MUX2_X1 U12736 ( .A(ram[3534]), .B(ram[3550]), .S(n8830), .Z(n3589) );
  MUX2_X1 U12737 ( .A(n3589), .B(n3588), .S(n4250), .Z(n3590) );
  MUX2_X1 U12738 ( .A(ram[3502]), .B(ram[3518]), .S(n8830), .Z(n3591) );
  MUX2_X1 U12739 ( .A(ram[3470]), .B(ram[3486]), .S(n8830), .Z(n3592) );
  MUX2_X1 U12740 ( .A(n3592), .B(n3591), .S(n4250), .Z(n3593) );
  MUX2_X1 U12741 ( .A(n3593), .B(n3590), .S(n4158), .Z(n3594) );
  MUX2_X1 U12742 ( .A(ram[3438]), .B(ram[3454]), .S(n8830), .Z(n3595) );
  MUX2_X1 U12743 ( .A(ram[3406]), .B(ram[3422]), .S(n8830), .Z(n3596) );
  MUX2_X1 U12744 ( .A(n3596), .B(n3595), .S(n4250), .Z(n3597) );
  MUX2_X1 U12745 ( .A(ram[3374]), .B(ram[3390]), .S(n8830), .Z(n3598) );
  MUX2_X1 U12746 ( .A(ram[3342]), .B(ram[3358]), .S(n8830), .Z(n3599) );
  MUX2_X1 U12747 ( .A(n3599), .B(n3598), .S(n4250), .Z(n3600) );
  MUX2_X1 U12748 ( .A(n3600), .B(n3597), .S(n4158), .Z(n3601) );
  MUX2_X1 U12749 ( .A(n3601), .B(n3594), .S(n4106), .Z(n3602) );
  MUX2_X1 U12750 ( .A(ram[3310]), .B(ram[3326]), .S(n8830), .Z(n3603) );
  MUX2_X1 U12751 ( .A(ram[3278]), .B(ram[3294]), .S(n8830), .Z(n3604) );
  MUX2_X1 U12752 ( .A(n3604), .B(n3603), .S(n4250), .Z(n3605) );
  MUX2_X1 U12753 ( .A(ram[3246]), .B(ram[3262]), .S(n8830), .Z(n3606) );
  MUX2_X1 U12754 ( .A(ram[3214]), .B(ram[3230]), .S(n8830), .Z(n3607) );
  MUX2_X1 U12755 ( .A(n3607), .B(n3606), .S(n4250), .Z(n3608) );
  MUX2_X1 U12756 ( .A(n3608), .B(n3605), .S(n4158), .Z(n3609) );
  MUX2_X1 U12757 ( .A(ram[3182]), .B(ram[3198]), .S(n8831), .Z(n3610) );
  MUX2_X1 U12758 ( .A(ram[3150]), .B(ram[3166]), .S(n8831), .Z(n3611) );
  MUX2_X1 U12759 ( .A(n3611), .B(n3610), .S(n4250), .Z(n3612) );
  MUX2_X1 U12760 ( .A(ram[3118]), .B(ram[3134]), .S(n8831), .Z(n3613) );
  MUX2_X1 U12761 ( .A(ram[3086]), .B(ram[3102]), .S(n8831), .Z(n3614) );
  MUX2_X1 U12762 ( .A(n3614), .B(n3613), .S(n4250), .Z(n3615) );
  MUX2_X1 U12763 ( .A(n3615), .B(n3612), .S(n4158), .Z(n3616) );
  MUX2_X1 U12764 ( .A(n3616), .B(n3609), .S(n4106), .Z(n3617) );
  MUX2_X1 U12765 ( .A(n3617), .B(n3602), .S(n4085), .Z(n3618) );
  MUX2_X1 U12766 ( .A(n3618), .B(n3587), .S(n4073), .Z(n3619) );
  MUX2_X1 U12767 ( .A(ram[3054]), .B(ram[3070]), .S(n8831), .Z(n3620) );
  MUX2_X1 U12768 ( .A(ram[3022]), .B(ram[3038]), .S(n8831), .Z(n3621) );
  MUX2_X1 U12769 ( .A(n3621), .B(n3620), .S(n4250), .Z(n3622) );
  MUX2_X1 U12770 ( .A(ram[2990]), .B(ram[3006]), .S(n8831), .Z(n3623) );
  MUX2_X1 U12771 ( .A(ram[2958]), .B(ram[2974]), .S(n8831), .Z(n3624) );
  MUX2_X1 U12772 ( .A(n3624), .B(n3623), .S(n4250), .Z(n3625) );
  MUX2_X1 U12773 ( .A(n3625), .B(n3622), .S(n4158), .Z(n3626) );
  MUX2_X1 U12774 ( .A(ram[2926]), .B(ram[2942]), .S(n8831), .Z(n3627) );
  MUX2_X1 U12775 ( .A(ram[2894]), .B(ram[2910]), .S(n8831), .Z(n3628) );
  MUX2_X1 U12776 ( .A(n3628), .B(n3627), .S(n4250), .Z(n3629) );
  MUX2_X1 U12777 ( .A(ram[2862]), .B(ram[2878]), .S(n8831), .Z(n3630) );
  MUX2_X1 U12778 ( .A(ram[2830]), .B(ram[2846]), .S(n8831), .Z(n3631) );
  MUX2_X1 U12779 ( .A(n3631), .B(n3630), .S(n4250), .Z(n3632) );
  MUX2_X1 U12780 ( .A(n3632), .B(n3629), .S(n4158), .Z(n3633) );
  MUX2_X1 U12781 ( .A(n3633), .B(n3626), .S(n4106), .Z(n3634) );
  MUX2_X1 U12782 ( .A(ram[2798]), .B(ram[2814]), .S(n8832), .Z(n3635) );
  MUX2_X1 U12783 ( .A(ram[2766]), .B(ram[2782]), .S(n8832), .Z(n3636) );
  MUX2_X1 U12784 ( .A(n3636), .B(n3635), .S(n4251), .Z(n3637) );
  MUX2_X1 U12785 ( .A(ram[2734]), .B(ram[2750]), .S(n8832), .Z(n3638) );
  MUX2_X1 U12786 ( .A(ram[2702]), .B(ram[2718]), .S(n8832), .Z(n3639) );
  MUX2_X1 U12787 ( .A(n3639), .B(n3638), .S(n4251), .Z(n3640) );
  MUX2_X1 U12788 ( .A(n3640), .B(n3637), .S(n4158), .Z(n3641) );
  MUX2_X1 U12789 ( .A(ram[2670]), .B(ram[2686]), .S(n8832), .Z(n3642) );
  MUX2_X1 U12790 ( .A(ram[2638]), .B(ram[2654]), .S(n8832), .Z(n3643) );
  MUX2_X1 U12791 ( .A(n3643), .B(n3642), .S(n4251), .Z(n3644) );
  MUX2_X1 U12792 ( .A(ram[2606]), .B(ram[2622]), .S(n8832), .Z(n3645) );
  MUX2_X1 U12793 ( .A(ram[2574]), .B(ram[2590]), .S(n8832), .Z(n3646) );
  MUX2_X1 U12794 ( .A(n3646), .B(n3645), .S(n4251), .Z(n3647) );
  MUX2_X1 U12795 ( .A(n3647), .B(n3644), .S(n4158), .Z(n3648) );
  MUX2_X1 U12796 ( .A(n3648), .B(n3641), .S(n4106), .Z(n3649) );
  MUX2_X1 U12797 ( .A(n3649), .B(n3634), .S(n4085), .Z(n3650) );
  MUX2_X1 U12798 ( .A(ram[2542]), .B(ram[2558]), .S(n8832), .Z(n3651) );
  MUX2_X1 U12799 ( .A(ram[2510]), .B(ram[2526]), .S(n8832), .Z(n3652) );
  MUX2_X1 U12800 ( .A(n3652), .B(n3651), .S(n4251), .Z(n3653) );
  MUX2_X1 U12801 ( .A(ram[2478]), .B(ram[2494]), .S(n8832), .Z(n3654) );
  MUX2_X1 U12802 ( .A(ram[2446]), .B(ram[2462]), .S(n8832), .Z(n3655) );
  MUX2_X1 U12803 ( .A(n3655), .B(n3654), .S(n4251), .Z(n3656) );
  MUX2_X1 U12804 ( .A(n3656), .B(n3653), .S(n4158), .Z(n3657) );
  MUX2_X1 U12805 ( .A(ram[2414]), .B(ram[2430]), .S(n8833), .Z(n3658) );
  MUX2_X1 U12806 ( .A(ram[2382]), .B(ram[2398]), .S(n8833), .Z(n3659) );
  MUX2_X1 U12807 ( .A(n3659), .B(n3658), .S(n4251), .Z(n3660) );
  MUX2_X1 U12808 ( .A(ram[2350]), .B(ram[2366]), .S(n8833), .Z(n3661) );
  MUX2_X1 U12809 ( .A(ram[2318]), .B(ram[2334]), .S(n8833), .Z(n3662) );
  MUX2_X1 U12810 ( .A(n3662), .B(n3661), .S(n4251), .Z(n3663) );
  MUX2_X1 U12811 ( .A(n3663), .B(n3660), .S(n4158), .Z(n3664) );
  MUX2_X1 U12812 ( .A(n3664), .B(n3657), .S(n4106), .Z(n3665) );
  MUX2_X1 U12813 ( .A(ram[2286]), .B(ram[2302]), .S(n8833), .Z(n3666) );
  MUX2_X1 U12814 ( .A(ram[2254]), .B(ram[2270]), .S(n8833), .Z(n3667) );
  MUX2_X1 U12815 ( .A(n3667), .B(n3666), .S(n4251), .Z(n3668) );
  MUX2_X1 U12816 ( .A(ram[2222]), .B(ram[2238]), .S(n8833), .Z(n3669) );
  MUX2_X1 U12817 ( .A(ram[2190]), .B(ram[2206]), .S(n8833), .Z(n3670) );
  MUX2_X1 U12818 ( .A(n3670), .B(n3669), .S(n4251), .Z(n3671) );
  MUX2_X1 U12819 ( .A(n3671), .B(n3668), .S(n4158), .Z(n3672) );
  MUX2_X1 U12820 ( .A(ram[2158]), .B(ram[2174]), .S(n8833), .Z(n3673) );
  MUX2_X1 U12821 ( .A(ram[2126]), .B(ram[2142]), .S(n8833), .Z(n3674) );
  MUX2_X1 U12822 ( .A(n3674), .B(n3673), .S(n4251), .Z(n3675) );
  MUX2_X1 U12823 ( .A(ram[2094]), .B(ram[2110]), .S(n8833), .Z(n3676) );
  MUX2_X1 U12824 ( .A(ram[2062]), .B(ram[2078]), .S(n8833), .Z(n3677) );
  MUX2_X1 U12825 ( .A(n3677), .B(n3676), .S(n4251), .Z(n3678) );
  MUX2_X1 U12826 ( .A(n3678), .B(n3675), .S(n4158), .Z(n3679) );
  MUX2_X1 U12827 ( .A(n3679), .B(n3672), .S(n4106), .Z(n3680) );
  MUX2_X1 U12828 ( .A(n3680), .B(n3665), .S(n4085), .Z(n3681) );
  MUX2_X1 U12829 ( .A(n3681), .B(n3650), .S(n4073), .Z(n3682) );
  MUX2_X1 U12830 ( .A(n3682), .B(n3619), .S(n4067), .Z(n3683) );
  MUX2_X1 U12831 ( .A(ram[2030]), .B(ram[2046]), .S(n8834), .Z(n3684) );
  MUX2_X1 U12832 ( .A(ram[1998]), .B(ram[2014]), .S(n8834), .Z(n3685) );
  MUX2_X1 U12833 ( .A(n3685), .B(n3684), .S(n4252), .Z(n3686) );
  MUX2_X1 U12834 ( .A(ram[1966]), .B(ram[1982]), .S(n8834), .Z(n3687) );
  MUX2_X1 U12835 ( .A(ram[1934]), .B(ram[1950]), .S(n8834), .Z(n3688) );
  MUX2_X1 U12836 ( .A(n3688), .B(n3687), .S(n4252), .Z(n3689) );
  MUX2_X1 U12837 ( .A(n3689), .B(n3686), .S(n4159), .Z(n3690) );
  MUX2_X1 U12838 ( .A(ram[1902]), .B(ram[1918]), .S(n8834), .Z(n3691) );
  MUX2_X1 U12839 ( .A(ram[1870]), .B(ram[1886]), .S(n8834), .Z(n3692) );
  MUX2_X1 U12840 ( .A(n3692), .B(n3691), .S(n4252), .Z(n3693) );
  MUX2_X1 U12841 ( .A(ram[1838]), .B(ram[1854]), .S(n8834), .Z(n3694) );
  MUX2_X1 U12842 ( .A(ram[1806]), .B(ram[1822]), .S(n8834), .Z(n3695) );
  MUX2_X1 U12843 ( .A(n3695), .B(n3694), .S(n4252), .Z(n3696) );
  MUX2_X1 U12844 ( .A(n3696), .B(n3693), .S(n4159), .Z(n3697) );
  MUX2_X1 U12845 ( .A(n3697), .B(n3690), .S(n4107), .Z(n3698) );
  MUX2_X1 U12846 ( .A(ram[1774]), .B(ram[1790]), .S(n8834), .Z(n3699) );
  MUX2_X1 U12847 ( .A(ram[1742]), .B(ram[1758]), .S(n8834), .Z(n3700) );
  MUX2_X1 U12848 ( .A(n3700), .B(n3699), .S(n4252), .Z(n3701) );
  MUX2_X1 U12849 ( .A(ram[1710]), .B(ram[1726]), .S(n8834), .Z(n3702) );
  MUX2_X1 U12850 ( .A(ram[1678]), .B(ram[1694]), .S(n8834), .Z(n3703) );
  MUX2_X1 U12851 ( .A(n3703), .B(n3702), .S(n4252), .Z(n3704) );
  MUX2_X1 U12852 ( .A(n3704), .B(n3701), .S(n4159), .Z(n3705) );
  MUX2_X1 U12853 ( .A(ram[1646]), .B(ram[1662]), .S(n8835), .Z(n3706) );
  MUX2_X1 U12854 ( .A(ram[1614]), .B(ram[1630]), .S(n8835), .Z(n3707) );
  MUX2_X1 U12855 ( .A(n3707), .B(n3706), .S(n4252), .Z(n3708) );
  MUX2_X1 U12856 ( .A(ram[1582]), .B(ram[1598]), .S(n8835), .Z(n3709) );
  MUX2_X1 U12857 ( .A(ram[1550]), .B(ram[1566]), .S(n8835), .Z(n3710) );
  MUX2_X1 U12858 ( .A(n3710), .B(n3709), .S(n4252), .Z(n3711) );
  MUX2_X1 U12859 ( .A(n3711), .B(n3708), .S(n4159), .Z(n3712) );
  MUX2_X1 U12860 ( .A(n3712), .B(n3705), .S(n4107), .Z(n3713) );
  MUX2_X1 U12861 ( .A(n3713), .B(n3698), .S(n4086), .Z(n3714) );
  MUX2_X1 U12862 ( .A(ram[1518]), .B(ram[1534]), .S(n8835), .Z(n3715) );
  MUX2_X1 U12863 ( .A(ram[1486]), .B(ram[1502]), .S(n8835), .Z(n3716) );
  MUX2_X1 U12864 ( .A(n3716), .B(n3715), .S(n4252), .Z(n3717) );
  MUX2_X1 U12865 ( .A(ram[1454]), .B(ram[1470]), .S(n8835), .Z(n3718) );
  MUX2_X1 U12866 ( .A(ram[1422]), .B(ram[1438]), .S(n8835), .Z(n3719) );
  MUX2_X1 U12867 ( .A(n3719), .B(n3718), .S(n4252), .Z(n3720) );
  MUX2_X1 U12868 ( .A(n3720), .B(n3717), .S(n4159), .Z(n3721) );
  MUX2_X1 U12869 ( .A(ram[1390]), .B(ram[1406]), .S(n8835), .Z(n3722) );
  MUX2_X1 U12870 ( .A(ram[1358]), .B(ram[1374]), .S(n8835), .Z(n3723) );
  MUX2_X1 U12871 ( .A(n3723), .B(n3722), .S(n4252), .Z(n3724) );
  MUX2_X1 U12872 ( .A(ram[1326]), .B(ram[1342]), .S(n8835), .Z(n3725) );
  MUX2_X1 U12873 ( .A(ram[1294]), .B(ram[1310]), .S(n8835), .Z(n3726) );
  MUX2_X1 U12874 ( .A(n3726), .B(n3725), .S(n4252), .Z(n3727) );
  MUX2_X1 U12875 ( .A(n3727), .B(n3724), .S(n4159), .Z(n3728) );
  MUX2_X1 U12876 ( .A(n3728), .B(n3721), .S(n4107), .Z(n3729) );
  MUX2_X1 U12877 ( .A(ram[1262]), .B(ram[1278]), .S(n8836), .Z(n3730) );
  MUX2_X1 U12878 ( .A(ram[1230]), .B(ram[1246]), .S(n8836), .Z(n3731) );
  MUX2_X1 U12879 ( .A(n3731), .B(n3730), .S(n4253), .Z(n3732) );
  MUX2_X1 U12880 ( .A(ram[1198]), .B(ram[1214]), .S(n8836), .Z(n3733) );
  MUX2_X1 U12881 ( .A(ram[1166]), .B(ram[1182]), .S(n8836), .Z(n3734) );
  MUX2_X1 U12882 ( .A(n3734), .B(n3733), .S(n4253), .Z(n3735) );
  MUX2_X1 U12883 ( .A(n3735), .B(n3732), .S(n4159), .Z(n3736) );
  MUX2_X1 U12884 ( .A(ram[1134]), .B(ram[1150]), .S(n8836), .Z(n3737) );
  MUX2_X1 U12885 ( .A(ram[1102]), .B(ram[1118]), .S(n8836), .Z(n3738) );
  MUX2_X1 U12886 ( .A(n3738), .B(n3737), .S(n4253), .Z(n3739) );
  MUX2_X1 U12887 ( .A(ram[1070]), .B(ram[1086]), .S(n8836), .Z(n3740) );
  MUX2_X1 U12888 ( .A(ram[1038]), .B(ram[1054]), .S(n8836), .Z(n3741) );
  MUX2_X1 U12889 ( .A(n3741), .B(n3740), .S(n4253), .Z(n3742) );
  MUX2_X1 U12890 ( .A(n3742), .B(n3739), .S(n4159), .Z(n3743) );
  MUX2_X1 U12891 ( .A(n3743), .B(n3736), .S(n4107), .Z(n3744) );
  MUX2_X1 U12892 ( .A(n3744), .B(n3729), .S(n4086), .Z(n3745) );
  MUX2_X1 U12893 ( .A(n3745), .B(n3714), .S(n4073), .Z(n3746) );
  MUX2_X1 U12894 ( .A(ram[1006]), .B(ram[1022]), .S(n8836), .Z(n3747) );
  MUX2_X1 U12895 ( .A(ram[974]), .B(ram[990]), .S(n8836), .Z(n3748) );
  MUX2_X1 U12896 ( .A(n3748), .B(n3747), .S(n4253), .Z(n3749) );
  MUX2_X1 U12897 ( .A(ram[942]), .B(ram[958]), .S(n8836), .Z(n3750) );
  MUX2_X1 U12898 ( .A(ram[910]), .B(ram[926]), .S(n8836), .Z(n3751) );
  MUX2_X1 U12899 ( .A(n3751), .B(n3750), .S(n4253), .Z(n3752) );
  MUX2_X1 U12900 ( .A(n3752), .B(n3749), .S(n4159), .Z(n3753) );
  MUX2_X1 U12901 ( .A(ram[878]), .B(ram[894]), .S(n8837), .Z(n3754) );
  MUX2_X1 U12902 ( .A(ram[846]), .B(ram[862]), .S(n8837), .Z(n3755) );
  MUX2_X1 U12903 ( .A(n3755), .B(n3754), .S(n4253), .Z(n3756) );
  MUX2_X1 U12904 ( .A(ram[814]), .B(ram[830]), .S(n8837), .Z(n3757) );
  MUX2_X1 U12905 ( .A(ram[782]), .B(ram[798]), .S(n8837), .Z(n3758) );
  MUX2_X1 U12906 ( .A(n3758), .B(n3757), .S(n4253), .Z(n3759) );
  MUX2_X1 U12907 ( .A(n3759), .B(n3756), .S(n4159), .Z(n3760) );
  MUX2_X1 U12908 ( .A(n3760), .B(n3753), .S(n4107), .Z(n3761) );
  MUX2_X1 U12909 ( .A(ram[750]), .B(ram[766]), .S(n8837), .Z(n3762) );
  MUX2_X1 U12910 ( .A(ram[718]), .B(ram[734]), .S(n8837), .Z(n3763) );
  MUX2_X1 U12911 ( .A(n3763), .B(n3762), .S(n4253), .Z(n3764) );
  MUX2_X1 U12912 ( .A(ram[686]), .B(ram[702]), .S(n8837), .Z(n3765) );
  MUX2_X1 U12913 ( .A(ram[654]), .B(ram[670]), .S(n8837), .Z(n3766) );
  MUX2_X1 U12914 ( .A(n3766), .B(n3765), .S(n4253), .Z(n3767) );
  MUX2_X1 U12915 ( .A(n3767), .B(n3764), .S(n4159), .Z(n3768) );
  MUX2_X1 U12916 ( .A(ram[622]), .B(ram[638]), .S(n8837), .Z(n3769) );
  MUX2_X1 U12917 ( .A(ram[590]), .B(ram[606]), .S(n8837), .Z(n3770) );
  MUX2_X1 U12918 ( .A(n3770), .B(n3769), .S(n4253), .Z(n3771) );
  MUX2_X1 U12919 ( .A(ram[558]), .B(ram[574]), .S(n8837), .Z(n3772) );
  MUX2_X1 U12920 ( .A(ram[526]), .B(ram[542]), .S(n8837), .Z(n3773) );
  MUX2_X1 U12921 ( .A(n3773), .B(n3772), .S(n4253), .Z(n3774) );
  MUX2_X1 U12922 ( .A(n3774), .B(n3771), .S(n4159), .Z(n3775) );
  MUX2_X1 U12923 ( .A(n3775), .B(n3768), .S(n4107), .Z(n3776) );
  MUX2_X1 U12924 ( .A(n3776), .B(n3761), .S(n4086), .Z(n3777) );
  MUX2_X1 U12925 ( .A(ram[494]), .B(ram[510]), .S(n8838), .Z(n3778) );
  MUX2_X1 U12926 ( .A(ram[462]), .B(ram[478]), .S(n8838), .Z(n3779) );
  MUX2_X1 U12927 ( .A(n3779), .B(n3778), .S(n4254), .Z(n3780) );
  MUX2_X1 U12928 ( .A(ram[430]), .B(ram[446]), .S(n8838), .Z(n3781) );
  MUX2_X1 U12929 ( .A(ram[398]), .B(ram[414]), .S(n8838), .Z(n3782) );
  MUX2_X1 U12930 ( .A(n3782), .B(n3781), .S(n4254), .Z(n3783) );
  MUX2_X1 U12931 ( .A(n3783), .B(n3780), .S(n4160), .Z(n3784) );
  MUX2_X1 U12932 ( .A(ram[366]), .B(ram[382]), .S(n8838), .Z(n3785) );
  MUX2_X1 U12933 ( .A(ram[334]), .B(ram[350]), .S(n8838), .Z(n3786) );
  MUX2_X1 U12934 ( .A(n3786), .B(n3785), .S(n4254), .Z(n3787) );
  MUX2_X1 U12935 ( .A(ram[302]), .B(ram[318]), .S(n8838), .Z(n3788) );
  MUX2_X1 U12936 ( .A(ram[270]), .B(ram[286]), .S(n8838), .Z(n3789) );
  MUX2_X1 U12937 ( .A(n3789), .B(n3788), .S(n4254), .Z(n3790) );
  MUX2_X1 U12938 ( .A(n3790), .B(n3787), .S(n4160), .Z(n3791) );
  MUX2_X1 U12939 ( .A(n3791), .B(n3784), .S(n4107), .Z(n3792) );
  MUX2_X1 U12940 ( .A(ram[238]), .B(ram[254]), .S(n8838), .Z(n3793) );
  MUX2_X1 U12941 ( .A(ram[206]), .B(ram[222]), .S(n8838), .Z(n3794) );
  MUX2_X1 U12942 ( .A(n3794), .B(n3793), .S(n4254), .Z(n3795) );
  MUX2_X1 U12943 ( .A(ram[174]), .B(ram[190]), .S(n8838), .Z(n3796) );
  MUX2_X1 U12944 ( .A(ram[142]), .B(ram[158]), .S(n8838), .Z(n3797) );
  MUX2_X1 U12945 ( .A(n3797), .B(n3796), .S(n4254), .Z(n3798) );
  MUX2_X1 U12946 ( .A(n3798), .B(n3795), .S(n4160), .Z(n3799) );
  MUX2_X1 U12947 ( .A(ram[110]), .B(ram[126]), .S(n8839), .Z(n3800) );
  MUX2_X1 U12948 ( .A(ram[78]), .B(ram[94]), .S(n8839), .Z(n3801) );
  MUX2_X1 U12949 ( .A(n3801), .B(n3800), .S(n4254), .Z(n3802) );
  MUX2_X1 U12950 ( .A(ram[46]), .B(ram[62]), .S(n8839), .Z(n3803) );
  MUX2_X1 U12951 ( .A(ram[14]), .B(ram[30]), .S(n8839), .Z(n3804) );
  MUX2_X1 U12952 ( .A(n3804), .B(n3803), .S(n4254), .Z(n3805) );
  MUX2_X1 U12953 ( .A(n3805), .B(n3802), .S(n4160), .Z(n3806) );
  MUX2_X1 U12954 ( .A(n3806), .B(n3799), .S(n4107), .Z(n3807) );
  MUX2_X1 U12955 ( .A(n3807), .B(n3792), .S(n4086), .Z(n3808) );
  MUX2_X1 U12956 ( .A(n3808), .B(n3777), .S(n4073), .Z(n3809) );
  MUX2_X1 U12957 ( .A(n3809), .B(n3746), .S(n4067), .Z(n3810) );
  MUX2_X1 U12958 ( .A(n3810), .B(n3683), .S(mem_access_addr[9]), .Z(N287) );
  MUX2_X1 U12959 ( .A(ram[4079]), .B(ram[4095]), .S(n8839), .Z(n3811) );
  MUX2_X1 U12960 ( .A(ram[4047]), .B(ram[4063]), .S(n8839), .Z(n3812) );
  MUX2_X1 U12961 ( .A(n3812), .B(n3811), .S(n4254), .Z(n3813) );
  MUX2_X1 U12962 ( .A(ram[4015]), .B(ram[4031]), .S(n8839), .Z(n3814) );
  MUX2_X1 U12963 ( .A(ram[3983]), .B(ram[3999]), .S(n8839), .Z(n3815) );
  MUX2_X1 U12964 ( .A(n3815), .B(n3814), .S(n4254), .Z(n3816) );
  MUX2_X1 U12965 ( .A(n3816), .B(n3813), .S(n4160), .Z(n3817) );
  MUX2_X1 U12966 ( .A(ram[3951]), .B(ram[3967]), .S(n8839), .Z(n3818) );
  MUX2_X1 U12967 ( .A(ram[3919]), .B(ram[3935]), .S(n8839), .Z(n3819) );
  MUX2_X1 U12968 ( .A(n3819), .B(n3818), .S(n4254), .Z(n3820) );
  MUX2_X1 U12969 ( .A(ram[3887]), .B(ram[3903]), .S(n8839), .Z(n3821) );
  MUX2_X1 U12970 ( .A(ram[3855]), .B(ram[3871]), .S(n8839), .Z(n3822) );
  MUX2_X1 U12971 ( .A(n3822), .B(n3821), .S(n4254), .Z(n3823) );
  MUX2_X1 U12972 ( .A(n3823), .B(n3820), .S(n4160), .Z(n3824) );
  MUX2_X1 U12973 ( .A(n3824), .B(n3817), .S(n4107), .Z(n3825) );
  MUX2_X1 U12974 ( .A(ram[3823]), .B(ram[3839]), .S(n8840), .Z(n3826) );
  MUX2_X1 U12975 ( .A(ram[3791]), .B(ram[3807]), .S(n8840), .Z(n3827) );
  MUX2_X1 U12976 ( .A(n3827), .B(n3826), .S(n4255), .Z(n3828) );
  MUX2_X1 U12977 ( .A(ram[3759]), .B(ram[3775]), .S(n8840), .Z(n3829) );
  MUX2_X1 U12978 ( .A(ram[3727]), .B(ram[3743]), .S(n8840), .Z(n3830) );
  MUX2_X1 U12979 ( .A(n3830), .B(n3829), .S(n4255), .Z(n3831) );
  MUX2_X1 U12980 ( .A(n3831), .B(n3828), .S(n4160), .Z(n3832) );
  MUX2_X1 U12981 ( .A(ram[3695]), .B(ram[3711]), .S(n8840), .Z(n3833) );
  MUX2_X1 U12982 ( .A(ram[3663]), .B(ram[3679]), .S(n8840), .Z(n3834) );
  MUX2_X1 U12983 ( .A(n3834), .B(n3833), .S(n4255), .Z(n3835) );
  MUX2_X1 U12984 ( .A(ram[3631]), .B(ram[3647]), .S(n8840), .Z(n3836) );
  MUX2_X1 U12985 ( .A(ram[3599]), .B(ram[3615]), .S(n8840), .Z(n3837) );
  MUX2_X1 U12986 ( .A(n3837), .B(n3836), .S(n4255), .Z(n3838) );
  MUX2_X1 U12987 ( .A(n3838), .B(n3835), .S(n4160), .Z(n3839) );
  MUX2_X1 U12988 ( .A(n3839), .B(n3832), .S(n4107), .Z(n3840) );
  MUX2_X1 U12989 ( .A(n3840), .B(n3825), .S(n4086), .Z(n3841) );
  MUX2_X1 U12990 ( .A(ram[3567]), .B(ram[3583]), .S(n8840), .Z(n3842) );
  MUX2_X1 U12991 ( .A(ram[3535]), .B(ram[3551]), .S(n8840), .Z(n3843) );
  MUX2_X1 U12992 ( .A(n3843), .B(n3842), .S(n4255), .Z(n3844) );
  MUX2_X1 U12993 ( .A(ram[3503]), .B(ram[3519]), .S(n8840), .Z(n3845) );
  MUX2_X1 U12994 ( .A(ram[3471]), .B(ram[3487]), .S(n8840), .Z(n3846) );
  MUX2_X1 U12995 ( .A(n3846), .B(n3845), .S(n4255), .Z(n3847) );
  MUX2_X1 U12996 ( .A(n3847), .B(n3844), .S(n4160), .Z(n3848) );
  MUX2_X1 U12997 ( .A(ram[3439]), .B(ram[3455]), .S(n8841), .Z(n3849) );
  MUX2_X1 U12998 ( .A(ram[3407]), .B(ram[3423]), .S(n8841), .Z(n3850) );
  MUX2_X1 U12999 ( .A(n3850), .B(n3849), .S(n4255), .Z(n3851) );
  MUX2_X1 U13000 ( .A(ram[3375]), .B(ram[3391]), .S(n8841), .Z(n3852) );
  MUX2_X1 U13001 ( .A(ram[3343]), .B(ram[3359]), .S(n8841), .Z(n3853) );
  MUX2_X1 U13002 ( .A(n3853), .B(n3852), .S(n4255), .Z(n3854) );
  MUX2_X1 U13003 ( .A(n3854), .B(n3851), .S(n4160), .Z(n3855) );
  MUX2_X1 U13004 ( .A(n3855), .B(n3848), .S(n4107), .Z(n3856) );
  MUX2_X1 U13005 ( .A(ram[3311]), .B(ram[3327]), .S(n8841), .Z(n3857) );
  MUX2_X1 U13006 ( .A(ram[3279]), .B(ram[3295]), .S(n8841), .Z(n3858) );
  MUX2_X1 U13007 ( .A(n3858), .B(n3857), .S(n4255), .Z(n3859) );
  MUX2_X1 U13008 ( .A(ram[3247]), .B(ram[3263]), .S(n8841), .Z(n3860) );
  MUX2_X1 U13009 ( .A(ram[3215]), .B(ram[3231]), .S(n8841), .Z(n3861) );
  MUX2_X1 U13010 ( .A(n3861), .B(n3860), .S(n4255), .Z(n3862) );
  MUX2_X1 U13011 ( .A(n3862), .B(n3859), .S(n4160), .Z(n3863) );
  MUX2_X1 U13012 ( .A(ram[3183]), .B(ram[3199]), .S(n8841), .Z(n3864) );
  MUX2_X1 U13013 ( .A(ram[3151]), .B(ram[3167]), .S(n8841), .Z(n3865) );
  MUX2_X1 U13014 ( .A(n3865), .B(n3864), .S(n4255), .Z(n3866) );
  MUX2_X1 U13015 ( .A(ram[3119]), .B(ram[3135]), .S(n8841), .Z(n3867) );
  MUX2_X1 U13016 ( .A(ram[3087]), .B(ram[3103]), .S(n8841), .Z(n3868) );
  MUX2_X1 U13017 ( .A(n3868), .B(n3867), .S(n4255), .Z(n3869) );
  MUX2_X1 U13018 ( .A(n3869), .B(n3866), .S(n4160), .Z(n3870) );
  MUX2_X1 U13019 ( .A(n3870), .B(n3863), .S(n4107), .Z(n3871) );
  MUX2_X1 U13020 ( .A(n3871), .B(n3856), .S(n4086), .Z(n3872) );
  MUX2_X1 U13021 ( .A(n3872), .B(n3841), .S(n4073), .Z(n3873) );
  MUX2_X1 U13022 ( .A(ram[3055]), .B(ram[3071]), .S(n8842), .Z(n3874) );
  MUX2_X1 U13023 ( .A(ram[3023]), .B(ram[3039]), .S(n8842), .Z(n3875) );
  MUX2_X1 U13024 ( .A(n3875), .B(n3874), .S(n4256), .Z(n3876) );
  MUX2_X1 U13025 ( .A(ram[2991]), .B(ram[3007]), .S(n8842), .Z(n3877) );
  MUX2_X1 U13026 ( .A(ram[2959]), .B(ram[2975]), .S(n8842), .Z(n3878) );
  MUX2_X1 U13027 ( .A(n3878), .B(n3877), .S(n4256), .Z(n3879) );
  MUX2_X1 U13028 ( .A(n3879), .B(n3876), .S(n4161), .Z(n3880) );
  MUX2_X1 U13029 ( .A(ram[2927]), .B(ram[2943]), .S(n8842), .Z(n3881) );
  MUX2_X1 U13030 ( .A(ram[2895]), .B(ram[2911]), .S(n8842), .Z(n3882) );
  MUX2_X1 U13031 ( .A(n3882), .B(n3881), .S(n4256), .Z(n3883) );
  MUX2_X1 U13032 ( .A(ram[2863]), .B(ram[2879]), .S(n8842), .Z(n3884) );
  MUX2_X1 U13033 ( .A(ram[2831]), .B(ram[2847]), .S(n8842), .Z(n3885) );
  MUX2_X1 U13034 ( .A(n3885), .B(n3884), .S(n4256), .Z(n3886) );
  MUX2_X1 U13035 ( .A(n3886), .B(n3883), .S(n4161), .Z(n3887) );
  MUX2_X1 U13036 ( .A(n3887), .B(n3880), .S(n4108), .Z(n3888) );
  MUX2_X1 U13037 ( .A(ram[2799]), .B(ram[2815]), .S(n8842), .Z(n3889) );
  MUX2_X1 U13038 ( .A(ram[2767]), .B(ram[2783]), .S(n8842), .Z(n3890) );
  MUX2_X1 U13039 ( .A(n3890), .B(n3889), .S(n4256), .Z(n3891) );
  MUX2_X1 U13040 ( .A(ram[2735]), .B(ram[2751]), .S(n8842), .Z(n3892) );
  MUX2_X1 U13041 ( .A(ram[2703]), .B(ram[2719]), .S(n8842), .Z(n3893) );
  MUX2_X1 U13042 ( .A(n3893), .B(n3892), .S(n4256), .Z(n3894) );
  MUX2_X1 U13043 ( .A(n3894), .B(n3891), .S(n4161), .Z(n3895) );
  MUX2_X1 U13044 ( .A(ram[2671]), .B(ram[2687]), .S(n8843), .Z(n3896) );
  MUX2_X1 U13045 ( .A(ram[2639]), .B(ram[2655]), .S(n8843), .Z(n3897) );
  MUX2_X1 U13046 ( .A(n3897), .B(n3896), .S(n4256), .Z(n3898) );
  MUX2_X1 U13047 ( .A(ram[2607]), .B(ram[2623]), .S(n8843), .Z(n3899) );
  MUX2_X1 U13048 ( .A(ram[2575]), .B(ram[2591]), .S(n8843), .Z(n3900) );
  MUX2_X1 U13049 ( .A(n3900), .B(n3899), .S(n4256), .Z(n3901) );
  MUX2_X1 U13050 ( .A(n3901), .B(n3898), .S(n4161), .Z(n3902) );
  MUX2_X1 U13051 ( .A(n3902), .B(n3895), .S(n4108), .Z(n3903) );
  MUX2_X1 U13052 ( .A(n3903), .B(n3888), .S(n4086), .Z(n3904) );
  MUX2_X1 U13053 ( .A(ram[2543]), .B(ram[2559]), .S(n8843), .Z(n3905) );
  MUX2_X1 U13054 ( .A(ram[2511]), .B(ram[2527]), .S(n8843), .Z(n3906) );
  MUX2_X1 U13055 ( .A(n3906), .B(n3905), .S(n4256), .Z(n3907) );
  MUX2_X1 U13056 ( .A(ram[2479]), .B(ram[2495]), .S(n8843), .Z(n3908) );
  MUX2_X1 U13057 ( .A(ram[2447]), .B(ram[2463]), .S(n8843), .Z(n3909) );
  MUX2_X1 U13058 ( .A(n3909), .B(n3908), .S(n4256), .Z(n3910) );
  MUX2_X1 U13059 ( .A(n3910), .B(n3907), .S(n4161), .Z(n3911) );
  MUX2_X1 U13060 ( .A(ram[2415]), .B(ram[2431]), .S(n8843), .Z(n3912) );
  MUX2_X1 U13061 ( .A(ram[2383]), .B(ram[2399]), .S(n8843), .Z(n3913) );
  MUX2_X1 U13062 ( .A(n3913), .B(n3912), .S(n4256), .Z(n3914) );
  MUX2_X1 U13063 ( .A(ram[2351]), .B(ram[2367]), .S(n8843), .Z(n3915) );
  MUX2_X1 U13064 ( .A(ram[2319]), .B(ram[2335]), .S(n8843), .Z(n3916) );
  MUX2_X1 U13065 ( .A(n3916), .B(n3915), .S(n4256), .Z(n3917) );
  MUX2_X1 U13066 ( .A(n3917), .B(n3914), .S(n4161), .Z(n3918) );
  MUX2_X1 U13067 ( .A(n3918), .B(n3911), .S(n4108), .Z(n3919) );
  MUX2_X1 U13068 ( .A(ram[2287]), .B(ram[2303]), .S(n8844), .Z(n3920) );
  MUX2_X1 U13069 ( .A(ram[2255]), .B(ram[2271]), .S(n8844), .Z(n3921) );
  MUX2_X1 U13070 ( .A(n3921), .B(n3920), .S(n4257), .Z(n3922) );
  MUX2_X1 U13071 ( .A(ram[2223]), .B(ram[2239]), .S(n8844), .Z(n3923) );
  MUX2_X1 U13072 ( .A(ram[2191]), .B(ram[2207]), .S(n8844), .Z(n3924) );
  MUX2_X1 U13073 ( .A(n3924), .B(n3923), .S(n4257), .Z(n3925) );
  MUX2_X1 U13074 ( .A(n3925), .B(n3922), .S(n4161), .Z(n3926) );
  MUX2_X1 U13075 ( .A(ram[2159]), .B(ram[2175]), .S(n8844), .Z(n3927) );
  MUX2_X1 U13076 ( .A(ram[2127]), .B(ram[2143]), .S(n8844), .Z(n3928) );
  MUX2_X1 U13077 ( .A(n3928), .B(n3927), .S(n4257), .Z(n3929) );
  MUX2_X1 U13078 ( .A(ram[2095]), .B(ram[2111]), .S(n8844), .Z(n3930) );
  MUX2_X1 U13079 ( .A(ram[2063]), .B(ram[2079]), .S(n8844), .Z(n3931) );
  MUX2_X1 U13080 ( .A(n3931), .B(n3930), .S(n4257), .Z(n3932) );
  MUX2_X1 U13081 ( .A(n3932), .B(n3929), .S(n4161), .Z(n3933) );
  MUX2_X1 U13082 ( .A(n3933), .B(n3926), .S(n4108), .Z(n3934) );
  MUX2_X1 U13083 ( .A(n3934), .B(n3919), .S(n4086), .Z(n3935) );
  MUX2_X1 U13084 ( .A(n3935), .B(n3904), .S(n4073), .Z(n3936) );
  MUX2_X1 U13085 ( .A(n3936), .B(n3873), .S(n4067), .Z(n3937) );
  MUX2_X1 U13086 ( .A(ram[2031]), .B(ram[2047]), .S(n8844), .Z(n3938) );
  MUX2_X1 U13087 ( .A(ram[1999]), .B(ram[2015]), .S(n8844), .Z(n3939) );
  MUX2_X1 U13088 ( .A(n3939), .B(n3938), .S(n4257), .Z(n3940) );
  MUX2_X1 U13089 ( .A(ram[1967]), .B(ram[1983]), .S(n8844), .Z(n3941) );
  MUX2_X1 U13090 ( .A(ram[1935]), .B(ram[1951]), .S(n8844), .Z(n3942) );
  MUX2_X1 U13091 ( .A(n3942), .B(n3941), .S(n4257), .Z(n3943) );
  MUX2_X1 U13092 ( .A(n3943), .B(n3940), .S(n4161), .Z(n3944) );
  MUX2_X1 U13093 ( .A(ram[1903]), .B(ram[1919]), .S(n8845), .Z(n3945) );
  MUX2_X1 U13094 ( .A(ram[1871]), .B(ram[1887]), .S(n8845), .Z(n3946) );
  MUX2_X1 U13095 ( .A(n3946), .B(n3945), .S(n4257), .Z(n3947) );
  MUX2_X1 U13096 ( .A(ram[1839]), .B(ram[1855]), .S(n8845), .Z(n3948) );
  MUX2_X1 U13097 ( .A(ram[1807]), .B(ram[1823]), .S(n8845), .Z(n3949) );
  MUX2_X1 U13098 ( .A(n3949), .B(n3948), .S(n4257), .Z(n3950) );
  MUX2_X1 U13099 ( .A(n3950), .B(n3947), .S(n4161), .Z(n3951) );
  MUX2_X1 U13100 ( .A(n3951), .B(n3944), .S(n4108), .Z(n3952) );
  MUX2_X1 U13101 ( .A(ram[1775]), .B(ram[1791]), .S(n8845), .Z(n3953) );
  MUX2_X1 U13102 ( .A(ram[1743]), .B(ram[1759]), .S(n8845), .Z(n3954) );
  MUX2_X1 U13103 ( .A(n3954), .B(n3953), .S(n4257), .Z(n3955) );
  MUX2_X1 U13104 ( .A(ram[1711]), .B(ram[1727]), .S(n8845), .Z(n3956) );
  MUX2_X1 U13105 ( .A(ram[1679]), .B(ram[1695]), .S(n8845), .Z(n3957) );
  MUX2_X1 U13106 ( .A(n3957), .B(n3956), .S(n4257), .Z(n3958) );
  MUX2_X1 U13107 ( .A(n3958), .B(n3955), .S(n4161), .Z(n3959) );
  MUX2_X1 U13108 ( .A(ram[1647]), .B(ram[1663]), .S(n8845), .Z(n3960) );
  MUX2_X1 U13109 ( .A(ram[1615]), .B(ram[1631]), .S(n8845), .Z(n3961) );
  MUX2_X1 U13110 ( .A(n3961), .B(n3960), .S(n4257), .Z(n3962) );
  MUX2_X1 U13111 ( .A(ram[1583]), .B(ram[1599]), .S(n8845), .Z(n3963) );
  MUX2_X1 U13112 ( .A(ram[1551]), .B(ram[1567]), .S(n8845), .Z(n3964) );
  MUX2_X1 U13113 ( .A(n3964), .B(n3963), .S(n4257), .Z(n3965) );
  MUX2_X1 U13114 ( .A(n3965), .B(n3962), .S(n4161), .Z(n3966) );
  MUX2_X1 U13115 ( .A(n3966), .B(n3959), .S(n4108), .Z(n3967) );
  MUX2_X1 U13116 ( .A(n3967), .B(n3952), .S(n4086), .Z(n3968) );
  MUX2_X1 U13117 ( .A(ram[1519]), .B(ram[1535]), .S(n8846), .Z(n3969) );
  MUX2_X1 U13118 ( .A(ram[1487]), .B(ram[1503]), .S(n8846), .Z(n3970) );
  MUX2_X1 U13119 ( .A(n3970), .B(n3969), .S(n4258), .Z(n3971) );
  MUX2_X1 U13120 ( .A(ram[1455]), .B(ram[1471]), .S(n8846), .Z(n3972) );
  MUX2_X1 U13121 ( .A(ram[1423]), .B(ram[1439]), .S(n8846), .Z(n3973) );
  MUX2_X1 U13122 ( .A(n3973), .B(n3972), .S(n4258), .Z(n3974) );
  MUX2_X1 U13123 ( .A(n3974), .B(n3971), .S(n4162), .Z(n3975) );
  MUX2_X1 U13124 ( .A(ram[1391]), .B(ram[1407]), .S(n8846), .Z(n3976) );
  MUX2_X1 U13125 ( .A(ram[1359]), .B(ram[1375]), .S(n8846), .Z(n3977) );
  MUX2_X1 U13126 ( .A(n3977), .B(n3976), .S(n4258), .Z(n3978) );
  MUX2_X1 U13127 ( .A(ram[1327]), .B(ram[1343]), .S(n8846), .Z(n3979) );
  MUX2_X1 U13128 ( .A(ram[1295]), .B(ram[1311]), .S(n8846), .Z(n3980) );
  MUX2_X1 U13129 ( .A(n3980), .B(n3979), .S(n4258), .Z(n3981) );
  MUX2_X1 U13130 ( .A(n3981), .B(n3978), .S(n4162), .Z(n3982) );
  MUX2_X1 U13131 ( .A(n3982), .B(n3975), .S(n4108), .Z(n3983) );
  MUX2_X1 U13132 ( .A(ram[1263]), .B(ram[1279]), .S(n8846), .Z(n3984) );
  MUX2_X1 U13133 ( .A(ram[1231]), .B(ram[1247]), .S(n8846), .Z(n3985) );
  MUX2_X1 U13134 ( .A(n3985), .B(n3984), .S(n4258), .Z(n3986) );
  MUX2_X1 U13135 ( .A(ram[1199]), .B(ram[1215]), .S(n8846), .Z(n3987) );
  MUX2_X1 U13136 ( .A(ram[1167]), .B(ram[1183]), .S(n8846), .Z(n3988) );
  MUX2_X1 U13137 ( .A(n3988), .B(n3987), .S(n4258), .Z(n3989) );
  MUX2_X1 U13138 ( .A(n3989), .B(n3986), .S(n4162), .Z(n3990) );
  MUX2_X1 U13139 ( .A(ram[1135]), .B(ram[1151]), .S(n8847), .Z(n3991) );
  MUX2_X1 U13140 ( .A(ram[1103]), .B(ram[1119]), .S(n8847), .Z(n3992) );
  MUX2_X1 U13141 ( .A(n3992), .B(n3991), .S(n4258), .Z(n3993) );
  MUX2_X1 U13142 ( .A(ram[1071]), .B(ram[1087]), .S(n8847), .Z(n3994) );
  MUX2_X1 U13143 ( .A(ram[1039]), .B(ram[1055]), .S(n8847), .Z(n3995) );
  MUX2_X1 U13144 ( .A(n3995), .B(n3994), .S(n4258), .Z(n3996) );
  MUX2_X1 U13145 ( .A(n3996), .B(n3993), .S(n4162), .Z(n3997) );
  MUX2_X1 U13146 ( .A(n3997), .B(n3990), .S(n4108), .Z(n3998) );
  MUX2_X1 U13147 ( .A(n3998), .B(n3983), .S(n4086), .Z(n3999) );
  MUX2_X1 U13148 ( .A(n3999), .B(n3968), .S(n4073), .Z(n4000) );
  MUX2_X1 U13149 ( .A(ram[1007]), .B(ram[1023]), .S(n8847), .Z(n4001) );
  MUX2_X1 U13150 ( .A(ram[975]), .B(ram[991]), .S(n8847), .Z(n4002) );
  MUX2_X1 U13151 ( .A(n4002), .B(n4001), .S(n4258), .Z(n4003) );
  MUX2_X1 U13152 ( .A(ram[943]), .B(ram[959]), .S(n8847), .Z(n4004) );
  MUX2_X1 U13153 ( .A(ram[911]), .B(ram[927]), .S(n8847), .Z(n4005) );
  MUX2_X1 U13154 ( .A(n4005), .B(n4004), .S(n4258), .Z(n4006) );
  MUX2_X1 U13155 ( .A(n4006), .B(n4003), .S(n4162), .Z(n4007) );
  MUX2_X1 U13156 ( .A(ram[879]), .B(ram[895]), .S(n8847), .Z(n4008) );
  MUX2_X1 U13157 ( .A(ram[847]), .B(ram[863]), .S(n8847), .Z(n4009) );
  MUX2_X1 U13158 ( .A(n4009), .B(n4008), .S(n4258), .Z(n4010) );
  MUX2_X1 U13159 ( .A(ram[815]), .B(ram[831]), .S(n8847), .Z(n4011) );
  MUX2_X1 U13160 ( .A(ram[783]), .B(ram[799]), .S(n8847), .Z(n4012) );
  MUX2_X1 U13161 ( .A(n4012), .B(n4011), .S(n4258), .Z(n4013) );
  MUX2_X1 U13162 ( .A(n4013), .B(n4010), .S(n4162), .Z(n4014) );
  MUX2_X1 U13163 ( .A(n4014), .B(n4007), .S(n4108), .Z(n4015) );
  MUX2_X1 U13164 ( .A(ram[751]), .B(ram[767]), .S(n8848), .Z(n4016) );
  MUX2_X1 U13165 ( .A(ram[719]), .B(ram[735]), .S(n8848), .Z(n4017) );
  MUX2_X1 U13166 ( .A(n4017), .B(n4016), .S(n4259), .Z(n4018) );
  MUX2_X1 U13167 ( .A(ram[687]), .B(ram[703]), .S(n8848), .Z(n4019) );
  MUX2_X1 U13168 ( .A(ram[655]), .B(ram[671]), .S(n8848), .Z(n4020) );
  MUX2_X1 U13169 ( .A(n4020), .B(n4019), .S(n4259), .Z(n4021) );
  MUX2_X1 U13170 ( .A(n4021), .B(n4018), .S(n4162), .Z(n4022) );
  MUX2_X1 U13171 ( .A(ram[623]), .B(ram[639]), .S(n8848), .Z(n4023) );
  MUX2_X1 U13172 ( .A(ram[591]), .B(ram[607]), .S(n8848), .Z(n4024) );
  MUX2_X1 U13173 ( .A(n4024), .B(n4023), .S(n4259), .Z(n4025) );
  MUX2_X1 U13174 ( .A(ram[559]), .B(ram[575]), .S(n8848), .Z(n4026) );
  MUX2_X1 U13175 ( .A(ram[527]), .B(ram[543]), .S(n8848), .Z(n4027) );
  MUX2_X1 U13176 ( .A(n4027), .B(n4026), .S(n4259), .Z(n4028) );
  MUX2_X1 U13177 ( .A(n4028), .B(n4025), .S(n4162), .Z(n4029) );
  MUX2_X1 U13178 ( .A(n4029), .B(n4022), .S(n4108), .Z(n4030) );
  MUX2_X1 U13179 ( .A(n4030), .B(n4015), .S(n4086), .Z(n4031) );
  MUX2_X1 U13180 ( .A(ram[495]), .B(ram[511]), .S(n8848), .Z(n4032) );
  MUX2_X1 U13181 ( .A(ram[463]), .B(ram[479]), .S(n8848), .Z(n4033) );
  MUX2_X1 U13182 ( .A(n4033), .B(n4032), .S(n4259), .Z(n4034) );
  MUX2_X1 U13183 ( .A(ram[431]), .B(ram[447]), .S(n8848), .Z(n4035) );
  MUX2_X1 U13184 ( .A(ram[399]), .B(ram[415]), .S(n8848), .Z(n4036) );
  MUX2_X1 U13185 ( .A(n4036), .B(n4035), .S(n4259), .Z(n4037) );
  MUX2_X1 U13186 ( .A(n4037), .B(n4034), .S(n4162), .Z(n4038) );
  MUX2_X1 U13187 ( .A(ram[367]), .B(ram[383]), .S(n8849), .Z(n4039) );
  MUX2_X1 U13188 ( .A(ram[335]), .B(ram[351]), .S(n8849), .Z(n4040) );
  MUX2_X1 U13189 ( .A(n4040), .B(n4039), .S(n4259), .Z(n4041) );
  MUX2_X1 U13190 ( .A(ram[303]), .B(ram[319]), .S(n8849), .Z(n4042) );
  MUX2_X1 U13191 ( .A(ram[271]), .B(ram[287]), .S(n8849), .Z(n4043) );
  MUX2_X1 U13192 ( .A(n4043), .B(n4042), .S(n4259), .Z(n4044) );
  MUX2_X1 U13193 ( .A(n4044), .B(n4041), .S(n4162), .Z(n4045) );
  MUX2_X1 U13194 ( .A(n4045), .B(n4038), .S(n4108), .Z(n4046) );
  MUX2_X1 U13195 ( .A(ram[239]), .B(ram[255]), .S(n8849), .Z(n4047) );
  MUX2_X1 U13196 ( .A(ram[207]), .B(ram[223]), .S(n8849), .Z(n4048) );
  MUX2_X1 U13197 ( .A(n4048), .B(n4047), .S(n4259), .Z(n4049) );
  MUX2_X1 U13198 ( .A(ram[175]), .B(ram[191]), .S(n8849), .Z(n4050) );
  MUX2_X1 U13199 ( .A(ram[143]), .B(ram[159]), .S(n8849), .Z(n4051) );
  MUX2_X1 U13200 ( .A(n4051), .B(n4050), .S(n4259), .Z(n4052) );
  MUX2_X1 U13201 ( .A(n4052), .B(n4049), .S(n4162), .Z(n4053) );
  MUX2_X1 U13202 ( .A(ram[111]), .B(ram[127]), .S(n8849), .Z(n4054) );
  MUX2_X1 U13203 ( .A(ram[79]), .B(ram[95]), .S(n8849), .Z(n4055) );
  MUX2_X1 U13204 ( .A(n4055), .B(n4054), .S(n4259), .Z(n4056) );
  MUX2_X1 U13205 ( .A(ram[47]), .B(ram[63]), .S(n8849), .Z(n4057) );
  MUX2_X1 U13206 ( .A(ram[15]), .B(ram[31]), .S(n8849), .Z(n4058) );
  MUX2_X1 U13207 ( .A(n4058), .B(n4057), .S(n4259), .Z(n4059) );
  MUX2_X1 U13208 ( .A(n4059), .B(n4056), .S(n4162), .Z(n4060) );
  MUX2_X1 U13209 ( .A(n4060), .B(n4053), .S(n4108), .Z(n4061) );
  MUX2_X1 U13210 ( .A(n4061), .B(n4046), .S(n4086), .Z(n4062) );
  MUX2_X1 U13211 ( .A(n4062), .B(n4031), .S(n4073), .Z(n4063) );
  MUX2_X1 U13212 ( .A(n4063), .B(n4000), .S(n4067), .Z(n4064) );
  MUX2_X1 U13213 ( .A(n4064), .B(n3937), .S(mem_access_addr[9]), .Z(N286) );
  BUF_X1 U13214 ( .A(n4074), .Z(n4068) );
  BUF_X1 U13215 ( .A(mem_access_addr[7]), .Z(n4074) );
  BUF_X1 U13216 ( .A(mem_access_addr[7]), .Z(n4075) );
  BUF_X1 U13217 ( .A(n9238), .Z(n4076) );
  BUF_X1 U13218 ( .A(n9238), .Z(n4081) );
  BUF_X1 U13219 ( .A(n9238), .Z(n4082) );
  BUF_X1 U13220 ( .A(n9238), .Z(n4083) );
  BUF_X1 U13221 ( .A(n9238), .Z(n4084) );
  BUF_X1 U13222 ( .A(n9238), .Z(n4085) );
  BUF_X1 U13223 ( .A(n9238), .Z(n4086) );
  BUF_X1 U13224 ( .A(n4109), .Z(n4087) );
  BUF_X1 U13225 ( .A(n4109), .Z(n4092) );
  BUF_X1 U13226 ( .A(n4109), .Z(n4093) );
  BUF_X1 U13227 ( .A(n4109), .Z(n4094) );
  BUF_X1 U13228 ( .A(n4109), .Z(n4095) );
  BUF_X1 U13229 ( .A(n4109), .Z(n4096) );
  BUF_X1 U13230 ( .A(n4109), .Z(n4097) );
  BUF_X1 U13231 ( .A(n4110), .Z(n4102) );
  BUF_X1 U13232 ( .A(n4110), .Z(n4103) );
  BUF_X1 U13233 ( .A(n4110), .Z(n4104) );
  BUF_X1 U13234 ( .A(n4110), .Z(n4105) );
  BUF_X1 U13235 ( .A(n4110), .Z(n4106) );
  BUF_X1 U13236 ( .A(n4110), .Z(n4107) );
  BUF_X1 U13237 ( .A(n4110), .Z(n4108) );
  BUF_X1 U13238 ( .A(n4119), .Z(n4120) );
  BUF_X1 U13239 ( .A(n4173), .Z(n4174) );
  BUF_X1 U13240 ( .A(n4173), .Z(n4179) );
  BUF_X1 U13241 ( .A(n4173), .Z(n4180) );
  BUF_X1 U13242 ( .A(n4173), .Z(n4181) );
  BUF_X1 U13243 ( .A(n4173), .Z(n4182) );
  BUF_X1 U13244 ( .A(n4173), .Z(n4183) );
  BUF_X1 U13245 ( .A(n4173), .Z(n4184) );
  BUF_X1 U13246 ( .A(n4172), .Z(n4189) );
  BUF_X1 U13247 ( .A(n4172), .Z(n4190) );
  BUF_X1 U13248 ( .A(n4172), .Z(n4191) );
  BUF_X1 U13249 ( .A(n4172), .Z(n4192) );
  BUF_X1 U13250 ( .A(n4172), .Z(n4193) );
  BUF_X1 U13251 ( .A(n4172), .Z(n4194) );
  BUF_X1 U13252 ( .A(n4172), .Z(n4195) );
  BUF_X1 U13253 ( .A(n4171), .Z(n4200) );
  BUF_X1 U13254 ( .A(n4171), .Z(n4201) );
  BUF_X1 U13255 ( .A(n4171), .Z(n4202) );
  BUF_X1 U13256 ( .A(n4171), .Z(n4203) );
  BUF_X1 U13257 ( .A(n4171), .Z(n4204) );
  BUF_X1 U13258 ( .A(n4171), .Z(n4205) );
  BUF_X1 U13259 ( .A(n4171), .Z(n4206) );
  BUF_X1 U13260 ( .A(n4170), .Z(n4211) );
  BUF_X1 U13261 ( .A(n4170), .Z(n4212) );
  BUF_X1 U13262 ( .A(n4170), .Z(n4213) );
  BUF_X1 U13263 ( .A(n4170), .Z(n4214) );
  BUF_X1 U13264 ( .A(n4170), .Z(n4215) );
  BUF_X1 U13265 ( .A(n4170), .Z(n4216) );
  BUF_X1 U13266 ( .A(n4170), .Z(n4217) );
  BUF_X1 U13267 ( .A(n4169), .Z(n4222) );
  BUF_X1 U13268 ( .A(n4169), .Z(n4223) );
  BUF_X1 U13269 ( .A(n4169), .Z(n4224) );
  BUF_X1 U13270 ( .A(n4169), .Z(n4225) );
  BUF_X1 U13271 ( .A(n4169), .Z(n4226) );
  BUF_X1 U13272 ( .A(n4169), .Z(n4227) );
  BUF_X1 U13273 ( .A(n4169), .Z(n4228) );
  BUF_X1 U13274 ( .A(n4168), .Z(n4233) );
  BUF_X1 U13275 ( .A(n4168), .Z(n4234) );
  BUF_X1 U13276 ( .A(n4168), .Z(n4235) );
  BUF_X1 U13277 ( .A(n4168), .Z(n4236) );
  BUF_X1 U13278 ( .A(n4168), .Z(n4237) );
  BUF_X1 U13279 ( .A(n4168), .Z(n4238) );
  BUF_X1 U13280 ( .A(n4168), .Z(n4239) );
  BUF_X1 U13281 ( .A(n4167), .Z(n4244) );
  BUF_X1 U13282 ( .A(n4167), .Z(n4245) );
  BUF_X1 U13283 ( .A(n4167), .Z(n4246) );
  BUF_X1 U13284 ( .A(n4167), .Z(n4247) );
  BUF_X1 U13285 ( .A(n4167), .Z(n4248) );
  BUF_X1 U13286 ( .A(n4167), .Z(n4249) );
  BUF_X1 U13287 ( .A(n4167), .Z(n4250) );
  BUF_X1 U13288 ( .A(n4166), .Z(n4255) );
  BUF_X1 U13289 ( .A(n4166), .Z(n4256) );
  BUF_X1 U13290 ( .A(n4166), .Z(n4257) );
  BUF_X1 U13291 ( .A(n4166), .Z(n4258) );
  BUF_X1 U13292 ( .A(n4166), .Z(n4259) );
  BUF_X1 U13293 ( .A(n4278), .Z(n4279) );
  BUF_X1 U13294 ( .A(n4278), .Z(n4284) );
  BUF_X1 U13295 ( .A(n4278), .Z(n4285) );
  BUF_X1 U13296 ( .A(n4278), .Z(n4286) );
  BUF_X1 U13297 ( .A(n4278), .Z(n4287) );
  BUF_X1 U13298 ( .A(n4278), .Z(n4288) );
  BUF_X1 U13299 ( .A(n4278), .Z(n4289) );
  BUF_X1 U13300 ( .A(n4277), .Z(n4294) );
  BUF_X1 U13301 ( .A(n4277), .Z(n4295) );
  BUF_X1 U13302 ( .A(n4277), .Z(n4296) );
  BUF_X1 U13303 ( .A(n4277), .Z(n4297) );
  BUF_X1 U13304 ( .A(n4277), .Z(n4298) );
  BUF_X1 U13305 ( .A(n4277), .Z(n4299) );
  BUF_X1 U13306 ( .A(n4277), .Z(n4300) );
  BUF_X1 U13307 ( .A(n4276), .Z(n4305) );
  BUF_X1 U13308 ( .A(n4276), .Z(n4306) );
  BUF_X1 U13309 ( .A(n4276), .Z(n4307) );
  BUF_X1 U13310 ( .A(n4276), .Z(n4308) );
  BUF_X1 U13311 ( .A(n4276), .Z(n4309) );
  BUF_X1 U13312 ( .A(n4276), .Z(n4310) );
  BUF_X1 U13313 ( .A(n4276), .Z(n4311) );
  BUF_X1 U13314 ( .A(n4275), .Z(n4316) );
  BUF_X1 U13315 ( .A(n4275), .Z(n4317) );
  BUF_X1 U13316 ( .A(n4275), .Z(n4318) );
  BUF_X1 U13317 ( .A(n4275), .Z(n4319) );
  BUF_X1 U13318 ( .A(n4275), .Z(n4320) );
  BUF_X1 U13319 ( .A(n4275), .Z(n4321) );
  BUF_X1 U13320 ( .A(n4275), .Z(n4322) );
  BUF_X1 U13321 ( .A(n4274), .Z(n4327) );
  BUF_X1 U13322 ( .A(n4274), .Z(n4328) );
  BUF_X1 U13323 ( .A(n4274), .Z(n4329) );
  BUF_X1 U13324 ( .A(n4274), .Z(n4330) );
  BUF_X1 U13325 ( .A(n4274), .Z(n4331) );
  BUF_X1 U13326 ( .A(n4274), .Z(n4332) );
  BUF_X1 U13327 ( .A(n4274), .Z(n4333) );
  BUF_X1 U13328 ( .A(n4273), .Z(n4338) );
  BUF_X1 U13329 ( .A(n4273), .Z(n4339) );
  BUF_X1 U13330 ( .A(n4273), .Z(n4340) );
  BUF_X1 U13331 ( .A(n4273), .Z(n4341) );
  BUF_X1 U13332 ( .A(n4273), .Z(n4342) );
  BUF_X1 U13333 ( .A(n4273), .Z(n4343) );
  BUF_X1 U13334 ( .A(n4273), .Z(n4344) );
  BUF_X1 U13335 ( .A(n4272), .Z(n4349) );
  BUF_X1 U13336 ( .A(n4272), .Z(n4350) );
  BUF_X1 U13337 ( .A(n4272), .Z(n4351) );
  BUF_X1 U13338 ( .A(n4272), .Z(n4352) );
  BUF_X1 U13339 ( .A(n4272), .Z(n4353) );
  BUF_X1 U13340 ( .A(n4272), .Z(n4354) );
  BUF_X1 U13341 ( .A(n4272), .Z(n4355) );
  BUF_X1 U13342 ( .A(n4271), .Z(n8760) );
  BUF_X1 U13343 ( .A(n4271), .Z(n8761) );
  BUF_X1 U13344 ( .A(n4271), .Z(n8762) );
  BUF_X1 U13345 ( .A(n4271), .Z(n8763) );
  BUF_X1 U13346 ( .A(n4271), .Z(n8764) );
  BUF_X1 U13347 ( .A(n4271), .Z(n8765) );
  BUF_X1 U13348 ( .A(n4271), .Z(n8766) );
  BUF_X1 U13349 ( .A(n4270), .Z(n8771) );
  BUF_X1 U13350 ( .A(n4270), .Z(n8772) );
  BUF_X1 U13351 ( .A(n4270), .Z(n8773) );
  BUF_X1 U13352 ( .A(n4270), .Z(n8774) );
  BUF_X1 U13353 ( .A(n4270), .Z(n8775) );
  BUF_X1 U13354 ( .A(n4270), .Z(n8776) );
  BUF_X1 U13355 ( .A(n4270), .Z(n8777) );
  BUF_X1 U13356 ( .A(n4269), .Z(n8782) );
  BUF_X1 U13357 ( .A(n4269), .Z(n8783) );
  BUF_X1 U13358 ( .A(n4269), .Z(n8784) );
  BUF_X1 U13359 ( .A(n4269), .Z(n8785) );
  BUF_X1 U13360 ( .A(n4269), .Z(n8786) );
  BUF_X1 U13361 ( .A(n4269), .Z(n8787) );
  BUF_X1 U13362 ( .A(n4269), .Z(n8788) );
  BUF_X1 U13363 ( .A(n4268), .Z(n8793) );
  BUF_X1 U13364 ( .A(n4268), .Z(n8794) );
  BUF_X1 U13365 ( .A(n4268), .Z(n8795) );
  BUF_X1 U13366 ( .A(n4268), .Z(n8796) );
  BUF_X1 U13367 ( .A(n4268), .Z(n8797) );
  BUF_X1 U13368 ( .A(n4268), .Z(n8798) );
  BUF_X1 U13369 ( .A(n4268), .Z(n8799) );
  BUF_X1 U13370 ( .A(n4267), .Z(n8804) );
  BUF_X1 U13371 ( .A(n4267), .Z(n8805) );
  BUF_X1 U13372 ( .A(n4267), .Z(n8806) );
  BUF_X1 U13373 ( .A(n4267), .Z(n8807) );
  BUF_X1 U13374 ( .A(n4267), .Z(n8808) );
  BUF_X1 U13375 ( .A(n4267), .Z(n8809) );
  BUF_X1 U13376 ( .A(n4267), .Z(n8810) );
  BUF_X1 U13377 ( .A(n4266), .Z(n8815) );
  BUF_X1 U13378 ( .A(n4266), .Z(n8816) );
  BUF_X1 U13379 ( .A(n4266), .Z(n8817) );
  BUF_X1 U13380 ( .A(n4266), .Z(n8818) );
  BUF_X1 U13381 ( .A(n4266), .Z(n8819) );
  BUF_X1 U13382 ( .A(n4266), .Z(n8820) );
  BUF_X1 U13383 ( .A(n4266), .Z(n8821) );
  BUF_X1 U13384 ( .A(n4265), .Z(n8826) );
  BUF_X1 U13385 ( .A(n4265), .Z(n8827) );
  BUF_X1 U13386 ( .A(n4265), .Z(n8828) );
  BUF_X1 U13387 ( .A(n4265), .Z(n8829) );
  BUF_X1 U13388 ( .A(n4265), .Z(n8830) );
  BUF_X1 U13389 ( .A(n4265), .Z(n8831) );
  BUF_X1 U13390 ( .A(n4265), .Z(n8832) );
  BUF_X1 U13391 ( .A(n4264), .Z(n8837) );
  BUF_X1 U13392 ( .A(n4264), .Z(n8838) );
  BUF_X1 U13393 ( .A(n4264), .Z(n8839) );
  BUF_X1 U13394 ( .A(n4264), .Z(n8840) );
  BUF_X1 U13395 ( .A(n4264), .Z(n8841) );
  BUF_X1 U13396 ( .A(n4264), .Z(n8842) );
  BUF_X1 U13397 ( .A(n4264), .Z(n8843) );
  BUF_X1 U13398 ( .A(n8852), .Z(n8854) );
  BUF_X1 U13399 ( .A(n8852), .Z(n8855) );
  BUF_X1 U13400 ( .A(n8852), .Z(n8856) );
  BUF_X1 U13401 ( .A(n8852), .Z(n8857) );
  BUF_X1 U13402 ( .A(n8852), .Z(n8858) );
  BUF_X1 U13403 ( .A(n8852), .Z(n8859) );
  BUF_X1 U13404 ( .A(n8852), .Z(n8860) );
  BUF_X1 U13405 ( .A(n8853), .Z(n8865) );
  BUF_X1 U13406 ( .A(n8853), .Z(n8866) );
  BUF_X1 U13407 ( .A(n8853), .Z(n8867) );
  BUF_X1 U13408 ( .A(n8853), .Z(n8868) );
  BUF_X1 U13409 ( .A(n8853), .Z(n8869) );
  BUF_X1 U13410 ( .A(n8853), .Z(n8870) );
  BUF_X1 U13411 ( .A(n8853), .Z(n8875) );
  BUF_X1 U13412 ( .A(n8876), .Z(n8878) );
  BUF_X1 U13413 ( .A(n8876), .Z(n8879) );
  BUF_X1 U13414 ( .A(n8876), .Z(n8880) );
  BUF_X1 U13415 ( .A(n8876), .Z(n8881) );
  BUF_X1 U13416 ( .A(n8876), .Z(n8882) );
  BUF_X1 U13417 ( .A(n8876), .Z(n8883) );
  BUF_X1 U13418 ( .A(n8876), .Z(n8884) );
  BUF_X1 U13419 ( .A(n8877), .Z(n8889) );
  BUF_X1 U13420 ( .A(n8877), .Z(n8890) );
  BUF_X1 U13421 ( .A(n8877), .Z(n8891) );
  BUF_X1 U13422 ( .A(n8877), .Z(n8892) );
  BUF_X1 U13423 ( .A(n8877), .Z(n8893) );
  BUF_X1 U13424 ( .A(n8877), .Z(n8894) );
  BUF_X1 U13425 ( .A(n8877), .Z(n8899) );
  BUF_X1 U13426 ( .A(n8900), .Z(n8902) );
  BUF_X1 U13427 ( .A(n8900), .Z(n8903) );
  BUF_X1 U13428 ( .A(n8900), .Z(n8904) );
  BUF_X1 U13429 ( .A(n8900), .Z(n8905) );
  BUF_X1 U13430 ( .A(n8900), .Z(n8906) );
  BUF_X1 U13431 ( .A(n8900), .Z(n8907) );
  BUF_X1 U13432 ( .A(n8900), .Z(n8908) );
  BUF_X1 U13433 ( .A(n8901), .Z(n8913) );
  BUF_X1 U13434 ( .A(n8901), .Z(n8914) );
  BUF_X1 U13435 ( .A(n8901), .Z(n8915) );
  BUF_X1 U13436 ( .A(n8901), .Z(n8916) );
  BUF_X1 U13437 ( .A(n8901), .Z(n8917) );
  BUF_X1 U13438 ( .A(n8901), .Z(n8918) );
  BUF_X1 U13439 ( .A(n8901), .Z(n8923) );
  BUF_X1 U13440 ( .A(n8924), .Z(n8926) );
  BUF_X1 U13441 ( .A(n8924), .Z(n8927) );
  BUF_X1 U13442 ( .A(n8924), .Z(n8928) );
  BUF_X1 U13443 ( .A(n8924), .Z(n8929) );
  BUF_X1 U13444 ( .A(n8924), .Z(n8930) );
  BUF_X1 U13445 ( .A(n8924), .Z(n8931) );
  BUF_X1 U13446 ( .A(n8924), .Z(n8932) );
  BUF_X1 U13447 ( .A(n8925), .Z(n8937) );
  BUF_X1 U13448 ( .A(n8925), .Z(n8938) );
  BUF_X1 U13449 ( .A(n8925), .Z(n8939) );
  BUF_X1 U13450 ( .A(n8925), .Z(n8940) );
  BUF_X1 U13451 ( .A(n8925), .Z(n8941) );
  BUF_X1 U13452 ( .A(n8925), .Z(n8942) );
  BUF_X1 U13453 ( .A(n8925), .Z(n8947) );
  BUF_X1 U13454 ( .A(n8948), .Z(n8950) );
  BUF_X1 U13455 ( .A(n8948), .Z(n8951) );
  BUF_X1 U13456 ( .A(n8948), .Z(n8952) );
  BUF_X1 U13457 ( .A(n8948), .Z(n8953) );
  BUF_X1 U13458 ( .A(n8948), .Z(n8954) );
  BUF_X1 U13459 ( .A(n8948), .Z(n8955) );
  BUF_X1 U13460 ( .A(n8948), .Z(n8956) );
  BUF_X1 U13461 ( .A(n8949), .Z(n8961) );
  BUF_X1 U13462 ( .A(n8949), .Z(n8962) );
  BUF_X1 U13463 ( .A(n8949), .Z(n8963) );
  BUF_X1 U13464 ( .A(n8949), .Z(n8964) );
  BUF_X1 U13465 ( .A(n8949), .Z(n8965) );
  BUF_X1 U13466 ( .A(n8949), .Z(n8966) );
  BUF_X1 U13467 ( .A(n8949), .Z(n8971) );
  BUF_X1 U13468 ( .A(n8972), .Z(n8974) );
  BUF_X1 U13469 ( .A(n8972), .Z(n8975) );
  BUF_X1 U13470 ( .A(n8972), .Z(n8976) );
  BUF_X1 U13471 ( .A(n8972), .Z(n8977) );
  BUF_X1 U13472 ( .A(n8972), .Z(n8978) );
  BUF_X1 U13473 ( .A(n8972), .Z(n8979) );
  BUF_X1 U13474 ( .A(n8972), .Z(n8980) );
  BUF_X1 U13475 ( .A(n8973), .Z(n8985) );
  BUF_X1 U13476 ( .A(n8973), .Z(n8986) );
  BUF_X1 U13477 ( .A(n8973), .Z(n8987) );
  BUF_X1 U13478 ( .A(n8973), .Z(n8988) );
  BUF_X1 U13479 ( .A(n8973), .Z(n8989) );
  BUF_X1 U13480 ( .A(n8973), .Z(n8990) );
  BUF_X1 U13481 ( .A(n8973), .Z(n8995) );
  BUF_X1 U13482 ( .A(n8996), .Z(n8998) );
  BUF_X1 U13483 ( .A(n8996), .Z(n8999) );
  BUF_X1 U13484 ( .A(n8996), .Z(n9000) );
  BUF_X1 U13485 ( .A(n8996), .Z(n9001) );
  BUF_X1 U13486 ( .A(n8996), .Z(n9002) );
  BUF_X1 U13487 ( .A(n8996), .Z(n9003) );
  BUF_X1 U13488 ( .A(n8996), .Z(n9004) );
  BUF_X1 U13489 ( .A(n8997), .Z(n9009) );
  BUF_X1 U13490 ( .A(n8997), .Z(n9010) );
  BUF_X1 U13491 ( .A(n8997), .Z(n9011) );
  BUF_X1 U13492 ( .A(n8997), .Z(n9012) );
  BUF_X1 U13493 ( .A(n8997), .Z(n9013) );
  BUF_X1 U13494 ( .A(n8997), .Z(n9014) );
  BUF_X1 U13495 ( .A(n8997), .Z(n9019) );
  BUF_X1 U13496 ( .A(n9020), .Z(n9022) );
  BUF_X1 U13497 ( .A(n9020), .Z(n9023) );
  BUF_X1 U13498 ( .A(n9020), .Z(n9024) );
  BUF_X1 U13499 ( .A(n9020), .Z(n9025) );
  BUF_X1 U13500 ( .A(n9020), .Z(n9026) );
  BUF_X1 U13501 ( .A(n9020), .Z(n9027) );
  BUF_X1 U13502 ( .A(n9020), .Z(n9028) );
  BUF_X1 U13503 ( .A(n9021), .Z(n9033) );
  BUF_X1 U13504 ( .A(n9021), .Z(n9034) );
  BUF_X1 U13505 ( .A(n9021), .Z(n9035) );
  BUF_X1 U13506 ( .A(n9021), .Z(n9036) );
  BUF_X1 U13507 ( .A(n9021), .Z(n9037) );
  BUF_X1 U13508 ( .A(n9021), .Z(n9038) );
  BUF_X1 U13509 ( .A(n9021), .Z(n9043) );
  BUF_X1 U13510 ( .A(n9044), .Z(n9046) );
  BUF_X1 U13511 ( .A(n9044), .Z(n9047) );
  BUF_X1 U13512 ( .A(n9044), .Z(n9048) );
  BUF_X1 U13513 ( .A(n9044), .Z(n9049) );
  BUF_X1 U13514 ( .A(n9044), .Z(n9050) );
  BUF_X1 U13515 ( .A(n9044), .Z(n9051) );
  BUF_X1 U13516 ( .A(n9044), .Z(n9052) );
  BUF_X1 U13517 ( .A(n9045), .Z(n9057) );
  BUF_X1 U13518 ( .A(n9045), .Z(n9058) );
  BUF_X1 U13519 ( .A(n9045), .Z(n9059) );
  BUF_X1 U13520 ( .A(n9045), .Z(n9060) );
  BUF_X1 U13521 ( .A(n9045), .Z(n9061) );
  BUF_X1 U13522 ( .A(n9045), .Z(n9062) );
  BUF_X1 U13523 ( .A(n9045), .Z(n9067) );
  BUF_X1 U13524 ( .A(n9068), .Z(n9070) );
  BUF_X1 U13525 ( .A(n9068), .Z(n9071) );
  BUF_X1 U13526 ( .A(n9068), .Z(n9072) );
  BUF_X1 U13527 ( .A(n9068), .Z(n9073) );
  BUF_X1 U13528 ( .A(n9068), .Z(n9074) );
  BUF_X1 U13529 ( .A(n9068), .Z(n9075) );
  BUF_X1 U13530 ( .A(n9068), .Z(n9076) );
  BUF_X1 U13531 ( .A(n9069), .Z(n9081) );
  BUF_X1 U13532 ( .A(n9069), .Z(n9082) );
  BUF_X1 U13533 ( .A(n9069), .Z(n9083) );
  BUF_X1 U13534 ( .A(n9069), .Z(n9084) );
  BUF_X1 U13535 ( .A(n9069), .Z(n9085) );
  BUF_X1 U13536 ( .A(n9069), .Z(n9086) );
  BUF_X1 U13537 ( .A(n9069), .Z(n9091) );
  BUF_X1 U13538 ( .A(n9092), .Z(n9094) );
  BUF_X1 U13539 ( .A(n9092), .Z(n9095) );
  BUF_X1 U13540 ( .A(n9092), .Z(n9096) );
  BUF_X1 U13541 ( .A(n9092), .Z(n9097) );
  BUF_X1 U13542 ( .A(n9092), .Z(n9098) );
  BUF_X1 U13543 ( .A(n9092), .Z(n9099) );
  BUF_X1 U13544 ( .A(n9092), .Z(n9100) );
  BUF_X1 U13545 ( .A(n9093), .Z(n9105) );
  BUF_X1 U13546 ( .A(n9093), .Z(n9106) );
  BUF_X1 U13547 ( .A(n9093), .Z(n9107) );
  BUF_X1 U13548 ( .A(n9093), .Z(n9108) );
  BUF_X1 U13549 ( .A(n9093), .Z(n9109) );
  BUF_X1 U13550 ( .A(n9093), .Z(n9110) );
  BUF_X1 U13551 ( .A(n9093), .Z(n9115) );
  BUF_X1 U13552 ( .A(n9116), .Z(n9118) );
  BUF_X1 U13553 ( .A(n9116), .Z(n9119) );
  BUF_X1 U13554 ( .A(n9116), .Z(n9120) );
  BUF_X1 U13555 ( .A(n9116), .Z(n9121) );
  BUF_X1 U13556 ( .A(n9116), .Z(n9122) );
  BUF_X1 U13557 ( .A(n9116), .Z(n9123) );
  BUF_X1 U13558 ( .A(n9116), .Z(n9124) );
  BUF_X1 U13559 ( .A(n9117), .Z(n9129) );
  BUF_X1 U13560 ( .A(n9117), .Z(n9130) );
  BUF_X1 U13561 ( .A(n9117), .Z(n9131) );
  BUF_X1 U13562 ( .A(n9117), .Z(n9132) );
  BUF_X1 U13563 ( .A(n9117), .Z(n9133) );
  BUF_X1 U13564 ( .A(n9117), .Z(n9134) );
  BUF_X1 U13565 ( .A(n9117), .Z(n9139) );
  BUF_X1 U13566 ( .A(n9140), .Z(n9142) );
  BUF_X1 U13567 ( .A(n9140), .Z(n9143) );
  BUF_X1 U13568 ( .A(n9140), .Z(n9144) );
  BUF_X1 U13569 ( .A(n9140), .Z(n9145) );
  BUF_X1 U13570 ( .A(n9140), .Z(n9146) );
  BUF_X1 U13571 ( .A(n9140), .Z(n9147) );
  BUF_X1 U13572 ( .A(n9140), .Z(n9148) );
  BUF_X1 U13573 ( .A(n9141), .Z(n9153) );
  BUF_X1 U13574 ( .A(n9141), .Z(n9154) );
  BUF_X1 U13575 ( .A(n9141), .Z(n9155) );
  BUF_X1 U13576 ( .A(n9141), .Z(n9156) );
  BUF_X1 U13577 ( .A(n9141), .Z(n9157) );
  BUF_X1 U13578 ( .A(n9141), .Z(n9158) );
  BUF_X1 U13579 ( .A(n9141), .Z(n9163) );
  BUF_X1 U13580 ( .A(n9164), .Z(n9166) );
  BUF_X1 U13581 ( .A(n9164), .Z(n9167) );
  BUF_X1 U13582 ( .A(n9164), .Z(n9168) );
  BUF_X1 U13583 ( .A(n9164), .Z(n9169) );
  BUF_X1 U13584 ( .A(n9164), .Z(n9170) );
  BUF_X1 U13585 ( .A(n9164), .Z(n9171) );
  BUF_X1 U13586 ( .A(n9164), .Z(n9172) );
  BUF_X1 U13587 ( .A(n9165), .Z(n9177) );
  BUF_X1 U13588 ( .A(n9165), .Z(n9178) );
  BUF_X1 U13589 ( .A(n9165), .Z(n9179) );
  BUF_X1 U13590 ( .A(n9165), .Z(n9180) );
  BUF_X1 U13591 ( .A(n9165), .Z(n9181) );
  BUF_X1 U13592 ( .A(n9165), .Z(n9182) );
  BUF_X1 U13593 ( .A(n9165), .Z(n9187) );
  BUF_X1 U13594 ( .A(n9188), .Z(n9190) );
  BUF_X1 U13595 ( .A(n9188), .Z(n9191) );
  BUF_X1 U13596 ( .A(n9188), .Z(n9192) );
  BUF_X1 U13597 ( .A(n9188), .Z(n9193) );
  BUF_X1 U13598 ( .A(n9188), .Z(n9194) );
  BUF_X1 U13599 ( .A(n9188), .Z(n9195) );
  BUF_X1 U13600 ( .A(n9188), .Z(n9196) );
  BUF_X1 U13601 ( .A(n9189), .Z(n9201) );
  BUF_X1 U13602 ( .A(n9189), .Z(n9202) );
  BUF_X1 U13603 ( .A(n9189), .Z(n9203) );
  BUF_X1 U13604 ( .A(n9189), .Z(n9204) );
  BUF_X1 U13605 ( .A(n9189), .Z(n9205) );
  BUF_X1 U13606 ( .A(n9189), .Z(n9206) );
  BUF_X1 U13607 ( .A(n9189), .Z(n9211) );
  BUF_X1 U13608 ( .A(n9212), .Z(n9214) );
  BUF_X1 U13609 ( .A(n9212), .Z(n9215) );
  BUF_X1 U13610 ( .A(n9212), .Z(n9216) );
  BUF_X1 U13611 ( .A(n9212), .Z(n9217) );
  BUF_X1 U13612 ( .A(n9212), .Z(n9218) );
  BUF_X1 U13613 ( .A(n9212), .Z(n9219) );
  BUF_X1 U13614 ( .A(n9212), .Z(n9220) );
  BUF_X1 U13615 ( .A(n9213), .Z(n9225) );
  BUF_X1 U13616 ( .A(n9213), .Z(n9226) );
  BUF_X1 U13617 ( .A(n9213), .Z(n9227) );
  BUF_X1 U13618 ( .A(n9213), .Z(n9228) );
  BUF_X1 U13619 ( .A(n9213), .Z(n9229) );
  BUF_X1 U13620 ( .A(n9213), .Z(n9230) );
  BUF_X1 U13621 ( .A(n9213), .Z(n9235) );
  INV_X1 U13622 ( .A(mem_access_addr[4]), .ZN(n9237) );
  INV_X1 U13623 ( .A(n9239), .ZN(n9238) );
  INV_X1 U13624 ( .A(mem_access_addr[6]), .ZN(n9239) );
  INV_X1 U13625 ( .A(mem_access_addr[8]), .ZN(n9240) );
endmodule


module mips_16 ( clk, reset, pc_out, alu_result );
  output [15:0] pc_out;
  output [15:0] alu_result;
  input clk, reset;
  wire   jump, branch, mem_read, mem_write, alu_src, reg_write,
         reg_write_dest_1_, JRControl, zero_flag, N54, n52, n530, n540, n55,
         n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69,
         n70, n71, n82, n83, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94,
         n95, n96, n97, n98, n99, n100, n101, n102, n103, n105, n106, n107,
         n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165,
         n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176,
         n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187,
         SYNOPSYS_UNCONNECTED_1, SYNOPSYS_UNCONNECTED_2,
         SYNOPSYS_UNCONNECTED_3, SYNOPSYS_UNCONNECTED_4,
         SYNOPSYS_UNCONNECTED_5, SYNOPSYS_UNCONNECTED_6,
         SYNOPSYS_UNCONNECTED_7, SYNOPSYS_UNCONNECTED_8,
         SYNOPSYS_UNCONNECTED_9, SYNOPSYS_UNCONNECTED_10,
         SYNOPSYS_UNCONNECTED_11, SYNOPSYS_UNCONNECTED_12,
         SYNOPSYS_UNCONNECTED_13, SYNOPSYS_UNCONNECTED_14,
         SYNOPSYS_UNCONNECTED_15, SYNOPSYS_UNCONNECTED_16;
  wire   [15:0] pc_next;
  wire   [15:0] instr;
  wire   [1:0] reg_dst;
  wire   [1:0] mem_to_reg;
  wire   [1:0] alu_op;
  wire   [15:0] reg_write_data;
  wire   [15:0] reg_read_data_1;
  wire   [15:0] reg_read_data_2;
  wire   [2:0] ALU_Control;
  wire   [6:0] read_data2;
  wire   [15:0] mem_read_data;

  DFFR_X1 pc_current_reg_15_ ( .D(pc_next[15]), .CK(clk), .RN(n186), .Q(
        pc_out[15]), .QN(n152) );
  NOR2_X2 U44 ( .A1(n185), .A2(mem_to_reg[1]), .ZN(n56) );
  instr_mem instrucion_memory ( .pc(pc_out), .instruction({
        SYNOPSYS_UNCONNECTED_1, SYNOPSYS_UNCONNECTED_2, SYNOPSYS_UNCONNECTED_3, 
        SYNOPSYS_UNCONNECTED_4, SYNOPSYS_UNCONNECTED_5, SYNOPSYS_UNCONNECTED_6, 
        SYNOPSYS_UNCONNECTED_7, SYNOPSYS_UNCONNECTED_8, SYNOPSYS_UNCONNECTED_9, 
        SYNOPSYS_UNCONNECTED_10, SYNOPSYS_UNCONNECTED_11, 
        SYNOPSYS_UNCONNECTED_12, SYNOPSYS_UNCONNECTED_13, 
        SYNOPSYS_UNCONNECTED_14, SYNOPSYS_UNCONNECTED_15, 
        SYNOPSYS_UNCONNECTED_16}) );
  control control_unit ( .opcode({1'b0, 1'b0, 1'b0}), .reset(reset), .reg_dst(
        reg_dst), .mem_to_reg(mem_to_reg), .alu_op(alu_op), .jump(jump), 
        .branch(branch), .mem_read(mem_read), .mem_write(mem_write), .alu_src(
        alu_src), .reg_write(reg_write) );
  register_file reg_file ( .clk(clk), .rst(reset), .reg_write_en(reg_write), 
        .reg_write_dest({reg_write_dest_1_, reg_write_dest_1_, 
        reg_write_dest_1_}), .reg_write_data(reg_write_data), 
        .reg_read_addr_1({1'b0, 1'b0, 1'b0}), .reg_read_data_1(reg_read_data_1), .reg_read_addr_2({1'b0, 1'b0, 1'b0}), .reg_read_data_2(reg_read_data_2) );
  JR_Control JRControl_unit ( .alu_op(alu_op), .funct({1'b0, 1'b0, 1'b0, 1'b0}), .JRControl(JRControl) );
  ALUControl ALU_Control_unit ( .ALU_Control(ALU_Control), .ALUOp(alu_op), 
        .Function({1'b0, 1'b0, 1'b0, 1'b0}) );
  alu alu_unit ( .a(reg_read_data_1), .b({n124, n132, n131, n127, n130, n126, 
        n129, n125, n128, read_data2}), .alu_control(ALU_Control), .result(
        alu_result), .zero(zero_flag) );
  data_memory datamem ( .clk(clk), .mem_access_addr(alu_result), 
        .mem_write_data(reg_read_data_2), .mem_write_en(mem_write), .mem_read(
        mem_read), .mem_read_data(mem_read_data) );
  DFFR_X1 pc_current_reg_0_ ( .D(pc_next[0]), .CK(clk), .RN(n186), .Q(
        pc_out[0]), .QN(n187) );
  DFFR_X1 pc_current_reg_1_ ( .D(pc_next[1]), .CK(clk), .RN(n186), .Q(
        pc_out[1]), .QN(N54) );
  DFFR_X1 pc_current_reg_2_ ( .D(pc_next[2]), .CK(clk), .RN(n186), .Q(
        pc_out[2]) );
  DFFR_X1 pc_current_reg_3_ ( .D(pc_next[3]), .CK(clk), .RN(n186), .Q(
        pc_out[3]) );
  DFFR_X1 pc_current_reg_4_ ( .D(pc_next[4]), .CK(clk), .RN(n186), .Q(
        pc_out[4]) );
  DFFR_X1 pc_current_reg_5_ ( .D(pc_next[5]), .CK(clk), .RN(n186), .Q(
        pc_out[5]) );
  DFFR_X1 pc_current_reg_6_ ( .D(pc_next[6]), .CK(clk), .RN(n186), .Q(
        pc_out[6]) );
  DFFR_X1 pc_current_reg_7_ ( .D(pc_next[7]), .CK(clk), .RN(n186), .Q(
        pc_out[7]) );
  DFFR_X1 pc_current_reg_8_ ( .D(pc_next[8]), .CK(clk), .RN(n186), .Q(
        pc_out[8]) );
  DFFR_X1 pc_current_reg_9_ ( .D(pc_next[9]), .CK(clk), .RN(n186), .Q(
        pc_out[9]) );
  DFFR_X1 pc_current_reg_10_ ( .D(pc_next[10]), .CK(clk), .RN(n186), .Q(
        pc_out[10]) );
  DFFR_X1 pc_current_reg_11_ ( .D(pc_next[11]), .CK(clk), .RN(n186), .Q(
        pc_out[11]) );
  DFFR_X1 pc_current_reg_12_ ( .D(pc_next[12]), .CK(clk), .RN(n186), .Q(
        pc_out[12]) );
  DFFR_X1 pc_current_reg_13_ ( .D(pc_next[13]), .CK(clk), .RN(n186), .Q(
        pc_out[13]) );
  DFFR_X1 pc_current_reg_14_ ( .D(pc_next[14]), .CK(clk), .RN(n186), .Q(
        pc_out[14]) );
  XNOR2_X1 U170 ( .A(n152), .B(n159), .ZN(n122) );
  NOR3_X4 U171 ( .A1(JRControl), .A2(jump), .A3(n167), .ZN(n86) );
  INV_X1 U172 ( .A(n123), .ZN(n168) );
  OAI21_X1 U173 ( .B1(n530), .B2(n122), .A(n65), .ZN(reg_write_data[15]) );
  AOI22_X1 U174 ( .A1(alu_result[15]), .A2(n55), .B1(mem_read_data[15]), .B2(
        n56), .ZN(n65) );
  INV_X1 U175 ( .A(n52), .ZN(reg_write_dest_1_) );
  INV_X1 U176 ( .A(mem_to_reg[0]), .ZN(n185) );
  AND2_X1 U177 ( .A1(jump), .A2(n182), .ZN(n85) );
  OAI221_X1 U178 ( .B1(n103), .B2(n122), .C1(n123), .C2(n122), .A(n105), .ZN(
        pc_next[15]) );
  AOI21_X1 U179 ( .B1(n106), .B2(n182), .A(n85), .ZN(n103) );
  NAND2_X1 U180 ( .A1(reg_read_data_1[15]), .A2(JRControl), .ZN(n105) );
  NAND2_X1 U181 ( .A1(n115), .A2(n116), .ZN(pc_next[10]) );
  NAND2_X1 U182 ( .A1(n136), .A2(n168), .ZN(n116) );
  AOI22_X1 U183 ( .A1(n86), .A2(n136), .B1(reg_read_data_1[10]), .B2(JRControl), .ZN(n115) );
  NAND2_X1 U184 ( .A1(n113), .A2(n114), .ZN(pc_next[11]) );
  NAND2_X1 U185 ( .A1(n137), .A2(n168), .ZN(n114) );
  AOI22_X1 U186 ( .A1(n86), .A2(n137), .B1(reg_read_data_1[11]), .B2(JRControl), .ZN(n113) );
  NAND2_X1 U187 ( .A1(n111), .A2(n112), .ZN(pc_next[12]) );
  NAND2_X1 U188 ( .A1(n138), .A2(n168), .ZN(n112) );
  AOI22_X1 U189 ( .A1(n86), .A2(n138), .B1(reg_read_data_1[12]), .B2(JRControl), .ZN(n111) );
  NAND2_X1 U190 ( .A1(n109), .A2(n110), .ZN(pc_next[13]) );
  NAND2_X1 U191 ( .A1(n139), .A2(n168), .ZN(n110) );
  AOI22_X1 U192 ( .A1(n86), .A2(n139), .B1(reg_read_data_1[13]), .B2(JRControl), .ZN(n109) );
  NAND2_X1 U193 ( .A1(n107), .A2(n108), .ZN(pc_next[14]) );
  NAND2_X1 U194 ( .A1(n140), .A2(n168), .ZN(n108) );
  AOI22_X1 U195 ( .A1(n86), .A2(n140), .B1(reg_read_data_1[14]), .B2(JRControl), .ZN(n107) );
  NAND2_X1 U196 ( .A1(n89), .A2(n90), .ZN(pc_next[7]) );
  NAND2_X1 U197 ( .A1(n133), .A2(n168), .ZN(n90) );
  AOI22_X1 U198 ( .A1(n86), .A2(n133), .B1(reg_read_data_1[7]), .B2(JRControl), 
        .ZN(n89) );
  NAND2_X1 U199 ( .A1(n87), .A2(n88), .ZN(pc_next[8]) );
  NAND2_X1 U200 ( .A1(n134), .A2(n168), .ZN(n88) );
  AOI22_X1 U201 ( .A1(n86), .A2(n134), .B1(reg_read_data_1[8]), .B2(JRControl), 
        .ZN(n87) );
  NAND2_X1 U202 ( .A1(n82), .A2(n83), .ZN(pc_next[9]) );
  NAND2_X1 U203 ( .A1(n135), .A2(n168), .ZN(n83) );
  AOI22_X1 U204 ( .A1(n86), .A2(n135), .B1(reg_read_data_1[9]), .B2(JRControl), 
        .ZN(n82) );
  NAND2_X1 U205 ( .A1(n99), .A2(n100), .ZN(pc_next[2]) );
  NAND2_X1 U206 ( .A1(n158), .A2(n168), .ZN(n100) );
  AOI22_X1 U207 ( .A1(n86), .A2(n158), .B1(reg_read_data_1[2]), .B2(JRControl), 
        .ZN(n99) );
  NAND2_X1 U208 ( .A1(n97), .A2(n98), .ZN(pc_next[3]) );
  NAND2_X1 U209 ( .A1(n154), .A2(n168), .ZN(n98) );
  AOI22_X1 U210 ( .A1(n86), .A2(n154), .B1(reg_read_data_1[3]), .B2(JRControl), 
        .ZN(n97) );
  NAND2_X1 U211 ( .A1(n93), .A2(n94), .ZN(pc_next[5]) );
  NAND2_X1 U212 ( .A1(n156), .A2(n168), .ZN(n94) );
  AOI22_X1 U213 ( .A1(n86), .A2(n156), .B1(reg_read_data_1[5]), .B2(JRControl), 
        .ZN(n93) );
  NAND2_X1 U214 ( .A1(n91), .A2(n92), .ZN(pc_next[6]) );
  NAND2_X1 U215 ( .A1(n157), .A2(n168), .ZN(n92) );
  AOI22_X1 U216 ( .A1(n86), .A2(n157), .B1(reg_read_data_1[6]), .B2(JRControl), 
        .ZN(n91) );
  NAND2_X1 U217 ( .A1(n95), .A2(n96), .ZN(pc_next[4]) );
  NAND2_X1 U218 ( .A1(n155), .A2(n168), .ZN(n96) );
  AOI22_X1 U219 ( .A1(n86), .A2(n155), .B1(reg_read_data_1[4]), .B2(JRControl), 
        .ZN(n95) );
  INV_X1 U220 ( .A(n106), .ZN(n167) );
  NAND2_X1 U221 ( .A1(mem_to_reg[1]), .A2(n185), .ZN(n530) );
  INV_X1 U222 ( .A(JRControl), .ZN(n182) );
  NOR2_X1 U223 ( .A1(alu_src), .A2(n160), .ZN(read_data2[0]) );
  NOR2_X1 U224 ( .A1(alu_src), .A2(n162), .ZN(read_data2[2]) );
  NOR2_X1 U225 ( .A1(alu_src), .A2(n164), .ZN(read_data2[4]) );
  NOR2_X1 U226 ( .A1(alu_src), .A2(n166), .ZN(read_data2[6]) );
  NOR2_X1 U227 ( .A1(alu_src), .A2(n163), .ZN(read_data2[3]) );
  NOR2_X1 U228 ( .A1(alu_src), .A2(n165), .ZN(read_data2[5]) );
  INV_X1 U229 ( .A(alu_src), .ZN(n184) );
  NOR2_X1 U230 ( .A1(alu_src), .A2(n161), .ZN(read_data2[1]) );
  OAI21_X1 U231 ( .B1(n530), .B2(n181), .A(n63), .ZN(reg_write_data[2]) );
  INV_X1 U232 ( .A(n158), .ZN(n181) );
  AOI22_X1 U233 ( .A1(alu_result[2]), .A2(n55), .B1(mem_read_data[2]), .B2(n56), .ZN(n63) );
  OAI21_X1 U234 ( .B1(n530), .B2(n180), .A(n62), .ZN(reg_write_data[3]) );
  INV_X1 U235 ( .A(n154), .ZN(n180) );
  AOI22_X1 U236 ( .A1(alu_result[3]), .A2(n55), .B1(mem_read_data[3]), .B2(n56), .ZN(n62) );
  OAI21_X1 U237 ( .B1(n530), .B2(n179), .A(n61), .ZN(reg_write_data[4]) );
  INV_X1 U238 ( .A(n155), .ZN(n179) );
  AOI22_X1 U239 ( .A1(alu_result[4]), .A2(n55), .B1(mem_read_data[4]), .B2(n56), .ZN(n61) );
  OAI21_X1 U240 ( .B1(n530), .B2(n178), .A(n60), .ZN(reg_write_data[5]) );
  INV_X1 U241 ( .A(n156), .ZN(n178) );
  AOI22_X1 U242 ( .A1(alu_result[5]), .A2(n55), .B1(mem_read_data[5]), .B2(n56), .ZN(n60) );
  OAI21_X1 U243 ( .B1(n530), .B2(n177), .A(n59), .ZN(reg_write_data[6]) );
  INV_X1 U244 ( .A(n157), .ZN(n177) );
  AOI22_X1 U245 ( .A1(alu_result[6]), .A2(n55), .B1(mem_read_data[6]), .B2(n56), .ZN(n59) );
  OAI21_X1 U246 ( .B1(n530), .B2(n176), .A(n58), .ZN(reg_write_data[7]) );
  INV_X1 U247 ( .A(n133), .ZN(n176) );
  AOI22_X1 U248 ( .A1(alu_result[7]), .A2(n55), .B1(mem_read_data[7]), .B2(n56), .ZN(n58) );
  OAI21_X1 U249 ( .B1(n530), .B2(n175), .A(n57), .ZN(reg_write_data[8]) );
  INV_X1 U250 ( .A(n134), .ZN(n175) );
  AOI22_X1 U251 ( .A1(alu_result[8]), .A2(n55), .B1(mem_read_data[8]), .B2(n56), .ZN(n57) );
  OAI21_X1 U252 ( .B1(n530), .B2(n174), .A(n540), .ZN(reg_write_data[9]) );
  INV_X1 U253 ( .A(n135), .ZN(n174) );
  AOI22_X1 U254 ( .A1(alu_result[9]), .A2(n55), .B1(mem_read_data[9]), .B2(n56), .ZN(n540) );
  OAI21_X1 U255 ( .B1(n530), .B2(n173), .A(n70), .ZN(reg_write_data[10]) );
  INV_X1 U256 ( .A(n136), .ZN(n173) );
  AOI22_X1 U257 ( .A1(alu_result[10]), .A2(n55), .B1(mem_read_data[10]), .B2(
        n56), .ZN(n70) );
  OAI21_X1 U258 ( .B1(n530), .B2(n172), .A(n69), .ZN(reg_write_data[11]) );
  INV_X1 U259 ( .A(n137), .ZN(n172) );
  AOI22_X1 U260 ( .A1(alu_result[11]), .A2(n55), .B1(mem_read_data[11]), .B2(
        n56), .ZN(n69) );
  OAI21_X1 U261 ( .B1(n530), .B2(n171), .A(n68), .ZN(reg_write_data[12]) );
  INV_X1 U262 ( .A(n138), .ZN(n171) );
  AOI22_X1 U263 ( .A1(alu_result[12]), .A2(n55), .B1(mem_read_data[12]), .B2(
        n56), .ZN(n68) );
  OAI21_X1 U264 ( .B1(n530), .B2(n170), .A(n67), .ZN(reg_write_data[13]) );
  INV_X1 U265 ( .A(n139), .ZN(n170) );
  AOI22_X1 U266 ( .A1(alu_result[13]), .A2(n55), .B1(mem_read_data[13]), .B2(
        n56), .ZN(n67) );
  OAI21_X1 U267 ( .B1(n530), .B2(n169), .A(n66), .ZN(reg_write_data[14]) );
  INV_X1 U268 ( .A(n140), .ZN(n169) );
  AOI22_X1 U269 ( .A1(alu_result[14]), .A2(n55), .B1(mem_read_data[14]), .B2(
        n56), .ZN(n66) );
  NAND2_X1 U270 ( .A1(reg_dst[1]), .A2(n183), .ZN(n52) );
  INV_X1 U271 ( .A(reg_dst[0]), .ZN(n183) );
  OR3_X1 U272 ( .A1(JRControl), .A2(jump), .A3(n106), .ZN(n123) );
  AND2_X1 U273 ( .A1(reg_read_data_2[15]), .A2(n184), .ZN(n124) );
  AND2_X1 U274 ( .A1(reg_read_data_2[8]), .A2(n184), .ZN(n125) );
  AND2_X1 U275 ( .A1(reg_read_data_2[10]), .A2(n184), .ZN(n126) );
  AND2_X1 U276 ( .A1(reg_read_data_2[12]), .A2(n184), .ZN(n127) );
  AND2_X1 U277 ( .A1(reg_read_data_2[7]), .A2(n184), .ZN(n128) );
  AND2_X1 U278 ( .A1(reg_read_data_2[9]), .A2(n184), .ZN(n129) );
  AND2_X1 U279 ( .A1(reg_read_data_2[11]), .A2(n184), .ZN(n130) );
  AND2_X1 U280 ( .A1(reg_read_data_2[13]), .A2(n184), .ZN(n131) );
  NAND2_X1 U281 ( .A1(zero_flag), .A2(branch), .ZN(n106) );
  AND2_X1 U282 ( .A1(reg_read_data_2[14]), .A2(n184), .ZN(n132) );
  XOR2_X1 U283 ( .A(pc_out[7]), .B(n144), .Z(n133) );
  XOR2_X1 U284 ( .A(pc_out[8]), .B(n145), .Z(n134) );
  XOR2_X1 U285 ( .A(pc_out[9]), .B(n146), .Z(n135) );
  XOR2_X1 U286 ( .A(pc_out[10]), .B(n147), .Z(n136) );
  XOR2_X1 U287 ( .A(pc_out[11]), .B(n148), .Z(n137) );
  XOR2_X1 U288 ( .A(pc_out[12]), .B(n149), .Z(n138) );
  XOR2_X1 U289 ( .A(pc_out[13]), .B(n150), .Z(n139) );
  XOR2_X1 U290 ( .A(pc_out[14]), .B(n151), .Z(n140) );
  AND2_X1 U291 ( .A1(pc_out[1]), .A2(pc_out[2]), .ZN(n141) );
  AND2_X1 U292 ( .A1(n141), .A2(pc_out[3]), .ZN(n142) );
  AND2_X1 U293 ( .A1(n142), .A2(pc_out[4]), .ZN(n143) );
  AND2_X1 U294 ( .A1(n153), .A2(pc_out[6]), .ZN(n144) );
  AND2_X1 U295 ( .A1(n144), .A2(pc_out[7]), .ZN(n145) );
  AND2_X1 U296 ( .A1(n145), .A2(pc_out[8]), .ZN(n146) );
  AND2_X1 U297 ( .A1(n146), .A2(pc_out[9]), .ZN(n147) );
  AND2_X1 U298 ( .A1(n147), .A2(pc_out[10]), .ZN(n148) );
  AND2_X1 U299 ( .A1(n148), .A2(pc_out[11]), .ZN(n149) );
  AND2_X1 U300 ( .A1(n149), .A2(pc_out[12]), .ZN(n150) );
  AND2_X1 U301 ( .A1(n150), .A2(pc_out[13]), .ZN(n151) );
  NAND2_X1 U302 ( .A1(n151), .A2(pc_out[14]), .ZN(n159) );
  AND2_X1 U303 ( .A1(n143), .A2(pc_out[5]), .ZN(n153) );
  XOR2_X1 U304 ( .A(pc_out[3]), .B(n141), .Z(n154) );
  XOR2_X1 U305 ( .A(pc_out[4]), .B(n142), .Z(n155) );
  XOR2_X1 U306 ( .A(pc_out[5]), .B(n143), .Z(n156) );
  XOR2_X1 U307 ( .A(pc_out[6]), .B(n153), .Z(n157) );
  XOR2_X1 U308 ( .A(pc_out[2]), .B(pc_out[1]), .Z(n158) );
  NAND2_X1 U309 ( .A1(n117), .A2(n118), .ZN(pc_next[0]) );
  NAND2_X1 U310 ( .A1(pc_out[0]), .A2(n168), .ZN(n118) );
  AOI22_X1 U311 ( .A1(n86), .A2(pc_out[0]), .B1(reg_read_data_1[0]), .B2(
        JRControl), .ZN(n117) );
  NAND2_X1 U312 ( .A1(n101), .A2(n102), .ZN(pc_next[1]) );
  NAND2_X1 U313 ( .A1(N54), .A2(n168), .ZN(n102) );
  AOI22_X1 U314 ( .A1(n86), .A2(N54), .B1(reg_read_data_1[1]), .B2(JRControl), 
        .ZN(n101) );
  INV_X1 U315 ( .A(reset), .ZN(n186) );
  OAI21_X1 U316 ( .B1(n530), .B2(n187), .A(n71), .ZN(reg_write_data[0]) );
  AOI22_X1 U317 ( .A1(alu_result[0]), .A2(n55), .B1(mem_read_data[0]), .B2(n56), .ZN(n71) );
  OAI21_X1 U318 ( .B1(n530), .B2(pc_out[1]), .A(n64), .ZN(reg_write_data[1])
         );
  AOI22_X1 U319 ( .A1(alu_result[1]), .A2(n55), .B1(mem_read_data[1]), .B2(n56), .ZN(n64) );
  XOR2_X2 U320 ( .A(n185), .B(mem_to_reg[1]), .Z(n55) );
  INV_X1 U321 ( .A(reg_read_data_2[0]), .ZN(n160) );
  INV_X1 U322 ( .A(reg_read_data_2[1]), .ZN(n161) );
  INV_X1 U323 ( .A(reg_read_data_2[2]), .ZN(n162) );
  INV_X1 U324 ( .A(reg_read_data_2[3]), .ZN(n163) );
  INV_X1 U325 ( .A(reg_read_data_2[4]), .ZN(n164) );
  INV_X1 U326 ( .A(reg_read_data_2[5]), .ZN(n165) );
  INV_X1 U327 ( .A(reg_read_data_2[6]), .ZN(n166) );
endmodule

