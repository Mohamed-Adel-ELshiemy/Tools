
module cortexm0ds_logic_DW01_inc_0 ( A, SUM );
  input [30:0] A;
  output [30:0] SUM;

  wire   [30:2] carry;

  HA_X1 U1_1_29 ( .A(A[29]), .B(carry[29]), .CO(carry[30]), .S(SUM[29]) );
  HA_X1 U1_1_28 ( .A(A[28]), .B(carry[28]), .CO(carry[29]), .S(SUM[28]) );
  HA_X1 U1_1_27 ( .A(A[27]), .B(carry[27]), .CO(carry[28]), .S(SUM[27]) );
  HA_X1 U1_1_26 ( .A(A[26]), .B(carry[26]), .CO(carry[27]), .S(SUM[26]) );
  HA_X1 U1_1_25 ( .A(A[25]), .B(carry[25]), .CO(carry[26]), .S(SUM[25]) );
  HA_X1 U1_1_24 ( .A(A[24]), .B(carry[24]), .CO(carry[25]), .S(SUM[24]) );
  HA_X1 U1_1_23 ( .A(A[23]), .B(carry[23]), .CO(carry[24]), .S(SUM[23]) );
  HA_X1 U1_1_22 ( .A(A[22]), .B(carry[22]), .CO(carry[23]), .S(SUM[22]) );
  HA_X1 U1_1_21 ( .A(A[21]), .B(carry[21]), .CO(carry[22]), .S(SUM[21]) );
  HA_X1 U1_1_20 ( .A(A[20]), .B(carry[20]), .CO(carry[21]), .S(SUM[20]) );
  HA_X1 U1_1_19 ( .A(A[19]), .B(carry[19]), .CO(carry[20]), .S(SUM[19]) );
  HA_X1 U1_1_18 ( .A(A[18]), .B(carry[18]), .CO(carry[19]), .S(SUM[18]) );
  HA_X1 U1_1_17 ( .A(A[17]), .B(carry[17]), .CO(carry[18]), .S(SUM[17]) );
  HA_X1 U1_1_16 ( .A(A[16]), .B(carry[16]), .CO(carry[17]), .S(SUM[16]) );
  HA_X1 U1_1_15 ( .A(A[15]), .B(carry[15]), .CO(carry[16]), .S(SUM[15]) );
  HA_X1 U1_1_14 ( .A(A[14]), .B(carry[14]), .CO(carry[15]), .S(SUM[14]) );
  HA_X1 U1_1_13 ( .A(A[13]), .B(carry[13]), .CO(carry[14]), .S(SUM[13]) );
  HA_X1 U1_1_12 ( .A(A[12]), .B(carry[12]), .CO(carry[13]), .S(SUM[12]) );
  HA_X1 U1_1_11 ( .A(A[11]), .B(carry[11]), .CO(carry[12]), .S(SUM[11]) );
  HA_X1 U1_1_10 ( .A(A[10]), .B(carry[10]), .CO(carry[11]), .S(SUM[10]) );
  HA_X1 U1_1_9 ( .A(A[9]), .B(carry[9]), .CO(carry[10]), .S(SUM[9]) );
  HA_X1 U1_1_8 ( .A(A[8]), .B(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  HA_X1 U1_1_7 ( .A(A[7]), .B(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  HA_X1 U1_1_6 ( .A(A[6]), .B(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  HA_X1 U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  HA_X1 U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  HA_X1 U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  HA_X1 U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  HA_X1 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .S(SUM[1]) );
  XOR2_X1 U1 ( .A(carry[30]), .B(A[30]), .Z(SUM[30]) );
  INV_X1 U2 ( .A(A[0]), .ZN(SUM[0]) );
endmodule


module cortexm0ds_logic_DW01_dec_1 ( A, SUM );
  input [23:0] A;
  output [23:0] SUM;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55;

  INV_X1 U1 ( .A(n49), .ZN(n8) );
  INV_X1 U2 ( .A(n48), .ZN(n7) );
  INV_X1 U3 ( .A(n40), .ZN(n14) );
  INV_X1 U4 ( .A(n39), .ZN(n13) );
  INV_X1 U5 ( .A(n38), .ZN(n12) );
  INV_X1 U6 ( .A(n37), .ZN(n11) );
  INV_X1 U7 ( .A(n47), .ZN(n6) );
  INV_X1 U8 ( .A(n46), .ZN(n5) );
  INV_X1 U9 ( .A(n45), .ZN(n4) );
  INV_X1 U10 ( .A(n36), .ZN(n10) );
  INV_X1 U11 ( .A(A[1]), .ZN(n26) );
  INV_X1 U12 ( .A(A[14]), .ZN(n29) );
  INV_X1 U13 ( .A(A[15]), .ZN(n28) );
  INV_X1 U14 ( .A(A[2]), .ZN(n25) );
  INV_X1 U15 ( .A(A[3]), .ZN(n24) );
  INV_X1 U16 ( .A(A[4]), .ZN(n23) );
  INV_X1 U17 ( .A(A[6]), .ZN(n22) );
  INV_X1 U18 ( .A(A[16]), .ZN(n20) );
  INV_X1 U19 ( .A(A[17]), .ZN(n19) );
  INV_X1 U20 ( .A(A[18]), .ZN(n18) );
  INV_X1 U21 ( .A(A[19]), .ZN(n17) );
  INV_X1 U22 ( .A(A[5]), .ZN(n3) );
  INV_X1 U23 ( .A(n50), .ZN(n9) );
  OR2_X1 U24 ( .A1(n10), .A2(A[6]), .ZN(n1) );
  OR2_X1 U25 ( .A1(n4), .A2(A[19]), .ZN(n2) );
  INV_X1 U26 ( .A(A[8]), .ZN(n21) );
  INV_X1 U27 ( .A(A[10]), .ZN(n27) );
  INV_X1 U28 ( .A(A[12]), .ZN(n16) );
  INV_X1 U29 ( .A(A[21]), .ZN(n30) );
  INV_X1 U30 ( .A(A[0]), .ZN(SUM[0]) );
  INV_X1 U31 ( .A(n31), .ZN(SUM[9]) );
  AOI21_X1 U32 ( .B1(n32), .B2(A[9]), .A(n33), .ZN(n31) );
  OAI21_X1 U33 ( .B1(n34), .B2(n21), .A(n32), .ZN(SUM[8]) );
  INV_X1 U34 ( .A(n35), .ZN(SUM[7]) );
  AOI21_X1 U35 ( .B1(n1), .B2(A[7]), .A(n34), .ZN(n35) );
  OAI21_X1 U36 ( .B1(n36), .B2(n22), .A(n1), .ZN(SUM[6]) );
  OAI21_X1 U37 ( .B1(n37), .B2(n3), .A(n10), .ZN(SUM[5]) );
  OAI21_X1 U38 ( .B1(n38), .B2(n23), .A(n11), .ZN(SUM[4]) );
  OAI21_X1 U39 ( .B1(n39), .B2(n24), .A(n12), .ZN(SUM[3]) );
  OAI21_X1 U40 ( .B1(n40), .B2(n25), .A(n13), .ZN(SUM[2]) );
  XOR2_X1 U41 ( .A(A[23]), .B(n41), .Z(SUM[23]) );
  NOR2_X1 U42 ( .A1(A[22]), .A2(n42), .ZN(n41) );
  XNOR2_X1 U43 ( .A(A[22]), .B(n42), .ZN(SUM[22]) );
  OAI21_X1 U44 ( .B1(n43), .B2(n30), .A(n42), .ZN(SUM[21]) );
  NAND2_X1 U45 ( .A1(n43), .A2(n30), .ZN(n42) );
  INV_X1 U46 ( .A(n44), .ZN(SUM[20]) );
  AOI21_X1 U47 ( .B1(n2), .B2(A[20]), .A(n43), .ZN(n44) );
  NOR2_X1 U48 ( .A1(n2), .A2(A[20]), .ZN(n43) );
  OAI21_X1 U49 ( .B1(SUM[0]), .B2(n26), .A(n14), .ZN(SUM[1]) );
  OAI21_X1 U50 ( .B1(n45), .B2(n17), .A(n2), .ZN(SUM[19]) );
  OAI21_X1 U51 ( .B1(n46), .B2(n18), .A(n4), .ZN(SUM[18]) );
  NOR2_X1 U52 ( .A1(n5), .A2(A[18]), .ZN(n45) );
  OAI21_X1 U53 ( .B1(n47), .B2(n19), .A(n5), .ZN(SUM[17]) );
  NOR2_X1 U54 ( .A1(n6), .A2(A[17]), .ZN(n46) );
  OAI21_X1 U55 ( .B1(n48), .B2(n20), .A(n6), .ZN(SUM[16]) );
  NOR2_X1 U56 ( .A1(n7), .A2(A[16]), .ZN(n47) );
  OAI21_X1 U57 ( .B1(n49), .B2(n28), .A(n7), .ZN(SUM[15]) );
  NOR2_X1 U58 ( .A1(n8), .A2(A[15]), .ZN(n48) );
  OAI21_X1 U59 ( .B1(n50), .B2(n29), .A(n8), .ZN(SUM[14]) );
  NOR2_X1 U60 ( .A1(n9), .A2(A[14]), .ZN(n49) );
  INV_X1 U61 ( .A(n51), .ZN(SUM[13]) );
  AOI21_X1 U62 ( .B1(n52), .B2(A[13]), .A(n50), .ZN(n51) );
  NOR2_X1 U63 ( .A1(n52), .A2(A[13]), .ZN(n50) );
  OAI21_X1 U64 ( .B1(n53), .B2(n16), .A(n52), .ZN(SUM[12]) );
  NAND2_X1 U65 ( .A1(n53), .A2(n16), .ZN(n52) );
  INV_X1 U66 ( .A(n54), .ZN(SUM[11]) );
  AOI21_X1 U67 ( .B1(n55), .B2(A[11]), .A(n53), .ZN(n54) );
  NOR2_X1 U68 ( .A1(n55), .A2(A[11]), .ZN(n53) );
  OAI21_X1 U69 ( .B1(n33), .B2(n27), .A(n55), .ZN(SUM[10]) );
  NAND2_X1 U70 ( .A1(n33), .A2(n27), .ZN(n55) );
  NOR2_X1 U71 ( .A1(n32), .A2(A[9]), .ZN(n33) );
  NAND2_X1 U72 ( .A1(n34), .A2(n21), .ZN(n32) );
  NOR2_X1 U73 ( .A1(n1), .A2(A[7]), .ZN(n34) );
  NOR2_X1 U74 ( .A1(n11), .A2(A[5]), .ZN(n36) );
  NOR2_X1 U75 ( .A1(n12), .A2(A[4]), .ZN(n37) );
  NOR2_X1 U76 ( .A1(n13), .A2(A[3]), .ZN(n38) );
  NOR2_X1 U77 ( .A1(n14), .A2(A[2]), .ZN(n39) );
  NOR2_X1 U78 ( .A1(A[1]), .A2(A[0]), .ZN(n40) );
endmodule


module cortexm0ds_logic_DW01_cmp6_4 ( A, B, TC, LT, GT, EQ, LE, GE, NE );
  input [31:0] A;
  input [31:0] B;
  input TC;
  output LT, GT, EQ, LE, GE, NE;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47;

  INV_X1 U1 ( .A(A[0]), .ZN(n2) );
  INV_X1 U2 ( .A(A[1]), .ZN(n1) );
  INV_X1 U3 ( .A(B[1]), .ZN(n3) );
  NOR4_X1 U4 ( .A1(n4), .A2(n5), .A3(n6), .A4(n7), .ZN(EQ) );
  NAND4_X1 U5 ( .A1(n8), .A2(n9), .A3(n10), .A4(n11), .ZN(n7) );
  XNOR2_X1 U6 ( .A(B[3]), .B(A[3]), .ZN(n11) );
  XNOR2_X1 U7 ( .A(B[4]), .B(A[4]), .ZN(n10) );
  XNOR2_X1 U8 ( .A(B[5]), .B(A[5]), .ZN(n9) );
  XNOR2_X1 U9 ( .A(B[6]), .B(A[6]), .ZN(n8) );
  NAND4_X1 U10 ( .A1(n12), .A2(n13), .A3(n14), .A4(n15), .ZN(n6) );
  OAI22_X1 U11 ( .A1(n16), .A2(n1), .B1(B[1]), .B2(n16), .ZN(n15) );
  AND2_X1 U12 ( .A1(B[0]), .A2(n2), .ZN(n16) );
  OAI22_X1 U13 ( .A1(A[1]), .A2(n17), .B1(n17), .B2(n3), .ZN(n14) );
  NOR2_X1 U14 ( .A1(n2), .A2(B[0]), .ZN(n17) );
  XNOR2_X1 U15 ( .A(B[31]), .B(A[31]), .ZN(n13) );
  XNOR2_X1 U16 ( .A(B[2]), .B(A[2]), .ZN(n12) );
  NAND2_X1 U17 ( .A1(n18), .A2(n19), .ZN(n5) );
  NOR4_X1 U18 ( .A1(n20), .A2(n21), .A3(n22), .A4(n23), .ZN(n19) );
  XOR2_X1 U19 ( .A(B[10]), .B(A[10]), .Z(n23) );
  XOR2_X1 U20 ( .A(B[9]), .B(A[9]), .Z(n22) );
  XOR2_X1 U21 ( .A(B[8]), .B(A[8]), .Z(n21) );
  XOR2_X1 U22 ( .A(B[7]), .B(A[7]), .Z(n20) );
  NOR4_X1 U23 ( .A1(n24), .A2(n25), .A3(n26), .A4(n27), .ZN(n18) );
  XOR2_X1 U24 ( .A(B[14]), .B(A[14]), .Z(n27) );
  XOR2_X1 U25 ( .A(B[13]), .B(A[13]), .Z(n26) );
  XOR2_X1 U26 ( .A(B[12]), .B(A[12]), .Z(n25) );
  XOR2_X1 U27 ( .A(B[11]), .B(A[11]), .Z(n24) );
  NAND4_X1 U28 ( .A1(n28), .A2(n29), .A3(n30), .A4(n31), .ZN(n4) );
  NOR4_X1 U29 ( .A1(n32), .A2(n33), .A3(n34), .A4(n35), .ZN(n31) );
  XOR2_X1 U30 ( .A(B[18]), .B(A[18]), .Z(n35) );
  XOR2_X1 U31 ( .A(B[17]), .B(A[17]), .Z(n34) );
  XOR2_X1 U32 ( .A(B[16]), .B(A[16]), .Z(n33) );
  XOR2_X1 U33 ( .A(B[15]), .B(A[15]), .Z(n32) );
  NOR4_X1 U34 ( .A1(n36), .A2(n37), .A3(n38), .A4(n39), .ZN(n30) );
  XOR2_X1 U35 ( .A(B[22]), .B(A[22]), .Z(n39) );
  XOR2_X1 U36 ( .A(B[21]), .B(A[21]), .Z(n38) );
  XOR2_X1 U37 ( .A(B[20]), .B(A[20]), .Z(n37) );
  XOR2_X1 U38 ( .A(B[19]), .B(A[19]), .Z(n36) );
  NOR4_X1 U39 ( .A1(n40), .A2(n41), .A3(n42), .A4(n43), .ZN(n29) );
  XOR2_X1 U40 ( .A(B[26]), .B(A[26]), .Z(n43) );
  XOR2_X1 U41 ( .A(B[25]), .B(A[25]), .Z(n42) );
  XOR2_X1 U42 ( .A(B[24]), .B(A[24]), .Z(n41) );
  XOR2_X1 U43 ( .A(B[23]), .B(A[23]), .Z(n40) );
  NOR4_X1 U44 ( .A1(n44), .A2(n45), .A3(n46), .A4(n47), .ZN(n28) );
  XOR2_X1 U45 ( .A(B[30]), .B(A[30]), .Z(n47) );
  XOR2_X1 U46 ( .A(B[29]), .B(A[29]), .Z(n46) );
  XOR2_X1 U47 ( .A(B[28]), .B(A[28]), .Z(n45) );
  XOR2_X1 U48 ( .A(B[27]), .B(A[27]), .Z(n44) );
endmodule


module cortexm0ds_logic_DW01_ash_0 ( A, DATA_TC, SH, SH_TC, B );
  input [30:0] A;
  input [4:0] SH;
  output [30:0] B;
  input DATA_TC, SH_TC;
  wire   \MR_int[1][30] , \ML_int[2][2] , \ML_int[3][6] , \ML_int[3][5] ,
         \ML_int[3][4] , \ML_int[3][2] , \ML_int[4][14] , \ML_int[4][13] ,
         \ML_int[4][12] , \ML_int[4][11] , \ML_int[4][10] , \ML_int[4][9] ,
         \ML_int[4][8] , \ML_int[5][30] , \ML_int[5][29] , \ML_int[5][28] ,
         \ML_int[5][27] , \ML_int[5][26] , \ML_int[5][25] , \ML_int[5][24] ,
         \ML_int[5][23] , \ML_int[5][22] , \ML_int[5][21] , \ML_int[5][20] ,
         \ML_int[5][19] , \ML_int[5][18] , \ML_int[5][17] , \ML_int[5][16] ,
         \ML_int[5][14] , \ML_int[5][13] , \ML_int[5][12] , \ML_int[5][11] ,
         \ML_int[5][10] , \ML_int[5][9] , \ML_int[5][8] , \ML_int[5][7] ,
         \ML_int[5][6] , \ML_int[5][5] , \ML_int[5][4] , \ML_int[5][3] ,
         \ML_int[5][2] , \ML_int[5][1] , \ML_int[5][0] , n1, n2, n3, n4, n5,
         n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n21,
         n22, n23, n24, n25, n26;
  assign \MR_int[1][30]  = SH[0];
  assign B[30] = \ML_int[5][30] ;
  assign B[29] = \ML_int[5][29] ;
  assign B[28] = \ML_int[5][28] ;
  assign B[27] = \ML_int[5][27] ;
  assign B[26] = \ML_int[5][26] ;
  assign B[25] = \ML_int[5][25] ;
  assign B[24] = \ML_int[5][24] ;
  assign B[23] = \ML_int[5][23] ;
  assign B[22] = \ML_int[5][22] ;
  assign B[21] = \ML_int[5][21] ;
  assign B[20] = \ML_int[5][20] ;
  assign B[19] = \ML_int[5][19] ;
  assign B[18] = \ML_int[5][18] ;
  assign B[17] = \ML_int[5][17] ;
  assign B[16] = \ML_int[5][16] ;
  assign B[14] = \ML_int[5][14] ;
  assign B[13] = \ML_int[5][13] ;
  assign B[12] = \ML_int[5][12] ;
  assign B[11] = \ML_int[5][11] ;
  assign B[10] = \ML_int[5][10] ;
  assign B[9] = \ML_int[5][9] ;
  assign B[8] = \ML_int[5][8] ;
  assign B[7] = \ML_int[5][7] ;
  assign B[6] = \ML_int[5][6] ;
  assign B[5] = \ML_int[5][5] ;
  assign B[4] = \ML_int[5][4] ;
  assign B[3] = \ML_int[5][3] ;
  assign B[2] = \ML_int[5][2] ;
  assign B[1] = \ML_int[5][1] ;
  assign B[0] = \ML_int[5][0] ;

  OR2_X1 U3 ( .A1(n2), .A2(SH[3]), .ZN(n1) );
  OR2_X1 U4 ( .A1(SH[1]), .A2(SH[2]), .ZN(n2) );
  OR2_X1 U5 ( .A1(SH[1]), .A2(\MR_int[1][30] ), .ZN(n3) );
  OR2_X1 U6 ( .A1(\MR_int[1][30] ), .A2(n2), .ZN(n4) );
  INV_X1 U7 ( .A(\ML_int[4][14] ), .ZN(n12) );
  INV_X1 U8 ( .A(\ML_int[4][10] ), .ZN(n8) );
  INV_X1 U9 ( .A(\ML_int[4][9] ), .ZN(n7) );
  INV_X1 U10 ( .A(\ML_int[4][8] ), .ZN(n6) );
  NAND2_X1 U11 ( .A1(SH[4]), .A2(n10), .ZN(\ML_int[5][28] ) );
  INV_X1 U12 ( .A(\ML_int[4][12] ), .ZN(n10) );
  NAND2_X1 U13 ( .A1(SH[4]), .A2(n9), .ZN(\ML_int[5][27] ) );
  INV_X1 U14 ( .A(\ML_int[4][11] ), .ZN(n9) );
  NAND2_X1 U15 ( .A1(SH[4]), .A2(n11), .ZN(\ML_int[5][29] ) );
  INV_X1 U16 ( .A(\ML_int[4][13] ), .ZN(n11) );
  INV_X1 U17 ( .A(SH[4]), .ZN(B[15]) );
  INV_X1 U18 ( .A(SH[3]), .ZN(n18) );
  NAND2_X1 U19 ( .A1(SH[3]), .A2(n15), .ZN(\ML_int[4][14] ) );
  INV_X1 U20 ( .A(\ML_int[3][6] ), .ZN(n15) );
  NAND2_X1 U21 ( .A1(SH[3]), .A2(n17), .ZN(\ML_int[4][13] ) );
  INV_X1 U22 ( .A(\ML_int[3][5] ), .ZN(n17) );
  NAND2_X1 U23 ( .A1(SH[3]), .A2(n14), .ZN(\ML_int[4][12] ) );
  INV_X1 U24 ( .A(\ML_int[3][4] ), .ZN(n14) );
  NAND2_X1 U25 ( .A1(SH[3]), .A2(SH[2]), .ZN(\ML_int[4][11] ) );
  NAND2_X1 U26 ( .A1(SH[3]), .A2(n16), .ZN(\ML_int[4][10] ) );
  INV_X1 U27 ( .A(\ML_int[3][2] ), .ZN(n16) );
  NAND2_X1 U28 ( .A1(SH[3]), .A2(n2), .ZN(\ML_int[4][9] ) );
  NAND2_X1 U29 ( .A1(SH[3]), .A2(n4), .ZN(\ML_int[4][8] ) );
  INV_X1 U30 ( .A(SH[2]), .ZN(n21) );
  NAND2_X1 U31 ( .A1(SH[2]), .A2(SH[1]), .ZN(\ML_int[3][5] ) );
  NAND2_X1 U32 ( .A1(SH[2]), .A2(n3), .ZN(\ML_int[3][4] ) );
  NAND2_X1 U33 ( .A1(SH[2]), .A2(n13), .ZN(\ML_int[3][6] ) );
  INV_X1 U34 ( .A(\ML_int[2][2] ), .ZN(n13) );
  NAND2_X1 U35 ( .A1(SH[1]), .A2(\MR_int[1][30] ), .ZN(\ML_int[2][2] ) );
  INV_X1 U36 ( .A(\MR_int[1][30] ), .ZN(n19) );
  OR2_X1 U37 ( .A1(\MR_int[1][30] ), .A2(n1), .ZN(n5) );
  NAND2_X1 U38 ( .A1(SH[4]), .A2(n6), .ZN(\ML_int[5][24] ) );
  NAND2_X1 U39 ( .A1(SH[4]), .A2(n7), .ZN(\ML_int[5][25] ) );
  NAND2_X1 U40 ( .A1(SH[4]), .A2(n8), .ZN(\ML_int[5][26] ) );
  NAND2_X1 U41 ( .A1(SH[4]), .A2(n22), .ZN(\ML_int[5][22] ) );
  NAND2_X1 U42 ( .A1(SH[4]), .A2(n12), .ZN(\ML_int[5][30] ) );
  NAND2_X1 U43 ( .A1(SH[4]), .A2(SH[3]), .ZN(\ML_int[5][23] ) );
  NAND2_X1 U44 ( .A1(SH[4]), .A2(n26), .ZN(\ML_int[5][18] ) );
  NAND2_X1 U45 ( .A1(SH[4]), .A2(n1), .ZN(\ML_int[5][17] ) );
  NAND2_X1 U46 ( .A1(SH[4]), .A2(n5), .ZN(\ML_int[5][16] ) );
  NAND2_X1 U47 ( .A1(SH[4]), .A2(n25), .ZN(\ML_int[5][19] ) );
  NAND2_X1 U48 ( .A1(SH[4]), .A2(n23), .ZN(\ML_int[5][21] ) );
  NAND2_X1 U49 ( .A1(SH[4]), .A2(n24), .ZN(\ML_int[5][20] ) );
  AND2_X1 U50 ( .A1(\ML_int[4][9] ), .A2(B[15]), .ZN(\ML_int[5][9] ) );
  AND2_X1 U51 ( .A1(\ML_int[4][8] ), .A2(B[15]), .ZN(\ML_int[5][8] ) );
  NOR2_X1 U52 ( .A1(SH[4]), .A2(SH[3]), .ZN(\ML_int[5][7] ) );
  NOR2_X1 U53 ( .A1(SH[4]), .A2(n22), .ZN(\ML_int[5][6] ) );
  NOR2_X1 U54 ( .A1(SH[4]), .A2(n23), .ZN(\ML_int[5][5] ) );
  NOR2_X1 U55 ( .A1(SH[4]), .A2(n24), .ZN(\ML_int[5][4] ) );
  NOR2_X1 U56 ( .A1(SH[4]), .A2(n25), .ZN(\ML_int[5][3] ) );
  NOR2_X1 U57 ( .A1(SH[4]), .A2(n26), .ZN(\ML_int[5][2] ) );
  AND2_X1 U58 ( .A1(\ML_int[4][14] ), .A2(B[15]), .ZN(\ML_int[5][14] ) );
  AND2_X1 U59 ( .A1(\ML_int[4][13] ), .A2(B[15]), .ZN(\ML_int[5][13] ) );
  AND2_X1 U60 ( .A1(\ML_int[4][12] ), .A2(B[15]), .ZN(\ML_int[5][12] ) );
  AND2_X1 U61 ( .A1(\ML_int[4][11] ), .A2(B[15]), .ZN(\ML_int[5][11] ) );
  AND2_X1 U62 ( .A1(\ML_int[4][10] ), .A2(B[15]), .ZN(\ML_int[5][10] ) );
  AND2_X1 U63 ( .A1(n19), .A2(\ML_int[5][1] ), .ZN(\ML_int[5][0] ) );
  NOR2_X1 U64 ( .A1(n1), .A2(SH[4]), .ZN(\ML_int[5][1] ) );
  NAND2_X1 U65 ( .A1(\ML_int[3][6] ), .A2(n18), .ZN(n22) );
  NAND2_X1 U66 ( .A1(\ML_int[3][5] ), .A2(n18), .ZN(n23) );
  NAND2_X1 U67 ( .A1(\ML_int[3][4] ), .A2(n18), .ZN(n24) );
  NAND2_X1 U68 ( .A1(n21), .A2(n18), .ZN(n25) );
  NAND2_X1 U69 ( .A1(\ML_int[3][2] ), .A2(n18), .ZN(n26) );
  AND2_X1 U70 ( .A1(\ML_int[2][2] ), .A2(n21), .ZN(\ML_int[3][2] ) );
endmodule


module cortexm0ds_logic_DW01_cmp6_5 ( A, B, TC, LT, GT, EQ, LE, GE, NE );
  input [31:0] A;
  input [31:0] B;
  input TC;
  output LT, GT, EQ, LE, GE, NE;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47;

  INV_X1 U1 ( .A(A[0]), .ZN(n2) );
  INV_X1 U2 ( .A(A[1]), .ZN(n1) );
  INV_X1 U3 ( .A(B[1]), .ZN(n3) );
  NOR4_X1 U4 ( .A1(n4), .A2(n5), .A3(n6), .A4(n7), .ZN(EQ) );
  NAND4_X1 U5 ( .A1(n8), .A2(n9), .A3(n10), .A4(n11), .ZN(n7) );
  XNOR2_X1 U6 ( .A(B[3]), .B(A[3]), .ZN(n11) );
  XNOR2_X1 U7 ( .A(B[4]), .B(A[4]), .ZN(n10) );
  XNOR2_X1 U8 ( .A(B[5]), .B(A[5]), .ZN(n9) );
  XNOR2_X1 U9 ( .A(B[6]), .B(A[6]), .ZN(n8) );
  NAND4_X1 U10 ( .A1(n12), .A2(n13), .A3(n14), .A4(n15), .ZN(n6) );
  OAI22_X1 U11 ( .A1(n16), .A2(n1), .B1(B[1]), .B2(n16), .ZN(n15) );
  AND2_X1 U12 ( .A1(B[0]), .A2(n2), .ZN(n16) );
  OAI22_X1 U13 ( .A1(A[1]), .A2(n17), .B1(n17), .B2(n3), .ZN(n14) );
  NOR2_X1 U14 ( .A1(n2), .A2(B[0]), .ZN(n17) );
  XNOR2_X1 U15 ( .A(B[31]), .B(A[31]), .ZN(n13) );
  XNOR2_X1 U16 ( .A(B[2]), .B(A[2]), .ZN(n12) );
  NAND2_X1 U17 ( .A1(n18), .A2(n19), .ZN(n5) );
  NOR4_X1 U18 ( .A1(n20), .A2(n21), .A3(n22), .A4(n23), .ZN(n19) );
  XOR2_X1 U19 ( .A(B[10]), .B(A[10]), .Z(n23) );
  XOR2_X1 U20 ( .A(B[9]), .B(A[9]), .Z(n22) );
  XOR2_X1 U21 ( .A(B[8]), .B(A[8]), .Z(n21) );
  XOR2_X1 U22 ( .A(B[7]), .B(A[7]), .Z(n20) );
  NOR4_X1 U23 ( .A1(n24), .A2(n25), .A3(n26), .A4(n27), .ZN(n18) );
  XOR2_X1 U24 ( .A(B[14]), .B(A[14]), .Z(n27) );
  XOR2_X1 U25 ( .A(B[13]), .B(A[13]), .Z(n26) );
  XOR2_X1 U26 ( .A(B[12]), .B(A[12]), .Z(n25) );
  XOR2_X1 U27 ( .A(B[11]), .B(A[11]), .Z(n24) );
  NAND4_X1 U28 ( .A1(n28), .A2(n29), .A3(n30), .A4(n31), .ZN(n4) );
  NOR4_X1 U29 ( .A1(n32), .A2(n33), .A3(n34), .A4(n35), .ZN(n31) );
  XOR2_X1 U30 ( .A(B[18]), .B(A[18]), .Z(n35) );
  XOR2_X1 U31 ( .A(B[17]), .B(A[17]), .Z(n34) );
  XOR2_X1 U32 ( .A(B[16]), .B(A[16]), .Z(n33) );
  XOR2_X1 U33 ( .A(B[15]), .B(A[15]), .Z(n32) );
  NOR4_X1 U34 ( .A1(n36), .A2(n37), .A3(n38), .A4(n39), .ZN(n30) );
  XOR2_X1 U35 ( .A(B[22]), .B(A[22]), .Z(n39) );
  XOR2_X1 U36 ( .A(B[21]), .B(A[21]), .Z(n38) );
  XOR2_X1 U37 ( .A(B[20]), .B(A[20]), .Z(n37) );
  XOR2_X1 U38 ( .A(B[19]), .B(A[19]), .Z(n36) );
  NOR4_X1 U39 ( .A1(n40), .A2(n41), .A3(n42), .A4(n43), .ZN(n29) );
  XOR2_X1 U40 ( .A(B[26]), .B(A[26]), .Z(n43) );
  XOR2_X1 U41 ( .A(B[25]), .B(A[25]), .Z(n42) );
  XOR2_X1 U42 ( .A(B[24]), .B(A[24]), .Z(n41) );
  XOR2_X1 U43 ( .A(B[23]), .B(A[23]), .Z(n40) );
  NOR4_X1 U44 ( .A1(n44), .A2(n45), .A3(n46), .A4(n47), .ZN(n28) );
  XOR2_X1 U45 ( .A(B[30]), .B(A[30]), .Z(n47) );
  XOR2_X1 U46 ( .A(B[29]), .B(A[29]), .Z(n46) );
  XOR2_X1 U47 ( .A(B[28]), .B(A[28]), .Z(n45) );
  XOR2_X1 U48 ( .A(B[27]), .B(A[27]), .Z(n44) );
endmodule


module cortexm0ds_logic_DW01_ash_1 ( A, DATA_TC, SH, SH_TC, B );
  input [30:0] A;
  input [4:0] SH;
  output [30:0] B;
  input DATA_TC, SH_TC;
  wire   \MR_int[1][30] , \ML_int[2][2] , \ML_int[3][6] , \ML_int[3][5] ,
         \ML_int[3][4] , \ML_int[3][2] , \ML_int[4][14] , \ML_int[4][13] ,
         \ML_int[4][12] , \ML_int[4][11] , \ML_int[4][10] , \ML_int[4][9] ,
         \ML_int[4][8] , \ML_int[5][30] , \ML_int[5][29] , \ML_int[5][28] ,
         \ML_int[5][27] , \ML_int[5][26] , \ML_int[5][25] , \ML_int[5][24] ,
         \ML_int[5][23] , \ML_int[5][22] , \ML_int[5][21] , \ML_int[5][20] ,
         \ML_int[5][19] , \ML_int[5][18] , \ML_int[5][17] , \ML_int[5][16] ,
         \ML_int[5][14] , \ML_int[5][13] , \ML_int[5][12] , \ML_int[5][11] ,
         \ML_int[5][10] , \ML_int[5][9] , \ML_int[5][8] , \ML_int[5][7] ,
         \ML_int[5][6] , \ML_int[5][5] , \ML_int[5][4] , \ML_int[5][3] ,
         \ML_int[5][2] , \ML_int[5][1] , \ML_int[5][0] , n1, n2, n3, n4, n5,
         n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n21,
         n22, n23, n24, n25, n26;
  assign \MR_int[1][30]  = SH[0];
  assign B[30] = \ML_int[5][30] ;
  assign B[29] = \ML_int[5][29] ;
  assign B[28] = \ML_int[5][28] ;
  assign B[27] = \ML_int[5][27] ;
  assign B[26] = \ML_int[5][26] ;
  assign B[25] = \ML_int[5][25] ;
  assign B[24] = \ML_int[5][24] ;
  assign B[23] = \ML_int[5][23] ;
  assign B[22] = \ML_int[5][22] ;
  assign B[21] = \ML_int[5][21] ;
  assign B[20] = \ML_int[5][20] ;
  assign B[19] = \ML_int[5][19] ;
  assign B[18] = \ML_int[5][18] ;
  assign B[17] = \ML_int[5][17] ;
  assign B[16] = \ML_int[5][16] ;
  assign B[14] = \ML_int[5][14] ;
  assign B[13] = \ML_int[5][13] ;
  assign B[12] = \ML_int[5][12] ;
  assign B[11] = \ML_int[5][11] ;
  assign B[10] = \ML_int[5][10] ;
  assign B[9] = \ML_int[5][9] ;
  assign B[8] = \ML_int[5][8] ;
  assign B[7] = \ML_int[5][7] ;
  assign B[6] = \ML_int[5][6] ;
  assign B[5] = \ML_int[5][5] ;
  assign B[4] = \ML_int[5][4] ;
  assign B[3] = \ML_int[5][3] ;
  assign B[2] = \ML_int[5][2] ;
  assign B[1] = \ML_int[5][1] ;
  assign B[0] = \ML_int[5][0] ;

  OR2_X1 U3 ( .A1(n2), .A2(SH[3]), .ZN(n1) );
  OR2_X1 U4 ( .A1(SH[1]), .A2(SH[2]), .ZN(n2) );
  OR2_X1 U5 ( .A1(SH[1]), .A2(\MR_int[1][30] ), .ZN(n3) );
  OR2_X1 U6 ( .A1(\MR_int[1][30] ), .A2(n2), .ZN(n4) );
  INV_X1 U7 ( .A(\ML_int[4][14] ), .ZN(n12) );
  INV_X1 U8 ( .A(\ML_int[4][10] ), .ZN(n8) );
  INV_X1 U9 ( .A(\ML_int[4][9] ), .ZN(n7) );
  INV_X1 U10 ( .A(\ML_int[4][8] ), .ZN(n6) );
  NAND2_X1 U11 ( .A1(SH[4]), .A2(n9), .ZN(\ML_int[5][27] ) );
  INV_X1 U12 ( .A(\ML_int[4][11] ), .ZN(n9) );
  NAND2_X1 U13 ( .A1(SH[4]), .A2(n10), .ZN(\ML_int[5][28] ) );
  INV_X1 U14 ( .A(\ML_int[4][12] ), .ZN(n10) );
  NAND2_X1 U15 ( .A1(SH[4]), .A2(n11), .ZN(\ML_int[5][29] ) );
  INV_X1 U16 ( .A(\ML_int[4][13] ), .ZN(n11) );
  INV_X1 U17 ( .A(SH[4]), .ZN(B[15]) );
  INV_X1 U18 ( .A(SH[3]), .ZN(n18) );
  NAND2_X1 U19 ( .A1(SH[3]), .A2(n15), .ZN(\ML_int[4][14] ) );
  INV_X1 U20 ( .A(\ML_int[3][6] ), .ZN(n15) );
  NAND2_X1 U21 ( .A1(SH[3]), .A2(n17), .ZN(\ML_int[4][13] ) );
  INV_X1 U22 ( .A(\ML_int[3][5] ), .ZN(n17) );
  NAND2_X1 U23 ( .A1(SH[3]), .A2(n14), .ZN(\ML_int[4][12] ) );
  INV_X1 U24 ( .A(\ML_int[3][4] ), .ZN(n14) );
  NAND2_X1 U25 ( .A1(SH[3]), .A2(SH[2]), .ZN(\ML_int[4][11] ) );
  NAND2_X1 U26 ( .A1(SH[3]), .A2(n16), .ZN(\ML_int[4][10] ) );
  INV_X1 U27 ( .A(\ML_int[3][2] ), .ZN(n16) );
  NAND2_X1 U28 ( .A1(SH[3]), .A2(n2), .ZN(\ML_int[4][9] ) );
  NAND2_X1 U29 ( .A1(SH[3]), .A2(n4), .ZN(\ML_int[4][8] ) );
  INV_X1 U30 ( .A(SH[2]), .ZN(n21) );
  NAND2_X1 U31 ( .A1(SH[2]), .A2(SH[1]), .ZN(\ML_int[3][5] ) );
  NAND2_X1 U32 ( .A1(SH[2]), .A2(n3), .ZN(\ML_int[3][4] ) );
  NAND2_X1 U33 ( .A1(SH[2]), .A2(n13), .ZN(\ML_int[3][6] ) );
  INV_X1 U34 ( .A(\ML_int[2][2] ), .ZN(n13) );
  NAND2_X1 U35 ( .A1(SH[1]), .A2(\MR_int[1][30] ), .ZN(\ML_int[2][2] ) );
  INV_X1 U36 ( .A(\MR_int[1][30] ), .ZN(n19) );
  OR2_X1 U37 ( .A1(\MR_int[1][30] ), .A2(n1), .ZN(n5) );
  NAND2_X1 U38 ( .A1(SH[4]), .A2(n7), .ZN(\ML_int[5][25] ) );
  NAND2_X1 U39 ( .A1(SH[4]), .A2(n22), .ZN(\ML_int[5][22] ) );
  NAND2_X1 U40 ( .A1(SH[4]), .A2(n8), .ZN(\ML_int[5][26] ) );
  NAND2_X1 U41 ( .A1(SH[4]), .A2(n6), .ZN(\ML_int[5][24] ) );
  NAND2_X1 U42 ( .A1(SH[4]), .A2(SH[3]), .ZN(\ML_int[5][23] ) );
  NAND2_X1 U43 ( .A1(SH[4]), .A2(n12), .ZN(\ML_int[5][30] ) );
  NAND2_X1 U44 ( .A1(SH[4]), .A2(n25), .ZN(\ML_int[5][19] ) );
  NAND2_X1 U45 ( .A1(SH[4]), .A2(n24), .ZN(\ML_int[5][20] ) );
  NAND2_X1 U46 ( .A1(SH[4]), .A2(n1), .ZN(\ML_int[5][17] ) );
  NAND2_X1 U47 ( .A1(SH[4]), .A2(n23), .ZN(\ML_int[5][21] ) );
  NAND2_X1 U48 ( .A1(SH[4]), .A2(n26), .ZN(\ML_int[5][18] ) );
  NAND2_X1 U49 ( .A1(SH[4]), .A2(n5), .ZN(\ML_int[5][16] ) );
  AND2_X1 U50 ( .A1(\ML_int[4][9] ), .A2(B[15]), .ZN(\ML_int[5][9] ) );
  AND2_X1 U51 ( .A1(\ML_int[4][8] ), .A2(B[15]), .ZN(\ML_int[5][8] ) );
  NOR2_X1 U52 ( .A1(SH[4]), .A2(SH[3]), .ZN(\ML_int[5][7] ) );
  NOR2_X1 U53 ( .A1(SH[4]), .A2(n22), .ZN(\ML_int[5][6] ) );
  NOR2_X1 U54 ( .A1(SH[4]), .A2(n23), .ZN(\ML_int[5][5] ) );
  NOR2_X1 U55 ( .A1(SH[4]), .A2(n24), .ZN(\ML_int[5][4] ) );
  NOR2_X1 U56 ( .A1(SH[4]), .A2(n25), .ZN(\ML_int[5][3] ) );
  NOR2_X1 U57 ( .A1(SH[4]), .A2(n26), .ZN(\ML_int[5][2] ) );
  AND2_X1 U58 ( .A1(\ML_int[4][14] ), .A2(B[15]), .ZN(\ML_int[5][14] ) );
  AND2_X1 U59 ( .A1(\ML_int[4][13] ), .A2(B[15]), .ZN(\ML_int[5][13] ) );
  AND2_X1 U60 ( .A1(\ML_int[4][12] ), .A2(B[15]), .ZN(\ML_int[5][12] ) );
  AND2_X1 U61 ( .A1(\ML_int[4][11] ), .A2(B[15]), .ZN(\ML_int[5][11] ) );
  AND2_X1 U62 ( .A1(\ML_int[4][10] ), .A2(B[15]), .ZN(\ML_int[5][10] ) );
  AND2_X1 U63 ( .A1(n19), .A2(\ML_int[5][1] ), .ZN(\ML_int[5][0] ) );
  NOR2_X1 U64 ( .A1(n1), .A2(SH[4]), .ZN(\ML_int[5][1] ) );
  NAND2_X1 U65 ( .A1(\ML_int[3][6] ), .A2(n18), .ZN(n22) );
  NAND2_X1 U66 ( .A1(\ML_int[3][5] ), .A2(n18), .ZN(n23) );
  NAND2_X1 U67 ( .A1(\ML_int[3][4] ), .A2(n18), .ZN(n24) );
  NAND2_X1 U68 ( .A1(n21), .A2(n18), .ZN(n25) );
  NAND2_X1 U69 ( .A1(\ML_int[3][2] ), .A2(n18), .ZN(n26) );
  AND2_X1 U70 ( .A1(\ML_int[2][2] ), .A2(n21), .ZN(\ML_int[3][2] ) );
endmodule


module cortexm0ds_logic_DW01_inc_1 ( A, SUM );
  input [29:0] A;
  output [29:0] SUM;

  wire   [29:2] carry;

  HA_X1 U1_1_28 ( .A(A[28]), .B(carry[28]), .CO(carry[29]), .S(SUM[28]) );
  HA_X1 U1_1_27 ( .A(A[27]), .B(carry[27]), .CO(carry[28]), .S(SUM[27]) );
  HA_X1 U1_1_26 ( .A(A[26]), .B(carry[26]), .CO(carry[27]), .S(SUM[26]) );
  HA_X1 U1_1_25 ( .A(A[25]), .B(carry[25]), .CO(carry[26]), .S(SUM[25]) );
  HA_X1 U1_1_24 ( .A(A[24]), .B(carry[24]), .CO(carry[25]), .S(SUM[24]) );
  HA_X1 U1_1_23 ( .A(A[23]), .B(carry[23]), .CO(carry[24]), .S(SUM[23]) );
  HA_X1 U1_1_22 ( .A(A[22]), .B(carry[22]), .CO(carry[23]), .S(SUM[22]) );
  HA_X1 U1_1_21 ( .A(A[21]), .B(carry[21]), .CO(carry[22]), .S(SUM[21]) );
  HA_X1 U1_1_20 ( .A(A[20]), .B(carry[20]), .CO(carry[21]), .S(SUM[20]) );
  HA_X1 U1_1_19 ( .A(A[19]), .B(carry[19]), .CO(carry[20]), .S(SUM[19]) );
  HA_X1 U1_1_18 ( .A(A[18]), .B(carry[18]), .CO(carry[19]), .S(SUM[18]) );
  HA_X1 U1_1_17 ( .A(A[17]), .B(carry[17]), .CO(carry[18]), .S(SUM[17]) );
  HA_X1 U1_1_16 ( .A(A[16]), .B(carry[16]), .CO(carry[17]), .S(SUM[16]) );
  HA_X1 U1_1_15 ( .A(A[15]), .B(carry[15]), .CO(carry[16]), .S(SUM[15]) );
  HA_X1 U1_1_14 ( .A(A[14]), .B(carry[14]), .CO(carry[15]), .S(SUM[14]) );
  HA_X1 U1_1_13 ( .A(A[13]), .B(carry[13]), .CO(carry[14]), .S(SUM[13]) );
  HA_X1 U1_1_12 ( .A(A[12]), .B(carry[12]), .CO(carry[13]), .S(SUM[12]) );
  HA_X1 U1_1_11 ( .A(A[11]), .B(carry[11]), .CO(carry[12]), .S(SUM[11]) );
  HA_X1 U1_1_10 ( .A(A[10]), .B(carry[10]), .CO(carry[11]), .S(SUM[10]) );
  HA_X1 U1_1_9 ( .A(A[9]), .B(carry[9]), .CO(carry[10]), .S(SUM[9]) );
  HA_X1 U1_1_8 ( .A(A[8]), .B(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  HA_X1 U1_1_7 ( .A(A[7]), .B(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  HA_X1 U1_1_6 ( .A(A[6]), .B(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  HA_X1 U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  HA_X1 U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  HA_X1 U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  HA_X1 U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  HA_X1 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .S(SUM[1]) );
  XOR2_X1 U1 ( .A(carry[29]), .B(A[29]), .Z(SUM[29]) );
endmodule


module cortexm0ds_logic_DW01_add_3 ( A, B, CI, SUM, CO );
  input [33:0] A;
  input [33:0] B;
  output [33:0] SUM;
  input CI;
  output CO;
  wire   n1;
  wire   [33:1] carry;

  FA_X1 U1_32 ( .A(A[32]), .B(B[32]), .CI(carry[32]), .CO(SUM[33]), .S(SUM[32]) );
  FA_X1 U1_31 ( .A(A[31]), .B(B[31]), .CI(carry[31]), .CO(carry[32]), .S(
        SUM[31]) );
  FA_X1 U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  FA_X1 U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  FA_X1 U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  FA_X1 U1_27 ( .A(A[27]), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  FA_X1 U1_26 ( .A(A[26]), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  FA_X1 U1_25 ( .A(A[25]), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  FA_X1 U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  FA_X1 U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  FA_X1 U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  FA_X1 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  FA_X1 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  FA_X1 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  FA_X1 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  FA_X1 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  FA_X1 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  FA_X1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  FA_X1 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  FA_X1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  FA_X1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  FA_X1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  FA_X1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  FA_X1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  FA_X1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  FA_X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  FA_X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  FA_X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  FA_X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  FA_X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  FA_X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(n1), .CO(carry[3]), .S(SUM[2]) );
  AND2_X1 U1 ( .A1(B[1]), .A2(A[1]), .ZN(n1) );
  XOR2_X1 U2 ( .A(B[1]), .B(A[1]), .Z(SUM[1]) );
endmodule


module cortexm0ds_logic_DW01_add_2 ( A, B, CI, SUM, CO );
  input [33:0] A;
  input [33:0] B;
  output [33:0] SUM;
  input CI;
  output CO;
  wire   n3, n4, n5, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21,
         n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35,
         n37, n61, n62, n65;

  XOR2_X1 U1 ( .A(A[28]), .B(n4), .Z(SUM[28]) );
  XOR2_X1 U2 ( .A(A[32]), .B(n35), .Z(SUM[32]) );
  AND2_X1 U3 ( .A1(A[26]), .A2(n32), .ZN(n3) );
  AND2_X1 U4 ( .A1(A[27]), .A2(n3), .ZN(n4) );
  AND2_X1 U5 ( .A1(A[28]), .A2(n4), .ZN(n5) );
  XOR2_X1 U6 ( .A(A[26]), .B(n32), .Z(SUM[26]) );
  XOR2_X1 U7 ( .A(A[27]), .B(n3), .Z(SUM[27]) );
  XNOR2_X1 U8 ( .A(A[33]), .B(n65), .ZN(SUM[33]) );
  NAND2_X1 U9 ( .A1(A[32]), .A2(n35), .ZN(n65) );
  XOR2_X1 U10 ( .A(A[29]), .B(n5), .Z(SUM[29]) );
  XOR2_X1 U11 ( .A(A[30]), .B(n33), .Z(SUM[30]) );
  AND2_X1 U12 ( .A1(A[18]), .A2(n25), .ZN(n11) );
  AND2_X1 U13 ( .A1(A[4]), .A2(n62), .ZN(n12) );
  AND2_X1 U14 ( .A1(A[5]), .A2(n12), .ZN(n13) );
  AND2_X1 U15 ( .A1(A[6]), .A2(n13), .ZN(n14) );
  AND2_X1 U16 ( .A1(A[7]), .A2(n14), .ZN(n15) );
  AND2_X1 U17 ( .A1(A[8]), .A2(n15), .ZN(n16) );
  AND2_X1 U18 ( .A1(A[9]), .A2(n16), .ZN(n17) );
  AND2_X1 U19 ( .A1(A[10]), .A2(n17), .ZN(n18) );
  AND2_X1 U20 ( .A1(A[11]), .A2(n18), .ZN(n19) );
  AND2_X1 U21 ( .A1(A[12]), .A2(n19), .ZN(n20) );
  AND2_X1 U22 ( .A1(A[13]), .A2(n20), .ZN(n21) );
  AND2_X1 U23 ( .A1(A[14]), .A2(n21), .ZN(n22) );
  AND2_X1 U24 ( .A1(A[15]), .A2(n22), .ZN(n23) );
  AND2_X1 U25 ( .A1(A[16]), .A2(n23), .ZN(n24) );
  AND2_X1 U26 ( .A1(A[17]), .A2(n24), .ZN(n25) );
  AND2_X1 U27 ( .A1(A[19]), .A2(n11), .ZN(n26) );
  AND2_X1 U28 ( .A1(A[20]), .A2(n26), .ZN(n27) );
  AND2_X1 U29 ( .A1(A[21]), .A2(n27), .ZN(n28) );
  AND2_X1 U30 ( .A1(A[22]), .A2(n28), .ZN(n29) );
  AND2_X1 U31 ( .A1(A[23]), .A2(n29), .ZN(n30) );
  AND2_X1 U32 ( .A1(A[24]), .A2(n30), .ZN(n31) );
  AND2_X1 U33 ( .A1(A[25]), .A2(n31), .ZN(n32) );
  AND2_X1 U34 ( .A1(A[29]), .A2(n5), .ZN(n33) );
  AND2_X1 U35 ( .A1(A[30]), .A2(n33), .ZN(n34) );
  AND2_X1 U36 ( .A1(A[31]), .A2(n34), .ZN(n35) );
  XOR2_X1 U37 ( .A(A[31]), .B(n34), .Z(SUM[31]) );
  AND2_X1 U38 ( .A1(A[2]), .A2(n61), .ZN(n37) );
  XOR2_X1 U39 ( .A(A[25]), .B(n31), .Z(SUM[25]) );
  XOR2_X1 U40 ( .A(A[20]), .B(n26), .Z(SUM[20]) );
  XOR2_X1 U41 ( .A(A[19]), .B(n11), .Z(SUM[19]) );
  XOR2_X1 U42 ( .A(A[18]), .B(n25), .Z(SUM[18]) );
  XOR2_X1 U43 ( .A(A[17]), .B(n24), .Z(SUM[17]) );
  XOR2_X1 U44 ( .A(A[23]), .B(n29), .Z(SUM[23]) );
  XOR2_X1 U45 ( .A(A[22]), .B(n28), .Z(SUM[22]) );
  XOR2_X1 U46 ( .A(A[21]), .B(n27), .Z(SUM[21]) );
  XOR2_X1 U47 ( .A(A[24]), .B(n30), .Z(SUM[24]) );
  XOR2_X1 U48 ( .A(A[16]), .B(n23), .Z(SUM[16]) );
  XOR2_X1 U49 ( .A(A[5]), .B(n12), .Z(SUM[5]) );
  XOR2_X1 U50 ( .A(A[2]), .B(n61), .Z(SUM[2]) );
  XOR2_X1 U51 ( .A(A[13]), .B(n20), .Z(SUM[13]) );
  XOR2_X1 U52 ( .A(A[12]), .B(n19), .Z(SUM[12]) );
  XOR2_X1 U53 ( .A(A[11]), .B(n18), .Z(SUM[11]) );
  XOR2_X1 U54 ( .A(A[10]), .B(n17), .Z(SUM[10]) );
  XOR2_X1 U55 ( .A(A[15]), .B(n22), .Z(SUM[15]) );
  XOR2_X1 U56 ( .A(A[14]), .B(n21), .Z(SUM[14]) );
  XOR2_X1 U57 ( .A(A[9]), .B(n16), .Z(SUM[9]) );
  XOR2_X1 U58 ( .A(A[8]), .B(n15), .Z(SUM[8]) );
  XOR2_X1 U59 ( .A(A[7]), .B(n14), .Z(SUM[7]) );
  XOR2_X1 U60 ( .A(A[4]), .B(n62), .Z(SUM[4]) );
  XOR2_X1 U61 ( .A(A[6]), .B(n13), .Z(SUM[6]) );
  AND2_X1 U62 ( .A1(B[1]), .A2(A[1]), .ZN(n61) );
  AND2_X1 U63 ( .A1(A[3]), .A2(n37), .ZN(n62) );
  XOR2_X1 U64 ( .A(A[3]), .B(n37), .Z(SUM[3]) );
  XOR2_X1 U65 ( .A(B[1]), .B(A[1]), .Z(SUM[1]) );
endmodule


module cortexm0ds_logic_DW02_mult_0 ( A, B, TC, PRODUCT );
  input [31:0] A;
  input [31:0] B;
  output [63:0] PRODUCT;
  input TC;
  wire   \ab[31][0] , \ab[30][1] , \ab[30][0] , \ab[29][2] , \ab[29][1] ,
         \ab[29][0] , \ab[28][3] , \ab[28][2] , \ab[28][1] , \ab[28][0] ,
         \ab[27][4] , \ab[27][3] , \ab[27][2] , \ab[27][1] , \ab[27][0] ,
         \ab[26][5] , \ab[26][4] , \ab[26][3] , \ab[26][2] , \ab[26][1] ,
         \ab[26][0] , \ab[25][6] , \ab[25][5] , \ab[25][4] , \ab[25][3] ,
         \ab[25][2] , \ab[25][1] , \ab[25][0] , \ab[24][7] , \ab[24][6] ,
         \ab[24][5] , \ab[24][4] , \ab[24][3] , \ab[24][2] , \ab[24][1] ,
         \ab[24][0] , \ab[23][8] , \ab[23][7] , \ab[23][6] , \ab[23][5] ,
         \ab[23][4] , \ab[23][3] , \ab[23][2] , \ab[23][1] , \ab[23][0] ,
         \ab[22][9] , \ab[22][8] , \ab[22][7] , \ab[22][6] , \ab[22][5] ,
         \ab[22][4] , \ab[22][3] , \ab[22][2] , \ab[22][1] , \ab[22][0] ,
         \ab[21][10] , \ab[21][9] , \ab[21][8] , \ab[21][7] , \ab[21][6] ,
         \ab[21][5] , \ab[21][4] , \ab[21][3] , \ab[21][2] , \ab[21][1] ,
         \ab[21][0] , \ab[20][11] , \ab[20][10] , \ab[20][9] , \ab[20][8] ,
         \ab[20][7] , \ab[20][6] , \ab[20][5] , \ab[20][4] , \ab[20][3] ,
         \ab[20][2] , \ab[20][1] , \ab[20][0] , \ab[19][12] , \ab[19][11] ,
         \ab[19][10] , \ab[19][9] , \ab[19][8] , \ab[19][7] , \ab[19][6] ,
         \ab[19][5] , \ab[19][4] , \ab[19][3] , \ab[19][2] , \ab[19][1] ,
         \ab[19][0] , \ab[18][13] , \ab[18][12] , \ab[18][11] , \ab[18][10] ,
         \ab[18][9] , \ab[18][8] , \ab[18][7] , \ab[18][6] , \ab[18][5] ,
         \ab[18][4] , \ab[18][3] , \ab[18][2] , \ab[18][1] , \ab[18][0] ,
         \ab[17][14] , \ab[17][13] , \ab[17][12] , \ab[17][11] , \ab[17][10] ,
         \ab[17][9] , \ab[17][8] , \ab[17][7] , \ab[17][6] , \ab[17][5] ,
         \ab[17][4] , \ab[17][3] , \ab[17][2] , \ab[17][1] , \ab[17][0] ,
         \ab[16][15] , \ab[16][14] , \ab[16][13] , \ab[16][12] , \ab[16][11] ,
         \ab[16][10] , \ab[16][9] , \ab[16][8] , \ab[16][7] , \ab[16][6] ,
         \ab[16][5] , \ab[16][4] , \ab[16][3] , \ab[16][2] , \ab[16][1] ,
         \ab[16][0] , \ab[15][16] , \ab[15][15] , \ab[15][14] , \ab[15][13] ,
         \ab[15][12] , \ab[15][11] , \ab[15][10] , \ab[15][9] , \ab[15][8] ,
         \ab[15][7] , \ab[15][6] , \ab[15][5] , \ab[15][4] , \ab[15][3] ,
         \ab[15][2] , \ab[15][1] , \ab[15][0] , \ab[14][17] , \ab[14][16] ,
         \ab[14][15] , \ab[14][14] , \ab[14][13] , \ab[14][12] , \ab[14][11] ,
         \ab[14][10] , \ab[14][9] , \ab[14][8] , \ab[14][7] , \ab[14][6] ,
         \ab[14][5] , \ab[14][4] , \ab[14][3] , \ab[14][2] , \ab[14][1] ,
         \ab[14][0] , \ab[13][18] , \ab[13][17] , \ab[13][16] , \ab[13][15] ,
         \ab[13][14] , \ab[13][13] , \ab[13][12] , \ab[13][11] , \ab[13][10] ,
         \ab[13][9] , \ab[13][8] , \ab[13][7] , \ab[13][6] , \ab[13][5] ,
         \ab[13][4] , \ab[13][3] , \ab[13][2] , \ab[13][1] , \ab[13][0] ,
         \ab[12][19] , \ab[12][18] , \ab[12][17] , \ab[12][16] , \ab[12][15] ,
         \ab[12][14] , \ab[12][13] , \ab[12][12] , \ab[12][11] , \ab[12][10] ,
         \ab[12][9] , \ab[12][8] , \ab[12][7] , \ab[12][6] , \ab[12][5] ,
         \ab[12][4] , \ab[12][3] , \ab[12][2] , \ab[12][1] , \ab[12][0] ,
         \ab[11][20] , \ab[11][19] , \ab[11][18] , \ab[11][17] , \ab[11][16] ,
         \ab[11][15] , \ab[11][14] , \ab[11][13] , \ab[11][12] , \ab[11][11] ,
         \ab[11][10] , \ab[11][9] , \ab[11][8] , \ab[11][7] , \ab[11][6] ,
         \ab[11][5] , \ab[11][4] , \ab[11][3] , \ab[11][2] , \ab[11][1] ,
         \ab[11][0] , \ab[10][21] , \ab[10][20] , \ab[10][19] , \ab[10][18] ,
         \ab[10][17] , \ab[10][16] , \ab[10][15] , \ab[10][14] , \ab[10][13] ,
         \ab[10][12] , \ab[10][11] , \ab[10][10] , \ab[10][9] , \ab[10][8] ,
         \ab[10][7] , \ab[10][6] , \ab[10][5] , \ab[10][4] , \ab[10][3] ,
         \ab[10][2] , \ab[10][1] , \ab[10][0] , \ab[9][22] , \ab[9][21] ,
         \ab[9][20] , \ab[9][19] , \ab[9][18] , \ab[9][17] , \ab[9][16] ,
         \ab[9][15] , \ab[9][14] , \ab[9][13] , \ab[9][12] , \ab[9][11] ,
         \ab[9][10] , \ab[9][9] , \ab[9][8] , \ab[9][7] , \ab[9][6] ,
         \ab[9][5] , \ab[9][4] , \ab[9][3] , \ab[9][2] , \ab[9][1] ,
         \ab[9][0] , \ab[8][23] , \ab[8][22] , \ab[8][21] , \ab[8][20] ,
         \ab[8][19] , \ab[8][18] , \ab[8][17] , \ab[8][16] , \ab[8][15] ,
         \ab[8][14] , \ab[8][13] , \ab[8][12] , \ab[8][11] , \ab[8][10] ,
         \ab[8][9] , \ab[8][8] , \ab[8][7] , \ab[8][6] , \ab[8][5] ,
         \ab[8][4] , \ab[8][3] , \ab[8][2] , \ab[8][1] , \ab[8][0] ,
         \ab[7][24] , \ab[7][23] , \ab[7][22] , \ab[7][21] , \ab[7][20] ,
         \ab[7][19] , \ab[7][18] , \ab[7][17] , \ab[7][16] , \ab[7][15] ,
         \ab[7][14] , \ab[7][13] , \ab[7][12] , \ab[7][11] , \ab[7][10] ,
         \ab[7][9] , \ab[7][8] , \ab[7][7] , \ab[7][6] , \ab[7][5] ,
         \ab[7][4] , \ab[7][3] , \ab[7][2] , \ab[7][1] , \ab[7][0] ,
         \ab[6][25] , \ab[6][24] , \ab[6][23] , \ab[6][22] , \ab[6][21] ,
         \ab[6][20] , \ab[6][19] , \ab[6][18] , \ab[6][17] , \ab[6][16] ,
         \ab[6][15] , \ab[6][14] , \ab[6][13] , \ab[6][12] , \ab[6][11] ,
         \ab[6][10] , \ab[6][9] , \ab[6][8] , \ab[6][7] , \ab[6][6] ,
         \ab[6][5] , \ab[6][4] , \ab[6][3] , \ab[6][2] , \ab[6][1] ,
         \ab[6][0] , \ab[5][26] , \ab[5][25] , \ab[5][24] , \ab[5][23] ,
         \ab[5][22] , \ab[5][21] , \ab[5][20] , \ab[5][19] , \ab[5][18] ,
         \ab[5][17] , \ab[5][16] , \ab[5][15] , \ab[5][14] , \ab[5][13] ,
         \ab[5][12] , \ab[5][11] , \ab[5][10] , \ab[5][9] , \ab[5][8] ,
         \ab[5][7] , \ab[5][6] , \ab[5][5] , \ab[5][4] , \ab[5][3] ,
         \ab[5][2] , \ab[5][1] , \ab[5][0] , \ab[4][27] , \ab[4][26] ,
         \ab[4][25] , \ab[4][24] , \ab[4][23] , \ab[4][22] , \ab[4][21] ,
         \ab[4][20] , \ab[4][19] , \ab[4][18] , \ab[4][17] , \ab[4][16] ,
         \ab[4][15] , \ab[4][14] , \ab[4][13] , \ab[4][12] , \ab[4][11] ,
         \ab[4][10] , \ab[4][9] , \ab[4][8] , \ab[4][7] , \ab[4][6] ,
         \ab[4][5] , \ab[4][4] , \ab[4][3] , \ab[4][2] , \ab[4][1] ,
         \ab[4][0] , \ab[3][28] , \ab[3][27] , \ab[3][26] , \ab[3][25] ,
         \ab[3][24] , \ab[3][23] , \ab[3][22] , \ab[3][21] , \ab[3][20] ,
         \ab[3][19] , \ab[3][18] , \ab[3][17] , \ab[3][16] , \ab[3][15] ,
         \ab[3][14] , \ab[3][13] , \ab[3][12] , \ab[3][11] , \ab[3][10] ,
         \ab[3][9] , \ab[3][8] , \ab[3][7] , \ab[3][6] , \ab[3][5] ,
         \ab[3][4] , \ab[3][3] , \ab[3][2] , \ab[3][1] , \ab[3][0] ,
         \ab[2][29] , \ab[2][28] , \ab[2][27] , \ab[2][26] , \ab[2][25] ,
         \ab[2][24] , \ab[2][23] , \ab[2][22] , \ab[2][21] , \ab[2][20] ,
         \ab[2][19] , \ab[2][18] , \ab[2][17] , \ab[2][16] , \ab[2][15] ,
         \ab[2][14] , \ab[2][13] , \ab[2][12] , \ab[2][11] , \ab[2][10] ,
         \ab[2][9] , \ab[2][8] , \ab[2][7] , \ab[2][6] , \ab[2][5] ,
         \ab[2][4] , \ab[2][3] , \ab[2][2] , \ab[2][1] , \ab[2][0] ,
         \ab[1][30] , \ab[1][29] , \ab[1][28] , \ab[1][27] , \ab[1][26] ,
         \ab[1][25] , \ab[1][24] , \ab[1][23] , \ab[1][22] , \ab[1][21] ,
         \ab[1][20] , \ab[1][19] , \ab[1][18] , \ab[1][17] , \ab[1][16] ,
         \ab[1][15] , \ab[1][14] , \ab[1][13] , \ab[1][12] , \ab[1][11] ,
         \ab[1][10] , \ab[1][9] , \ab[1][8] , \ab[1][7] , \ab[1][6] ,
         \ab[1][5] , \ab[1][4] , \ab[1][3] , \ab[1][2] , \ab[1][1] ,
         \ab[1][0] , \ab[0][31] , \ab[0][30] , \ab[0][29] , \ab[0][28] ,
         \ab[0][27] , \ab[0][26] , \ab[0][25] , \ab[0][24] , \ab[0][23] ,
         \ab[0][22] , \ab[0][21] , \ab[0][20] , \ab[0][19] , \ab[0][18] ,
         \ab[0][17] , \ab[0][16] , \ab[0][15] , \ab[0][14] , \ab[0][13] ,
         \ab[0][12] , \ab[0][11] , \ab[0][10] , \ab[0][9] , \ab[0][8] ,
         \ab[0][7] , \ab[0][6] , \ab[0][5] , \ab[0][4] , \ab[0][3] ,
         \ab[0][2] , \ab[0][1] , \CARRYB[15][15] , \CARRYB[15][14] ,
         \CARRYB[15][13] , \CARRYB[15][12] , \CARRYB[15][11] ,
         \CARRYB[15][10] , \CARRYB[15][9] , \CARRYB[15][8] , \CARRYB[15][7] ,
         \CARRYB[15][6] , \CARRYB[15][5] , \CARRYB[15][4] , \CARRYB[15][3] ,
         \CARRYB[15][2] , \CARRYB[15][1] , \CARRYB[15][0] , \CARRYB[14][16] ,
         \CARRYB[14][15] , \CARRYB[14][14] , \CARRYB[14][13] ,
         \CARRYB[14][12] , \CARRYB[14][11] , \CARRYB[14][10] , \CARRYB[14][9] ,
         \CARRYB[14][8] , \CARRYB[14][7] , \CARRYB[14][6] , \CARRYB[14][5] ,
         \CARRYB[14][4] , \CARRYB[14][3] , \CARRYB[14][2] , \CARRYB[14][1] ,
         \CARRYB[14][0] , \CARRYB[13][17] , \CARRYB[13][16] , \CARRYB[13][15] ,
         \CARRYB[13][14] , \CARRYB[13][13] , \CARRYB[13][12] ,
         \CARRYB[13][11] , \CARRYB[13][10] , \CARRYB[13][9] , \CARRYB[13][8] ,
         \CARRYB[13][7] , \CARRYB[13][6] , \CARRYB[13][5] , \CARRYB[13][4] ,
         \CARRYB[13][3] , \CARRYB[13][2] , \CARRYB[13][1] , \CARRYB[13][0] ,
         \CARRYB[12][18] , \CARRYB[12][17] , \CARRYB[12][16] ,
         \CARRYB[12][15] , \CARRYB[12][14] , \CARRYB[12][13] ,
         \CARRYB[12][12] , \CARRYB[12][11] , \CARRYB[12][10] , \CARRYB[12][9] ,
         \CARRYB[12][8] , \CARRYB[12][7] , \CARRYB[12][6] , \CARRYB[12][5] ,
         \CARRYB[12][4] , \CARRYB[12][3] , \CARRYB[12][2] , \CARRYB[12][1] ,
         \CARRYB[12][0] , \CARRYB[11][19] , \CARRYB[11][18] , \CARRYB[11][17] ,
         \CARRYB[11][16] , \CARRYB[11][15] , \CARRYB[11][14] ,
         \CARRYB[11][13] , \CARRYB[11][12] , \CARRYB[11][11] ,
         \CARRYB[11][10] , \CARRYB[11][9] , \CARRYB[11][8] , \CARRYB[11][7] ,
         \CARRYB[11][6] , \CARRYB[11][5] , \CARRYB[11][4] , \CARRYB[11][3] ,
         \CARRYB[11][2] , \CARRYB[11][1] , \CARRYB[11][0] , \CARRYB[10][20] ,
         \CARRYB[10][19] , \CARRYB[10][18] , \CARRYB[10][17] ,
         \CARRYB[10][16] , \CARRYB[10][15] , \CARRYB[10][14] ,
         \CARRYB[10][13] , \CARRYB[10][12] , \CARRYB[10][11] ,
         \CARRYB[10][10] , \CARRYB[10][9] , \CARRYB[10][8] , \CARRYB[10][7] ,
         \CARRYB[10][6] , \CARRYB[10][5] , \CARRYB[10][4] , \CARRYB[10][3] ,
         \CARRYB[10][2] , \CARRYB[10][1] , \CARRYB[10][0] , \CARRYB[9][21] ,
         \CARRYB[9][20] , \CARRYB[9][19] , \CARRYB[9][18] , \CARRYB[9][17] ,
         \CARRYB[9][16] , \CARRYB[9][15] , \CARRYB[9][14] , \CARRYB[9][13] ,
         \CARRYB[9][12] , \CARRYB[9][11] , \CARRYB[9][10] , \CARRYB[9][9] ,
         \CARRYB[9][8] , \CARRYB[9][7] , \CARRYB[9][6] , \CARRYB[9][5] ,
         \CARRYB[9][4] , \CARRYB[9][3] , \CARRYB[9][2] , \CARRYB[9][1] ,
         \CARRYB[9][0] , \CARRYB[8][22] , \CARRYB[8][21] , \CARRYB[8][20] ,
         \CARRYB[8][19] , \CARRYB[8][18] , \CARRYB[8][17] , \CARRYB[8][16] ,
         \CARRYB[8][15] , \CARRYB[8][14] , \CARRYB[8][13] , \CARRYB[8][12] ,
         \CARRYB[8][11] , \CARRYB[8][10] , \CARRYB[8][9] , \CARRYB[8][8] ,
         \CARRYB[8][7] , \CARRYB[8][6] , \CARRYB[8][5] , \CARRYB[8][4] ,
         \CARRYB[8][3] , \CARRYB[8][2] , \CARRYB[8][1] , \CARRYB[8][0] ,
         \CARRYB[7][23] , \CARRYB[7][22] , \CARRYB[7][21] , \CARRYB[7][20] ,
         \CARRYB[7][19] , \CARRYB[7][18] , \CARRYB[7][17] , \CARRYB[7][16] ,
         \CARRYB[7][15] , \CARRYB[7][14] , \CARRYB[7][13] , \CARRYB[7][12] ,
         \CARRYB[7][11] , \CARRYB[7][10] , \CARRYB[7][9] , \CARRYB[7][8] ,
         \CARRYB[7][7] , \CARRYB[7][6] , \CARRYB[7][5] , \CARRYB[7][4] ,
         \CARRYB[7][3] , \CARRYB[7][2] , \CARRYB[7][1] , \CARRYB[7][0] ,
         \CARRYB[6][24] , \CARRYB[6][23] , \CARRYB[6][22] , \CARRYB[6][21] ,
         \CARRYB[6][20] , \CARRYB[6][19] , \CARRYB[6][18] , \CARRYB[6][17] ,
         \CARRYB[6][16] , \CARRYB[6][15] , \CARRYB[6][14] , \CARRYB[6][13] ,
         \CARRYB[6][12] , \CARRYB[6][11] , \CARRYB[6][10] , \CARRYB[6][9] ,
         \CARRYB[6][8] , \CARRYB[6][7] , \CARRYB[6][6] , \CARRYB[6][5] ,
         \CARRYB[6][4] , \CARRYB[6][3] , \CARRYB[6][2] , \CARRYB[6][1] ,
         \CARRYB[6][0] , \CARRYB[5][25] , \CARRYB[5][24] , \CARRYB[5][23] ,
         \CARRYB[5][22] , \CARRYB[5][21] , \CARRYB[5][20] , \CARRYB[5][19] ,
         \CARRYB[5][18] , \CARRYB[5][17] , \CARRYB[5][16] , \CARRYB[5][15] ,
         \CARRYB[5][14] , \CARRYB[5][13] , \CARRYB[5][12] , \CARRYB[5][11] ,
         \CARRYB[5][10] , \CARRYB[5][9] , \CARRYB[5][8] , \CARRYB[5][7] ,
         \CARRYB[5][6] , \CARRYB[5][5] , \CARRYB[5][4] , \CARRYB[5][3] ,
         \CARRYB[5][2] , \CARRYB[5][1] , \CARRYB[5][0] , \CARRYB[4][26] ,
         \CARRYB[4][25] , \CARRYB[4][24] , \CARRYB[4][23] , \CARRYB[4][22] ,
         \CARRYB[4][21] , \CARRYB[4][20] , \CARRYB[4][19] , \CARRYB[4][18] ,
         \CARRYB[4][17] , \CARRYB[4][16] , \CARRYB[4][15] , \CARRYB[4][14] ,
         \CARRYB[4][13] , \CARRYB[4][12] , \CARRYB[4][11] , \CARRYB[4][10] ,
         \CARRYB[4][9] , \CARRYB[4][8] , \CARRYB[4][7] , \CARRYB[4][6] ,
         \CARRYB[4][5] , \CARRYB[4][4] , \CARRYB[4][3] , \CARRYB[4][2] ,
         \CARRYB[4][1] , \CARRYB[4][0] , \CARRYB[3][27] , \CARRYB[3][26] ,
         \CARRYB[3][25] , \CARRYB[3][24] , \CARRYB[3][23] , \CARRYB[3][22] ,
         \CARRYB[3][21] , \CARRYB[3][20] , \CARRYB[3][19] , \CARRYB[3][18] ,
         \CARRYB[3][17] , \CARRYB[3][16] , \CARRYB[3][15] , \CARRYB[3][14] ,
         \CARRYB[3][13] , \CARRYB[3][12] , \CARRYB[3][11] , \CARRYB[3][10] ,
         \CARRYB[3][9] , \CARRYB[3][8] , \CARRYB[3][7] , \CARRYB[3][6] ,
         \CARRYB[3][5] , \CARRYB[3][4] , \CARRYB[3][3] , \CARRYB[3][2] ,
         \CARRYB[3][1] , \CARRYB[3][0] , \CARRYB[2][28] , \CARRYB[2][27] ,
         \CARRYB[2][26] , \CARRYB[2][25] , \CARRYB[2][24] , \CARRYB[2][23] ,
         \CARRYB[2][22] , \CARRYB[2][21] , \CARRYB[2][20] , \CARRYB[2][19] ,
         \CARRYB[2][18] , \CARRYB[2][17] , \CARRYB[2][16] , \CARRYB[2][15] ,
         \CARRYB[2][14] , \CARRYB[2][13] , \CARRYB[2][12] , \CARRYB[2][11] ,
         \CARRYB[2][10] , \CARRYB[2][9] , \CARRYB[2][8] , \CARRYB[2][7] ,
         \CARRYB[2][6] , \CARRYB[2][5] , \CARRYB[2][4] , \CARRYB[2][3] ,
         \CARRYB[2][2] , \CARRYB[2][1] , \CARRYB[2][0] , \SUMB[15][16] ,
         \SUMB[15][15] , \SUMB[15][14] , \SUMB[15][13] , \SUMB[15][12] ,
         \SUMB[15][11] , \SUMB[15][10] , \SUMB[15][9] , \SUMB[15][8] ,
         \SUMB[15][7] , \SUMB[15][6] , \SUMB[15][5] , \SUMB[15][4] ,
         \SUMB[15][3] , \SUMB[15][2] , \SUMB[15][1] , \SUMB[14][17] ,
         \SUMB[14][16] , \SUMB[14][15] , \SUMB[14][14] , \SUMB[14][13] ,
         \SUMB[14][12] , \SUMB[14][11] , \SUMB[14][10] , \SUMB[14][9] ,
         \SUMB[14][8] , \SUMB[14][7] , \SUMB[14][6] , \SUMB[14][5] ,
         \SUMB[14][4] , \SUMB[14][3] , \SUMB[14][2] , \SUMB[14][1] ,
         \SUMB[13][18] , \SUMB[13][17] , \SUMB[13][16] , \SUMB[13][15] ,
         \SUMB[13][14] , \SUMB[13][13] , \SUMB[13][12] , \SUMB[13][11] ,
         \SUMB[13][10] , \SUMB[13][9] , \SUMB[13][8] , \SUMB[13][7] ,
         \SUMB[13][6] , \SUMB[13][5] , \SUMB[13][4] , \SUMB[13][3] ,
         \SUMB[13][2] , \SUMB[13][1] , \SUMB[12][19] , \SUMB[12][18] ,
         \SUMB[12][17] , \SUMB[12][16] , \SUMB[12][15] , \SUMB[12][14] ,
         \SUMB[12][13] , \SUMB[12][12] , \SUMB[12][11] , \SUMB[12][10] ,
         \SUMB[12][9] , \SUMB[12][8] , \SUMB[12][7] , \SUMB[12][6] ,
         \SUMB[12][5] , \SUMB[12][4] , \SUMB[12][3] , \SUMB[12][2] ,
         \SUMB[12][1] , \SUMB[11][20] , \SUMB[11][19] , \SUMB[11][18] ,
         \SUMB[11][17] , \SUMB[11][16] , \SUMB[11][15] , \SUMB[11][14] ,
         \SUMB[11][13] , \SUMB[11][12] , \SUMB[11][11] , \SUMB[11][10] ,
         \SUMB[11][9] , \SUMB[11][8] , \SUMB[11][7] , \SUMB[11][6] ,
         \SUMB[11][5] , \SUMB[11][4] , \SUMB[11][3] , \SUMB[11][2] ,
         \SUMB[11][1] , \SUMB[10][21] , \SUMB[10][20] , \SUMB[10][19] ,
         \SUMB[10][18] , \SUMB[10][17] , \SUMB[10][16] , \SUMB[10][15] ,
         \SUMB[10][14] , \SUMB[10][13] , \SUMB[10][12] , \SUMB[10][11] ,
         \SUMB[10][10] , \SUMB[10][9] , \SUMB[10][8] , \SUMB[10][7] ,
         \SUMB[10][6] , \SUMB[10][5] , \SUMB[10][4] , \SUMB[10][3] ,
         \SUMB[10][2] , \SUMB[10][1] , \SUMB[9][22] , \SUMB[9][21] ,
         \SUMB[9][20] , \SUMB[9][19] , \SUMB[9][18] , \SUMB[9][17] ,
         \SUMB[9][16] , \SUMB[9][15] , \SUMB[9][14] , \SUMB[9][13] ,
         \SUMB[9][12] , \SUMB[9][11] , \SUMB[9][10] , \SUMB[9][9] ,
         \SUMB[9][8] , \SUMB[9][7] , \SUMB[9][6] , \SUMB[9][5] , \SUMB[9][4] ,
         \SUMB[9][3] , \SUMB[9][2] , \SUMB[9][1] , \SUMB[8][23] ,
         \SUMB[8][22] , \SUMB[8][21] , \SUMB[8][20] , \SUMB[8][19] ,
         \SUMB[8][18] , \SUMB[8][17] , \SUMB[8][16] , \SUMB[8][15] ,
         \SUMB[8][14] , \SUMB[8][13] , \SUMB[8][12] , \SUMB[8][11] ,
         \SUMB[8][10] , \SUMB[8][9] , \SUMB[8][8] , \SUMB[8][7] , \SUMB[8][6] ,
         \SUMB[8][5] , \SUMB[8][4] , \SUMB[8][3] , \SUMB[8][2] , \SUMB[8][1] ,
         \SUMB[7][24] , \SUMB[7][23] , \SUMB[7][22] , \SUMB[7][21] ,
         \SUMB[7][20] , \SUMB[7][19] , \SUMB[7][18] , \SUMB[7][17] ,
         \SUMB[7][16] , \SUMB[7][15] , \SUMB[7][14] , \SUMB[7][13] ,
         \SUMB[7][12] , \SUMB[7][11] , \SUMB[7][10] , \SUMB[7][9] ,
         \SUMB[7][8] , \SUMB[7][7] , \SUMB[7][6] , \SUMB[7][5] , \SUMB[7][4] ,
         \SUMB[7][3] , \SUMB[7][2] , \SUMB[7][1] , \SUMB[6][25] ,
         \SUMB[6][24] , \SUMB[6][23] , \SUMB[6][22] , \SUMB[6][21] ,
         \SUMB[6][20] , \SUMB[6][19] , \SUMB[6][18] , \SUMB[6][17] ,
         \SUMB[6][16] , \SUMB[6][15] , \SUMB[6][14] , \SUMB[6][13] ,
         \SUMB[6][12] , \SUMB[6][11] , \SUMB[6][10] , \SUMB[6][9] ,
         \SUMB[6][8] , \SUMB[6][7] , \SUMB[6][6] , \SUMB[6][5] , \SUMB[6][4] ,
         \SUMB[6][3] , \SUMB[6][2] , \SUMB[6][1] , \SUMB[5][26] ,
         \SUMB[5][25] , \SUMB[5][24] , \SUMB[5][23] , \SUMB[5][22] ,
         \SUMB[5][21] , \SUMB[5][20] , \SUMB[5][19] , \SUMB[5][18] ,
         \SUMB[5][17] , \SUMB[5][16] , \SUMB[5][15] , \SUMB[5][14] ,
         \SUMB[5][13] , \SUMB[5][12] , \SUMB[5][11] , \SUMB[5][10] ,
         \SUMB[5][9] , \SUMB[5][8] , \SUMB[5][7] , \SUMB[5][6] , \SUMB[5][5] ,
         \SUMB[5][4] , \SUMB[5][3] , \SUMB[5][2] , \SUMB[5][1] , \SUMB[4][27] ,
         \SUMB[4][26] , \SUMB[4][25] , \SUMB[4][24] , \SUMB[4][23] ,
         \SUMB[4][22] , \SUMB[4][21] , \SUMB[4][20] , \SUMB[4][19] ,
         \SUMB[4][18] , \SUMB[4][17] , \SUMB[4][16] , \SUMB[4][15] ,
         \SUMB[4][14] , \SUMB[4][13] , \SUMB[4][12] , \SUMB[4][11] ,
         \SUMB[4][10] , \SUMB[4][9] , \SUMB[4][8] , \SUMB[4][7] , \SUMB[4][6] ,
         \SUMB[4][5] , \SUMB[4][4] , \SUMB[4][3] , \SUMB[4][2] , \SUMB[4][1] ,
         \SUMB[3][28] , \SUMB[3][27] , \SUMB[3][26] , \SUMB[3][25] ,
         \SUMB[3][24] , \SUMB[3][23] , \SUMB[3][22] , \SUMB[3][21] ,
         \SUMB[3][20] , \SUMB[3][19] , \SUMB[3][18] , \SUMB[3][17] ,
         \SUMB[3][16] , \SUMB[3][15] , \SUMB[3][14] , \SUMB[3][13] ,
         \SUMB[3][12] , \SUMB[3][11] , \SUMB[3][10] , \SUMB[3][9] ,
         \SUMB[3][8] , \SUMB[3][7] , \SUMB[3][6] , \SUMB[3][5] , \SUMB[3][4] ,
         \SUMB[3][3] , \SUMB[3][2] , \SUMB[3][1] , \SUMB[2][29] ,
         \SUMB[2][28] , \SUMB[2][27] , \SUMB[2][26] , \SUMB[2][25] ,
         \SUMB[2][24] , \SUMB[2][23] , \SUMB[2][22] , \SUMB[2][21] ,
         \SUMB[2][20] , \SUMB[2][19] , \SUMB[2][18] , \SUMB[2][17] ,
         \SUMB[2][16] , \SUMB[2][15] , \SUMB[2][14] , \SUMB[2][13] ,
         \SUMB[2][12] , \SUMB[2][11] , \SUMB[2][10] , \SUMB[2][9] ,
         \SUMB[2][8] , \SUMB[2][7] , \SUMB[2][6] , \SUMB[2][5] , \SUMB[2][4] ,
         \SUMB[2][3] , \SUMB[2][2] , \SUMB[2][1] , \CARRYB[30][0] ,
         \CARRYB[29][1] , \CARRYB[29][0] , \CARRYB[28][2] , \CARRYB[28][1] ,
         \CARRYB[28][0] , \CARRYB[27][3] , \CARRYB[27][2] , \CARRYB[27][1] ,
         \CARRYB[27][0] , \CARRYB[26][4] , \CARRYB[26][3] , \CARRYB[26][2] ,
         \CARRYB[26][1] , \CARRYB[26][0] , \CARRYB[25][5] , \CARRYB[25][4] ,
         \CARRYB[25][3] , \CARRYB[25][2] , \CARRYB[25][1] , \CARRYB[25][0] ,
         \CARRYB[24][6] , \CARRYB[24][5] , \CARRYB[24][4] , \CARRYB[24][3] ,
         \CARRYB[24][2] , \CARRYB[24][1] , \CARRYB[24][0] , \CARRYB[23][7] ,
         \CARRYB[23][6] , \CARRYB[23][5] , \CARRYB[23][4] , \CARRYB[23][3] ,
         \CARRYB[23][2] , \CARRYB[23][1] , \CARRYB[23][0] , \CARRYB[22][8] ,
         \CARRYB[22][7] , \CARRYB[22][6] , \CARRYB[22][5] , \CARRYB[22][4] ,
         \CARRYB[22][3] , \CARRYB[22][2] , \CARRYB[22][1] , \CARRYB[22][0] ,
         \CARRYB[21][9] , \CARRYB[21][8] , \CARRYB[21][7] , \CARRYB[21][6] ,
         \CARRYB[21][5] , \CARRYB[21][4] , \CARRYB[21][3] , \CARRYB[21][2] ,
         \CARRYB[21][1] , \CARRYB[21][0] , \CARRYB[20][10] , \CARRYB[20][9] ,
         \CARRYB[20][8] , \CARRYB[20][7] , \CARRYB[20][6] , \CARRYB[20][5] ,
         \CARRYB[20][4] , \CARRYB[20][3] , \CARRYB[20][2] , \CARRYB[20][1] ,
         \CARRYB[20][0] , \CARRYB[19][11] , \CARRYB[19][10] , \CARRYB[19][9] ,
         \CARRYB[19][8] , \CARRYB[19][7] , \CARRYB[19][6] , \CARRYB[19][5] ,
         \CARRYB[19][4] , \CARRYB[19][3] , \CARRYB[19][2] , \CARRYB[19][1] ,
         \CARRYB[19][0] , \CARRYB[18][12] , \CARRYB[18][11] , \CARRYB[18][10] ,
         \CARRYB[18][9] , \CARRYB[18][8] , \CARRYB[18][7] , \CARRYB[18][6] ,
         \CARRYB[18][5] , \CARRYB[18][4] , \CARRYB[18][3] , \CARRYB[18][2] ,
         \CARRYB[18][1] , \CARRYB[18][0] , \CARRYB[17][13] , \CARRYB[17][12] ,
         \CARRYB[17][11] , \CARRYB[17][10] , \CARRYB[17][9] , \CARRYB[17][8] ,
         \CARRYB[17][7] , \CARRYB[17][6] , \CARRYB[17][5] , \CARRYB[17][4] ,
         \CARRYB[17][3] , \CARRYB[17][2] , \CARRYB[17][1] , \CARRYB[17][0] ,
         \CARRYB[16][14] , \CARRYB[16][13] , \CARRYB[16][12] ,
         \CARRYB[16][11] , \CARRYB[16][10] , \CARRYB[16][9] , \CARRYB[16][8] ,
         \CARRYB[16][7] , \CARRYB[16][6] , \CARRYB[16][5] , \CARRYB[16][4] ,
         \CARRYB[16][3] , \CARRYB[16][2] , \CARRYB[16][1] , \CARRYB[16][0] ,
         \SUMB[30][1] , \SUMB[29][2] , \SUMB[29][1] , \SUMB[28][3] ,
         \SUMB[28][2] , \SUMB[28][1] , \SUMB[27][4] , \SUMB[27][3] ,
         \SUMB[27][2] , \SUMB[27][1] , \SUMB[26][5] , \SUMB[26][4] ,
         \SUMB[26][3] , \SUMB[26][2] , \SUMB[26][1] , \SUMB[25][6] ,
         \SUMB[25][5] , \SUMB[25][4] , \SUMB[25][3] , \SUMB[25][2] ,
         \SUMB[25][1] , \SUMB[24][7] , \SUMB[24][6] , \SUMB[24][5] ,
         \SUMB[24][4] , \SUMB[24][3] , \SUMB[24][2] , \SUMB[24][1] ,
         \SUMB[23][8] , \SUMB[23][7] , \SUMB[23][6] , \SUMB[23][5] ,
         \SUMB[23][4] , \SUMB[23][3] , \SUMB[23][2] , \SUMB[23][1] ,
         \SUMB[22][9] , \SUMB[22][8] , \SUMB[22][7] , \SUMB[22][6] ,
         \SUMB[22][5] , \SUMB[22][4] , \SUMB[22][3] , \SUMB[22][2] ,
         \SUMB[22][1] , \SUMB[21][10] , \SUMB[21][9] , \SUMB[21][8] ,
         \SUMB[21][7] , \SUMB[21][6] , \SUMB[21][5] , \SUMB[21][4] ,
         \SUMB[21][3] , \SUMB[21][2] , \SUMB[21][1] , \SUMB[20][11] ,
         \SUMB[20][10] , \SUMB[20][9] , \SUMB[20][8] , \SUMB[20][7] ,
         \SUMB[20][6] , \SUMB[20][5] , \SUMB[20][4] , \SUMB[20][3] ,
         \SUMB[20][2] , \SUMB[20][1] , \SUMB[19][12] , \SUMB[19][11] ,
         \SUMB[19][10] , \SUMB[19][9] , \SUMB[19][8] , \SUMB[19][7] ,
         \SUMB[19][6] , \SUMB[19][5] , \SUMB[19][4] , \SUMB[19][3] ,
         \SUMB[19][2] , \SUMB[19][1] , \SUMB[18][13] , \SUMB[18][12] ,
         \SUMB[18][11] , \SUMB[18][10] , \SUMB[18][9] , \SUMB[18][8] ,
         \SUMB[18][7] , \SUMB[18][6] , \SUMB[18][5] , \SUMB[18][4] ,
         \SUMB[18][3] , \SUMB[18][2] , \SUMB[18][1] , \SUMB[17][14] ,
         \SUMB[17][13] , \SUMB[17][12] , \SUMB[17][11] , \SUMB[17][10] ,
         \SUMB[17][9] , \SUMB[17][8] , \SUMB[17][7] , \SUMB[17][6] ,
         \SUMB[17][5] , \SUMB[17][4] , \SUMB[17][3] , \SUMB[17][2] ,
         \SUMB[17][1] , \SUMB[16][15] , \SUMB[16][14] , \SUMB[16][13] ,
         \SUMB[16][12] , \SUMB[16][11] , \SUMB[16][10] , \SUMB[16][9] ,
         \SUMB[16][8] , \SUMB[16][7] , \SUMB[16][6] , \SUMB[16][5] ,
         \SUMB[16][4] , \SUMB[16][3] , \SUMB[16][2] , \SUMB[16][1] , n3, n4,
         n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19,
         n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47,
         n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n62,
         n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76,
         n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90,
         n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103,
         n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114,
         n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125,
         n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136,
         n137, n138;

  FA_X1 S4_0 ( .A(\ab[31][0] ), .B(\CARRYB[30][0] ), .CI(\SUMB[30][1] ), .S(
        PRODUCT[31]) );
  FA_X1 S1_30_0 ( .A(\ab[30][0] ), .B(\CARRYB[29][0] ), .CI(\SUMB[29][1] ), 
        .CO(\CARRYB[30][0] ), .S(PRODUCT[30]) );
  FA_X1 S2_30_1 ( .A(\ab[30][1] ), .B(\CARRYB[29][1] ), .CI(\SUMB[29][2] ), 
        .S(\SUMB[30][1] ) );
  FA_X1 S1_29_0 ( .A(\ab[29][0] ), .B(\CARRYB[28][0] ), .CI(\SUMB[28][1] ), 
        .CO(\CARRYB[29][0] ), .S(PRODUCT[29]) );
  FA_X1 S2_29_1 ( .A(\ab[29][1] ), .B(\CARRYB[28][1] ), .CI(\SUMB[28][2] ), 
        .CO(\CARRYB[29][1] ), .S(\SUMB[29][1] ) );
  FA_X1 S2_29_2 ( .A(\ab[29][2] ), .B(\CARRYB[28][2] ), .CI(\SUMB[28][3] ), 
        .S(\SUMB[29][2] ) );
  FA_X1 S1_28_0 ( .A(\ab[28][0] ), .B(\CARRYB[27][0] ), .CI(\SUMB[27][1] ), 
        .CO(\CARRYB[28][0] ), .S(PRODUCT[28]) );
  FA_X1 S2_28_1 ( .A(\ab[28][1] ), .B(\CARRYB[27][1] ), .CI(\SUMB[27][2] ), 
        .CO(\CARRYB[28][1] ), .S(\SUMB[28][1] ) );
  FA_X1 S2_28_2 ( .A(\ab[28][2] ), .B(\CARRYB[27][2] ), .CI(\SUMB[27][3] ), 
        .CO(\CARRYB[28][2] ), .S(\SUMB[28][2] ) );
  FA_X1 S2_28_3 ( .A(\ab[28][3] ), .B(\CARRYB[27][3] ), .CI(\SUMB[27][4] ), 
        .S(\SUMB[28][3] ) );
  FA_X1 S1_27_0 ( .A(\ab[27][0] ), .B(\CARRYB[26][0] ), .CI(\SUMB[26][1] ), 
        .CO(\CARRYB[27][0] ), .S(PRODUCT[27]) );
  FA_X1 S2_27_1 ( .A(\ab[27][1] ), .B(\CARRYB[26][1] ), .CI(\SUMB[26][2] ), 
        .CO(\CARRYB[27][1] ), .S(\SUMB[27][1] ) );
  FA_X1 S2_27_2 ( .A(\ab[27][2] ), .B(\CARRYB[26][2] ), .CI(\SUMB[26][3] ), 
        .CO(\CARRYB[27][2] ), .S(\SUMB[27][2] ) );
  FA_X1 S2_27_3 ( .A(\ab[27][3] ), .B(\CARRYB[26][3] ), .CI(\SUMB[26][4] ), 
        .CO(\CARRYB[27][3] ), .S(\SUMB[27][3] ) );
  FA_X1 S2_27_4 ( .A(\ab[27][4] ), .B(\CARRYB[26][4] ), .CI(\SUMB[26][5] ), 
        .S(\SUMB[27][4] ) );
  FA_X1 S1_26_0 ( .A(\ab[26][0] ), .B(\CARRYB[25][0] ), .CI(\SUMB[25][1] ), 
        .CO(\CARRYB[26][0] ), .S(PRODUCT[26]) );
  FA_X1 S2_26_1 ( .A(\ab[26][1] ), .B(\CARRYB[25][1] ), .CI(\SUMB[25][2] ), 
        .CO(\CARRYB[26][1] ), .S(\SUMB[26][1] ) );
  FA_X1 S2_26_2 ( .A(\ab[26][2] ), .B(\CARRYB[25][2] ), .CI(\SUMB[25][3] ), 
        .CO(\CARRYB[26][2] ), .S(\SUMB[26][2] ) );
  FA_X1 S2_26_3 ( .A(\ab[26][3] ), .B(\CARRYB[25][3] ), .CI(\SUMB[25][4] ), 
        .CO(\CARRYB[26][3] ), .S(\SUMB[26][3] ) );
  FA_X1 S2_26_4 ( .A(\ab[26][4] ), .B(\CARRYB[25][4] ), .CI(\SUMB[25][5] ), 
        .CO(\CARRYB[26][4] ), .S(\SUMB[26][4] ) );
  FA_X1 S2_26_5 ( .A(\ab[26][5] ), .B(\CARRYB[25][5] ), .CI(\SUMB[25][6] ), 
        .S(\SUMB[26][5] ) );
  FA_X1 S1_25_0 ( .A(\ab[25][0] ), .B(\CARRYB[24][0] ), .CI(\SUMB[24][1] ), 
        .CO(\CARRYB[25][0] ), .S(PRODUCT[25]) );
  FA_X1 S2_25_1 ( .A(\ab[25][1] ), .B(\CARRYB[24][1] ), .CI(\SUMB[24][2] ), 
        .CO(\CARRYB[25][1] ), .S(\SUMB[25][1] ) );
  FA_X1 S2_25_2 ( .A(\ab[25][2] ), .B(\CARRYB[24][2] ), .CI(\SUMB[24][3] ), 
        .CO(\CARRYB[25][2] ), .S(\SUMB[25][2] ) );
  FA_X1 S2_25_3 ( .A(\ab[25][3] ), .B(\CARRYB[24][3] ), .CI(\SUMB[24][4] ), 
        .CO(\CARRYB[25][3] ), .S(\SUMB[25][3] ) );
  FA_X1 S2_25_4 ( .A(\ab[25][4] ), .B(\CARRYB[24][4] ), .CI(\SUMB[24][5] ), 
        .CO(\CARRYB[25][4] ), .S(\SUMB[25][4] ) );
  FA_X1 S2_25_5 ( .A(\ab[25][5] ), .B(\CARRYB[24][5] ), .CI(\SUMB[24][6] ), 
        .CO(\CARRYB[25][5] ), .S(\SUMB[25][5] ) );
  FA_X1 S2_25_6 ( .A(\ab[25][6] ), .B(\CARRYB[24][6] ), .CI(\SUMB[24][7] ), 
        .S(\SUMB[25][6] ) );
  FA_X1 S1_24_0 ( .A(\ab[24][0] ), .B(\CARRYB[23][0] ), .CI(\SUMB[23][1] ), 
        .CO(\CARRYB[24][0] ), .S(PRODUCT[24]) );
  FA_X1 S2_24_1 ( .A(\ab[24][1] ), .B(\CARRYB[23][1] ), .CI(\SUMB[23][2] ), 
        .CO(\CARRYB[24][1] ), .S(\SUMB[24][1] ) );
  FA_X1 S2_24_2 ( .A(\ab[24][2] ), .B(\CARRYB[23][2] ), .CI(\SUMB[23][3] ), 
        .CO(\CARRYB[24][2] ), .S(\SUMB[24][2] ) );
  FA_X1 S2_24_3 ( .A(\ab[24][3] ), .B(\CARRYB[23][3] ), .CI(\SUMB[23][4] ), 
        .CO(\CARRYB[24][3] ), .S(\SUMB[24][3] ) );
  FA_X1 S2_24_4 ( .A(\ab[24][4] ), .B(\CARRYB[23][4] ), .CI(\SUMB[23][5] ), 
        .CO(\CARRYB[24][4] ), .S(\SUMB[24][4] ) );
  FA_X1 S2_24_5 ( .A(\ab[24][5] ), .B(\CARRYB[23][5] ), .CI(\SUMB[23][6] ), 
        .CO(\CARRYB[24][5] ), .S(\SUMB[24][5] ) );
  FA_X1 S2_24_6 ( .A(\ab[24][6] ), .B(\CARRYB[23][6] ), .CI(\SUMB[23][7] ), 
        .CO(\CARRYB[24][6] ), .S(\SUMB[24][6] ) );
  FA_X1 S2_24_7 ( .A(\ab[24][7] ), .B(\CARRYB[23][7] ), .CI(\SUMB[23][8] ), 
        .S(\SUMB[24][7] ) );
  FA_X1 S1_23_0 ( .A(\ab[23][0] ), .B(\CARRYB[22][0] ), .CI(\SUMB[22][1] ), 
        .CO(\CARRYB[23][0] ), .S(PRODUCT[23]) );
  FA_X1 S2_23_1 ( .A(\ab[23][1] ), .B(\CARRYB[22][1] ), .CI(\SUMB[22][2] ), 
        .CO(\CARRYB[23][1] ), .S(\SUMB[23][1] ) );
  FA_X1 S2_23_2 ( .A(\ab[23][2] ), .B(\CARRYB[22][2] ), .CI(\SUMB[22][3] ), 
        .CO(\CARRYB[23][2] ), .S(\SUMB[23][2] ) );
  FA_X1 S2_23_3 ( .A(\ab[23][3] ), .B(\CARRYB[22][3] ), .CI(\SUMB[22][4] ), 
        .CO(\CARRYB[23][3] ), .S(\SUMB[23][3] ) );
  FA_X1 S2_23_4 ( .A(\ab[23][4] ), .B(\CARRYB[22][4] ), .CI(\SUMB[22][5] ), 
        .CO(\CARRYB[23][4] ), .S(\SUMB[23][4] ) );
  FA_X1 S2_23_5 ( .A(\ab[23][5] ), .B(\CARRYB[22][5] ), .CI(\SUMB[22][6] ), 
        .CO(\CARRYB[23][5] ), .S(\SUMB[23][5] ) );
  FA_X1 S2_23_6 ( .A(\ab[23][6] ), .B(\CARRYB[22][6] ), .CI(\SUMB[22][7] ), 
        .CO(\CARRYB[23][6] ), .S(\SUMB[23][6] ) );
  FA_X1 S2_23_7 ( .A(\ab[23][7] ), .B(\CARRYB[22][7] ), .CI(\SUMB[22][8] ), 
        .CO(\CARRYB[23][7] ), .S(\SUMB[23][7] ) );
  FA_X1 S2_23_8 ( .A(\ab[23][8] ), .B(\CARRYB[22][8] ), .CI(\SUMB[22][9] ), 
        .S(\SUMB[23][8] ) );
  FA_X1 S1_22_0 ( .A(\ab[22][0] ), .B(\CARRYB[21][0] ), .CI(\SUMB[21][1] ), 
        .CO(\CARRYB[22][0] ), .S(PRODUCT[22]) );
  FA_X1 S2_22_1 ( .A(\ab[22][1] ), .B(\CARRYB[21][1] ), .CI(\SUMB[21][2] ), 
        .CO(\CARRYB[22][1] ), .S(\SUMB[22][1] ) );
  FA_X1 S2_22_2 ( .A(\ab[22][2] ), .B(\CARRYB[21][2] ), .CI(\SUMB[21][3] ), 
        .CO(\CARRYB[22][2] ), .S(\SUMB[22][2] ) );
  FA_X1 S2_22_3 ( .A(\ab[22][3] ), .B(\CARRYB[21][3] ), .CI(\SUMB[21][4] ), 
        .CO(\CARRYB[22][3] ), .S(\SUMB[22][3] ) );
  FA_X1 S2_22_4 ( .A(\ab[22][4] ), .B(\CARRYB[21][4] ), .CI(\SUMB[21][5] ), 
        .CO(\CARRYB[22][4] ), .S(\SUMB[22][4] ) );
  FA_X1 S2_22_5 ( .A(\ab[22][5] ), .B(\CARRYB[21][5] ), .CI(\SUMB[21][6] ), 
        .CO(\CARRYB[22][5] ), .S(\SUMB[22][5] ) );
  FA_X1 S2_22_6 ( .A(\ab[22][6] ), .B(\CARRYB[21][6] ), .CI(\SUMB[21][7] ), 
        .CO(\CARRYB[22][6] ), .S(\SUMB[22][6] ) );
  FA_X1 S2_22_7 ( .A(\ab[22][7] ), .B(\CARRYB[21][7] ), .CI(\SUMB[21][8] ), 
        .CO(\CARRYB[22][7] ), .S(\SUMB[22][7] ) );
  FA_X1 S2_22_8 ( .A(\ab[22][8] ), .B(\CARRYB[21][8] ), .CI(\SUMB[21][9] ), 
        .CO(\CARRYB[22][8] ), .S(\SUMB[22][8] ) );
  FA_X1 S2_22_9 ( .A(\ab[22][9] ), .B(\CARRYB[21][9] ), .CI(\SUMB[21][10] ), 
        .S(\SUMB[22][9] ) );
  FA_X1 S1_21_0 ( .A(\ab[21][0] ), .B(\CARRYB[20][0] ), .CI(\SUMB[20][1] ), 
        .CO(\CARRYB[21][0] ), .S(PRODUCT[21]) );
  FA_X1 S2_21_1 ( .A(\ab[21][1] ), .B(\CARRYB[20][1] ), .CI(\SUMB[20][2] ), 
        .CO(\CARRYB[21][1] ), .S(\SUMB[21][1] ) );
  FA_X1 S2_21_2 ( .A(\ab[21][2] ), .B(\CARRYB[20][2] ), .CI(\SUMB[20][3] ), 
        .CO(\CARRYB[21][2] ), .S(\SUMB[21][2] ) );
  FA_X1 S2_21_3 ( .A(\ab[21][3] ), .B(\CARRYB[20][3] ), .CI(\SUMB[20][4] ), 
        .CO(\CARRYB[21][3] ), .S(\SUMB[21][3] ) );
  FA_X1 S2_21_4 ( .A(\ab[21][4] ), .B(\CARRYB[20][4] ), .CI(\SUMB[20][5] ), 
        .CO(\CARRYB[21][4] ), .S(\SUMB[21][4] ) );
  FA_X1 S2_21_5 ( .A(\ab[21][5] ), .B(\CARRYB[20][5] ), .CI(\SUMB[20][6] ), 
        .CO(\CARRYB[21][5] ), .S(\SUMB[21][5] ) );
  FA_X1 S2_21_6 ( .A(\ab[21][6] ), .B(\CARRYB[20][6] ), .CI(\SUMB[20][7] ), 
        .CO(\CARRYB[21][6] ), .S(\SUMB[21][6] ) );
  FA_X1 S2_21_7 ( .A(\ab[21][7] ), .B(\CARRYB[20][7] ), .CI(\SUMB[20][8] ), 
        .CO(\CARRYB[21][7] ), .S(\SUMB[21][7] ) );
  FA_X1 S2_21_8 ( .A(\ab[21][8] ), .B(\CARRYB[20][8] ), .CI(\SUMB[20][9] ), 
        .CO(\CARRYB[21][8] ), .S(\SUMB[21][8] ) );
  FA_X1 S2_21_9 ( .A(\ab[21][9] ), .B(\CARRYB[20][9] ), .CI(\SUMB[20][10] ), 
        .CO(\CARRYB[21][9] ), .S(\SUMB[21][9] ) );
  FA_X1 S2_21_10 ( .A(\ab[21][10] ), .B(\CARRYB[20][10] ), .CI(\SUMB[20][11] ), 
        .S(\SUMB[21][10] ) );
  FA_X1 S1_20_0 ( .A(\ab[20][0] ), .B(\CARRYB[19][0] ), .CI(\SUMB[19][1] ), 
        .CO(\CARRYB[20][0] ), .S(PRODUCT[20]) );
  FA_X1 S2_20_1 ( .A(\ab[20][1] ), .B(\CARRYB[19][1] ), .CI(\SUMB[19][2] ), 
        .CO(\CARRYB[20][1] ), .S(\SUMB[20][1] ) );
  FA_X1 S2_20_2 ( .A(\ab[20][2] ), .B(\CARRYB[19][2] ), .CI(\SUMB[19][3] ), 
        .CO(\CARRYB[20][2] ), .S(\SUMB[20][2] ) );
  FA_X1 S2_20_3 ( .A(\ab[20][3] ), .B(\CARRYB[19][3] ), .CI(\SUMB[19][4] ), 
        .CO(\CARRYB[20][3] ), .S(\SUMB[20][3] ) );
  FA_X1 S2_20_4 ( .A(\ab[20][4] ), .B(\CARRYB[19][4] ), .CI(\SUMB[19][5] ), 
        .CO(\CARRYB[20][4] ), .S(\SUMB[20][4] ) );
  FA_X1 S2_20_5 ( .A(\ab[20][5] ), .B(\CARRYB[19][5] ), .CI(\SUMB[19][6] ), 
        .CO(\CARRYB[20][5] ), .S(\SUMB[20][5] ) );
  FA_X1 S2_20_6 ( .A(\ab[20][6] ), .B(\CARRYB[19][6] ), .CI(\SUMB[19][7] ), 
        .CO(\CARRYB[20][6] ), .S(\SUMB[20][6] ) );
  FA_X1 S2_20_7 ( .A(\ab[20][7] ), .B(\CARRYB[19][7] ), .CI(\SUMB[19][8] ), 
        .CO(\CARRYB[20][7] ), .S(\SUMB[20][7] ) );
  FA_X1 S2_20_8 ( .A(\ab[20][8] ), .B(\CARRYB[19][8] ), .CI(\SUMB[19][9] ), 
        .CO(\CARRYB[20][8] ), .S(\SUMB[20][8] ) );
  FA_X1 S2_20_9 ( .A(\ab[20][9] ), .B(\CARRYB[19][9] ), .CI(\SUMB[19][10] ), 
        .CO(\CARRYB[20][9] ), .S(\SUMB[20][9] ) );
  FA_X1 S2_20_10 ( .A(\ab[20][10] ), .B(\CARRYB[19][10] ), .CI(\SUMB[19][11] ), 
        .CO(\CARRYB[20][10] ), .S(\SUMB[20][10] ) );
  FA_X1 S2_20_11 ( .A(\ab[20][11] ), .B(\CARRYB[19][11] ), .CI(\SUMB[19][12] ), 
        .S(\SUMB[20][11] ) );
  FA_X1 S1_19_0 ( .A(\ab[19][0] ), .B(\CARRYB[18][0] ), .CI(\SUMB[18][1] ), 
        .CO(\CARRYB[19][0] ), .S(PRODUCT[19]) );
  FA_X1 S2_19_1 ( .A(\ab[19][1] ), .B(\CARRYB[18][1] ), .CI(\SUMB[18][2] ), 
        .CO(\CARRYB[19][1] ), .S(\SUMB[19][1] ) );
  FA_X1 S2_19_2 ( .A(\ab[19][2] ), .B(\CARRYB[18][2] ), .CI(\SUMB[18][3] ), 
        .CO(\CARRYB[19][2] ), .S(\SUMB[19][2] ) );
  FA_X1 S2_19_3 ( .A(\ab[19][3] ), .B(\CARRYB[18][3] ), .CI(\SUMB[18][4] ), 
        .CO(\CARRYB[19][3] ), .S(\SUMB[19][3] ) );
  FA_X1 S2_19_4 ( .A(\ab[19][4] ), .B(\CARRYB[18][4] ), .CI(\SUMB[18][5] ), 
        .CO(\CARRYB[19][4] ), .S(\SUMB[19][4] ) );
  FA_X1 S2_19_5 ( .A(\ab[19][5] ), .B(\CARRYB[18][5] ), .CI(\SUMB[18][6] ), 
        .CO(\CARRYB[19][5] ), .S(\SUMB[19][5] ) );
  FA_X1 S2_19_6 ( .A(\ab[19][6] ), .B(\CARRYB[18][6] ), .CI(\SUMB[18][7] ), 
        .CO(\CARRYB[19][6] ), .S(\SUMB[19][6] ) );
  FA_X1 S2_19_7 ( .A(\ab[19][7] ), .B(\CARRYB[18][7] ), .CI(\SUMB[18][8] ), 
        .CO(\CARRYB[19][7] ), .S(\SUMB[19][7] ) );
  FA_X1 S2_19_8 ( .A(\ab[19][8] ), .B(\CARRYB[18][8] ), .CI(\SUMB[18][9] ), 
        .CO(\CARRYB[19][8] ), .S(\SUMB[19][8] ) );
  FA_X1 S2_19_9 ( .A(\ab[19][9] ), .B(\CARRYB[18][9] ), .CI(\SUMB[18][10] ), 
        .CO(\CARRYB[19][9] ), .S(\SUMB[19][9] ) );
  FA_X1 S2_19_10 ( .A(\ab[19][10] ), .B(\CARRYB[18][10] ), .CI(\SUMB[18][11] ), 
        .CO(\CARRYB[19][10] ), .S(\SUMB[19][10] ) );
  FA_X1 S2_19_11 ( .A(\ab[19][11] ), .B(\CARRYB[18][11] ), .CI(\SUMB[18][12] ), 
        .CO(\CARRYB[19][11] ), .S(\SUMB[19][11] ) );
  FA_X1 S2_19_12 ( .A(\ab[19][12] ), .B(\CARRYB[18][12] ), .CI(\SUMB[18][13] ), 
        .S(\SUMB[19][12] ) );
  FA_X1 S1_18_0 ( .A(\ab[18][0] ), .B(\CARRYB[17][0] ), .CI(\SUMB[17][1] ), 
        .CO(\CARRYB[18][0] ), .S(PRODUCT[18]) );
  FA_X1 S2_18_1 ( .A(\ab[18][1] ), .B(\CARRYB[17][1] ), .CI(\SUMB[17][2] ), 
        .CO(\CARRYB[18][1] ), .S(\SUMB[18][1] ) );
  FA_X1 S2_18_2 ( .A(\ab[18][2] ), .B(\CARRYB[17][2] ), .CI(\SUMB[17][3] ), 
        .CO(\CARRYB[18][2] ), .S(\SUMB[18][2] ) );
  FA_X1 S2_18_3 ( .A(\ab[18][3] ), .B(\CARRYB[17][3] ), .CI(\SUMB[17][4] ), 
        .CO(\CARRYB[18][3] ), .S(\SUMB[18][3] ) );
  FA_X1 S2_18_4 ( .A(\ab[18][4] ), .B(\CARRYB[17][4] ), .CI(\SUMB[17][5] ), 
        .CO(\CARRYB[18][4] ), .S(\SUMB[18][4] ) );
  FA_X1 S2_18_5 ( .A(\ab[18][5] ), .B(\CARRYB[17][5] ), .CI(\SUMB[17][6] ), 
        .CO(\CARRYB[18][5] ), .S(\SUMB[18][5] ) );
  FA_X1 S2_18_6 ( .A(\ab[18][6] ), .B(\CARRYB[17][6] ), .CI(\SUMB[17][7] ), 
        .CO(\CARRYB[18][6] ), .S(\SUMB[18][6] ) );
  FA_X1 S2_18_7 ( .A(\ab[18][7] ), .B(\CARRYB[17][7] ), .CI(\SUMB[17][8] ), 
        .CO(\CARRYB[18][7] ), .S(\SUMB[18][7] ) );
  FA_X1 S2_18_8 ( .A(\ab[18][8] ), .B(\CARRYB[17][8] ), .CI(\SUMB[17][9] ), 
        .CO(\CARRYB[18][8] ), .S(\SUMB[18][8] ) );
  FA_X1 S2_18_9 ( .A(\ab[18][9] ), .B(\CARRYB[17][9] ), .CI(\SUMB[17][10] ), 
        .CO(\CARRYB[18][9] ), .S(\SUMB[18][9] ) );
  FA_X1 S2_18_10 ( .A(\ab[18][10] ), .B(\CARRYB[17][10] ), .CI(\SUMB[17][11] ), 
        .CO(\CARRYB[18][10] ), .S(\SUMB[18][10] ) );
  FA_X1 S2_18_11 ( .A(\ab[18][11] ), .B(\CARRYB[17][11] ), .CI(\SUMB[17][12] ), 
        .CO(\CARRYB[18][11] ), .S(\SUMB[18][11] ) );
  FA_X1 S2_18_12 ( .A(\ab[18][12] ), .B(\CARRYB[17][12] ), .CI(\SUMB[17][13] ), 
        .CO(\CARRYB[18][12] ), .S(\SUMB[18][12] ) );
  FA_X1 S2_18_13 ( .A(\ab[18][13] ), .B(\CARRYB[17][13] ), .CI(\SUMB[17][14] ), 
        .S(\SUMB[18][13] ) );
  FA_X1 S1_17_0 ( .A(\ab[17][0] ), .B(\CARRYB[16][0] ), .CI(\SUMB[16][1] ), 
        .CO(\CARRYB[17][0] ), .S(PRODUCT[17]) );
  FA_X1 S2_17_1 ( .A(\ab[17][1] ), .B(\CARRYB[16][1] ), .CI(\SUMB[16][2] ), 
        .CO(\CARRYB[17][1] ), .S(\SUMB[17][1] ) );
  FA_X1 S2_17_2 ( .A(\ab[17][2] ), .B(\CARRYB[16][2] ), .CI(\SUMB[16][3] ), 
        .CO(\CARRYB[17][2] ), .S(\SUMB[17][2] ) );
  FA_X1 S2_17_3 ( .A(\ab[17][3] ), .B(\CARRYB[16][3] ), .CI(\SUMB[16][4] ), 
        .CO(\CARRYB[17][3] ), .S(\SUMB[17][3] ) );
  FA_X1 S2_17_4 ( .A(\ab[17][4] ), .B(\CARRYB[16][4] ), .CI(\SUMB[16][5] ), 
        .CO(\CARRYB[17][4] ), .S(\SUMB[17][4] ) );
  FA_X1 S2_17_5 ( .A(\ab[17][5] ), .B(\CARRYB[16][5] ), .CI(\SUMB[16][6] ), 
        .CO(\CARRYB[17][5] ), .S(\SUMB[17][5] ) );
  FA_X1 S2_17_6 ( .A(\ab[17][6] ), .B(\CARRYB[16][6] ), .CI(\SUMB[16][7] ), 
        .CO(\CARRYB[17][6] ), .S(\SUMB[17][6] ) );
  FA_X1 S2_17_7 ( .A(\ab[17][7] ), .B(\CARRYB[16][7] ), .CI(\SUMB[16][8] ), 
        .CO(\CARRYB[17][7] ), .S(\SUMB[17][7] ) );
  FA_X1 S2_17_8 ( .A(\ab[17][8] ), .B(\CARRYB[16][8] ), .CI(\SUMB[16][9] ), 
        .CO(\CARRYB[17][8] ), .S(\SUMB[17][8] ) );
  FA_X1 S2_17_9 ( .A(\ab[17][9] ), .B(\CARRYB[16][9] ), .CI(\SUMB[16][10] ), 
        .CO(\CARRYB[17][9] ), .S(\SUMB[17][9] ) );
  FA_X1 S2_17_10 ( .A(\ab[17][10] ), .B(\CARRYB[16][10] ), .CI(\SUMB[16][11] ), 
        .CO(\CARRYB[17][10] ), .S(\SUMB[17][10] ) );
  FA_X1 S2_17_11 ( .A(\ab[17][11] ), .B(\CARRYB[16][11] ), .CI(\SUMB[16][12] ), 
        .CO(\CARRYB[17][11] ), .S(\SUMB[17][11] ) );
  FA_X1 S2_17_12 ( .A(\ab[17][12] ), .B(\CARRYB[16][12] ), .CI(\SUMB[16][13] ), 
        .CO(\CARRYB[17][12] ), .S(\SUMB[17][12] ) );
  FA_X1 S2_17_13 ( .A(\ab[17][13] ), .B(\CARRYB[16][13] ), .CI(\SUMB[16][14] ), 
        .CO(\CARRYB[17][13] ), .S(\SUMB[17][13] ) );
  FA_X1 S2_17_14 ( .A(\ab[17][14] ), .B(\CARRYB[16][14] ), .CI(\SUMB[16][15] ), 
        .S(\SUMB[17][14] ) );
  FA_X1 S1_16_0 ( .A(\ab[16][0] ), .B(\CARRYB[15][0] ), .CI(\SUMB[15][1] ), 
        .CO(\CARRYB[16][0] ), .S(PRODUCT[16]) );
  FA_X1 S2_16_1 ( .A(\ab[16][1] ), .B(\CARRYB[15][1] ), .CI(\SUMB[15][2] ), 
        .CO(\CARRYB[16][1] ), .S(\SUMB[16][1] ) );
  FA_X1 S2_16_2 ( .A(\ab[16][2] ), .B(\CARRYB[15][2] ), .CI(\SUMB[15][3] ), 
        .CO(\CARRYB[16][2] ), .S(\SUMB[16][2] ) );
  FA_X1 S2_16_3 ( .A(\ab[16][3] ), .B(\CARRYB[15][3] ), .CI(\SUMB[15][4] ), 
        .CO(\CARRYB[16][3] ), .S(\SUMB[16][3] ) );
  FA_X1 S2_16_4 ( .A(\ab[16][4] ), .B(\CARRYB[15][4] ), .CI(\SUMB[15][5] ), 
        .CO(\CARRYB[16][4] ), .S(\SUMB[16][4] ) );
  FA_X1 S2_16_5 ( .A(\ab[16][5] ), .B(\CARRYB[15][5] ), .CI(\SUMB[15][6] ), 
        .CO(\CARRYB[16][5] ), .S(\SUMB[16][5] ) );
  FA_X1 S2_16_6 ( .A(\ab[16][6] ), .B(\CARRYB[15][6] ), .CI(\SUMB[15][7] ), 
        .CO(\CARRYB[16][6] ), .S(\SUMB[16][6] ) );
  FA_X1 S2_16_7 ( .A(\ab[16][7] ), .B(\CARRYB[15][7] ), .CI(\SUMB[15][8] ), 
        .CO(\CARRYB[16][7] ), .S(\SUMB[16][7] ) );
  FA_X1 S2_16_8 ( .A(\ab[16][8] ), .B(\CARRYB[15][8] ), .CI(\SUMB[15][9] ), 
        .CO(\CARRYB[16][8] ), .S(\SUMB[16][8] ) );
  FA_X1 S2_16_9 ( .A(\ab[16][9] ), .B(\CARRYB[15][9] ), .CI(\SUMB[15][10] ), 
        .CO(\CARRYB[16][9] ), .S(\SUMB[16][9] ) );
  FA_X1 S2_16_10 ( .A(\ab[16][10] ), .B(\CARRYB[15][10] ), .CI(\SUMB[15][11] ), 
        .CO(\CARRYB[16][10] ), .S(\SUMB[16][10] ) );
  FA_X1 S2_16_11 ( .A(\ab[16][11] ), .B(\CARRYB[15][11] ), .CI(\SUMB[15][12] ), 
        .CO(\CARRYB[16][11] ), .S(\SUMB[16][11] ) );
  FA_X1 S2_16_12 ( .A(\ab[16][12] ), .B(\CARRYB[15][12] ), .CI(\SUMB[15][13] ), 
        .CO(\CARRYB[16][12] ), .S(\SUMB[16][12] ) );
  FA_X1 S2_16_13 ( .A(\ab[16][13] ), .B(\CARRYB[15][13] ), .CI(\SUMB[15][14] ), 
        .CO(\CARRYB[16][13] ), .S(\SUMB[16][13] ) );
  FA_X1 S2_16_14 ( .A(\ab[16][14] ), .B(\CARRYB[15][14] ), .CI(\SUMB[15][15] ), 
        .CO(\CARRYB[16][14] ), .S(\SUMB[16][14] ) );
  FA_X1 S2_16_15 ( .A(\ab[16][15] ), .B(\CARRYB[15][15] ), .CI(\SUMB[15][16] ), 
        .S(\SUMB[16][15] ) );
  FA_X1 S1_15_0 ( .A(\ab[15][0] ), .B(\CARRYB[14][0] ), .CI(\SUMB[14][1] ), 
        .CO(\CARRYB[15][0] ), .S(PRODUCT[15]) );
  FA_X1 S2_15_1 ( .A(\ab[15][1] ), .B(\CARRYB[14][1] ), .CI(\SUMB[14][2] ), 
        .CO(\CARRYB[15][1] ), .S(\SUMB[15][1] ) );
  FA_X1 S2_15_2 ( .A(\ab[15][2] ), .B(\CARRYB[14][2] ), .CI(\SUMB[14][3] ), 
        .CO(\CARRYB[15][2] ), .S(\SUMB[15][2] ) );
  FA_X1 S2_15_3 ( .A(\ab[15][3] ), .B(\CARRYB[14][3] ), .CI(\SUMB[14][4] ), 
        .CO(\CARRYB[15][3] ), .S(\SUMB[15][3] ) );
  FA_X1 S2_15_4 ( .A(\ab[15][4] ), .B(\CARRYB[14][4] ), .CI(\SUMB[14][5] ), 
        .CO(\CARRYB[15][4] ), .S(\SUMB[15][4] ) );
  FA_X1 S2_15_5 ( .A(\ab[15][5] ), .B(\CARRYB[14][5] ), .CI(\SUMB[14][6] ), 
        .CO(\CARRYB[15][5] ), .S(\SUMB[15][5] ) );
  FA_X1 S2_15_6 ( .A(\ab[15][6] ), .B(\CARRYB[14][6] ), .CI(\SUMB[14][7] ), 
        .CO(\CARRYB[15][6] ), .S(\SUMB[15][6] ) );
  FA_X1 S2_15_7 ( .A(\ab[15][7] ), .B(\CARRYB[14][7] ), .CI(\SUMB[14][8] ), 
        .CO(\CARRYB[15][7] ), .S(\SUMB[15][7] ) );
  FA_X1 S2_15_8 ( .A(\ab[15][8] ), .B(\CARRYB[14][8] ), .CI(\SUMB[14][9] ), 
        .CO(\CARRYB[15][8] ), .S(\SUMB[15][8] ) );
  FA_X1 S2_15_9 ( .A(\ab[15][9] ), .B(\CARRYB[14][9] ), .CI(\SUMB[14][10] ), 
        .CO(\CARRYB[15][9] ), .S(\SUMB[15][9] ) );
  FA_X1 S2_15_10 ( .A(\ab[15][10] ), .B(\CARRYB[14][10] ), .CI(\SUMB[14][11] ), 
        .CO(\CARRYB[15][10] ), .S(\SUMB[15][10] ) );
  FA_X1 S2_15_11 ( .A(\ab[15][11] ), .B(\CARRYB[14][11] ), .CI(\SUMB[14][12] ), 
        .CO(\CARRYB[15][11] ), .S(\SUMB[15][11] ) );
  FA_X1 S2_15_12 ( .A(\ab[15][12] ), .B(\CARRYB[14][12] ), .CI(\SUMB[14][13] ), 
        .CO(\CARRYB[15][12] ), .S(\SUMB[15][12] ) );
  FA_X1 S2_15_13 ( .A(\ab[15][13] ), .B(\CARRYB[14][13] ), .CI(\SUMB[14][14] ), 
        .CO(\CARRYB[15][13] ), .S(\SUMB[15][13] ) );
  FA_X1 S2_15_14 ( .A(\ab[15][14] ), .B(\CARRYB[14][14] ), .CI(\SUMB[14][15] ), 
        .CO(\CARRYB[15][14] ), .S(\SUMB[15][14] ) );
  FA_X1 S2_15_15 ( .A(\ab[15][15] ), .B(\CARRYB[14][15] ), .CI(\SUMB[14][16] ), 
        .CO(\CARRYB[15][15] ), .S(\SUMB[15][15] ) );
  FA_X1 S2_15_16 ( .A(\ab[15][16] ), .B(\CARRYB[14][16] ), .CI(\SUMB[14][17] ), 
        .S(\SUMB[15][16] ) );
  FA_X1 S1_14_0 ( .A(\ab[14][0] ), .B(\CARRYB[13][0] ), .CI(\SUMB[13][1] ), 
        .CO(\CARRYB[14][0] ), .S(PRODUCT[14]) );
  FA_X1 S2_14_1 ( .A(\ab[14][1] ), .B(\CARRYB[13][1] ), .CI(\SUMB[13][2] ), 
        .CO(\CARRYB[14][1] ), .S(\SUMB[14][1] ) );
  FA_X1 S2_14_2 ( .A(\ab[14][2] ), .B(\CARRYB[13][2] ), .CI(\SUMB[13][3] ), 
        .CO(\CARRYB[14][2] ), .S(\SUMB[14][2] ) );
  FA_X1 S2_14_3 ( .A(\ab[14][3] ), .B(\CARRYB[13][3] ), .CI(\SUMB[13][4] ), 
        .CO(\CARRYB[14][3] ), .S(\SUMB[14][3] ) );
  FA_X1 S2_14_4 ( .A(\ab[14][4] ), .B(\CARRYB[13][4] ), .CI(\SUMB[13][5] ), 
        .CO(\CARRYB[14][4] ), .S(\SUMB[14][4] ) );
  FA_X1 S2_14_5 ( .A(\ab[14][5] ), .B(\CARRYB[13][5] ), .CI(\SUMB[13][6] ), 
        .CO(\CARRYB[14][5] ), .S(\SUMB[14][5] ) );
  FA_X1 S2_14_6 ( .A(\ab[14][6] ), .B(\CARRYB[13][6] ), .CI(\SUMB[13][7] ), 
        .CO(\CARRYB[14][6] ), .S(\SUMB[14][6] ) );
  FA_X1 S2_14_7 ( .A(\ab[14][7] ), .B(\CARRYB[13][7] ), .CI(\SUMB[13][8] ), 
        .CO(\CARRYB[14][7] ), .S(\SUMB[14][7] ) );
  FA_X1 S2_14_8 ( .A(\ab[14][8] ), .B(\CARRYB[13][8] ), .CI(\SUMB[13][9] ), 
        .CO(\CARRYB[14][8] ), .S(\SUMB[14][8] ) );
  FA_X1 S2_14_9 ( .A(\ab[14][9] ), .B(\CARRYB[13][9] ), .CI(\SUMB[13][10] ), 
        .CO(\CARRYB[14][9] ), .S(\SUMB[14][9] ) );
  FA_X1 S2_14_10 ( .A(\ab[14][10] ), .B(\CARRYB[13][10] ), .CI(\SUMB[13][11] ), 
        .CO(\CARRYB[14][10] ), .S(\SUMB[14][10] ) );
  FA_X1 S2_14_11 ( .A(\ab[14][11] ), .B(\CARRYB[13][11] ), .CI(\SUMB[13][12] ), 
        .CO(\CARRYB[14][11] ), .S(\SUMB[14][11] ) );
  FA_X1 S2_14_12 ( .A(\ab[14][12] ), .B(\CARRYB[13][12] ), .CI(\SUMB[13][13] ), 
        .CO(\CARRYB[14][12] ), .S(\SUMB[14][12] ) );
  FA_X1 S2_14_13 ( .A(\ab[14][13] ), .B(\CARRYB[13][13] ), .CI(\SUMB[13][14] ), 
        .CO(\CARRYB[14][13] ), .S(\SUMB[14][13] ) );
  FA_X1 S2_14_14 ( .A(\ab[14][14] ), .B(\CARRYB[13][14] ), .CI(\SUMB[13][15] ), 
        .CO(\CARRYB[14][14] ), .S(\SUMB[14][14] ) );
  FA_X1 S2_14_15 ( .A(\ab[14][15] ), .B(\CARRYB[13][15] ), .CI(\SUMB[13][16] ), 
        .CO(\CARRYB[14][15] ), .S(\SUMB[14][15] ) );
  FA_X1 S2_14_16 ( .A(\ab[14][16] ), .B(\CARRYB[13][16] ), .CI(\SUMB[13][17] ), 
        .CO(\CARRYB[14][16] ), .S(\SUMB[14][16] ) );
  FA_X1 S2_14_17 ( .A(\ab[14][17] ), .B(\CARRYB[13][17] ), .CI(\SUMB[13][18] ), 
        .S(\SUMB[14][17] ) );
  FA_X1 S1_13_0 ( .A(\ab[13][0] ), .B(\CARRYB[12][0] ), .CI(\SUMB[12][1] ), 
        .CO(\CARRYB[13][0] ), .S(PRODUCT[13]) );
  FA_X1 S2_13_1 ( .A(\ab[13][1] ), .B(\CARRYB[12][1] ), .CI(\SUMB[12][2] ), 
        .CO(\CARRYB[13][1] ), .S(\SUMB[13][1] ) );
  FA_X1 S2_13_2 ( .A(\ab[13][2] ), .B(\CARRYB[12][2] ), .CI(\SUMB[12][3] ), 
        .CO(\CARRYB[13][2] ), .S(\SUMB[13][2] ) );
  FA_X1 S2_13_3 ( .A(\ab[13][3] ), .B(\CARRYB[12][3] ), .CI(\SUMB[12][4] ), 
        .CO(\CARRYB[13][3] ), .S(\SUMB[13][3] ) );
  FA_X1 S2_13_4 ( .A(\ab[13][4] ), .B(\CARRYB[12][4] ), .CI(\SUMB[12][5] ), 
        .CO(\CARRYB[13][4] ), .S(\SUMB[13][4] ) );
  FA_X1 S2_13_5 ( .A(\ab[13][5] ), .B(\CARRYB[12][5] ), .CI(\SUMB[12][6] ), 
        .CO(\CARRYB[13][5] ), .S(\SUMB[13][5] ) );
  FA_X1 S2_13_6 ( .A(\ab[13][6] ), .B(\CARRYB[12][6] ), .CI(\SUMB[12][7] ), 
        .CO(\CARRYB[13][6] ), .S(\SUMB[13][6] ) );
  FA_X1 S2_13_7 ( .A(\ab[13][7] ), .B(\CARRYB[12][7] ), .CI(\SUMB[12][8] ), 
        .CO(\CARRYB[13][7] ), .S(\SUMB[13][7] ) );
  FA_X1 S2_13_8 ( .A(\ab[13][8] ), .B(\CARRYB[12][8] ), .CI(\SUMB[12][9] ), 
        .CO(\CARRYB[13][8] ), .S(\SUMB[13][8] ) );
  FA_X1 S2_13_9 ( .A(\ab[13][9] ), .B(\CARRYB[12][9] ), .CI(\SUMB[12][10] ), 
        .CO(\CARRYB[13][9] ), .S(\SUMB[13][9] ) );
  FA_X1 S2_13_10 ( .A(\ab[13][10] ), .B(\CARRYB[12][10] ), .CI(\SUMB[12][11] ), 
        .CO(\CARRYB[13][10] ), .S(\SUMB[13][10] ) );
  FA_X1 S2_13_11 ( .A(\ab[13][11] ), .B(\CARRYB[12][11] ), .CI(\SUMB[12][12] ), 
        .CO(\CARRYB[13][11] ), .S(\SUMB[13][11] ) );
  FA_X1 S2_13_12 ( .A(\ab[13][12] ), .B(\CARRYB[12][12] ), .CI(\SUMB[12][13] ), 
        .CO(\CARRYB[13][12] ), .S(\SUMB[13][12] ) );
  FA_X1 S2_13_13 ( .A(\ab[13][13] ), .B(\CARRYB[12][13] ), .CI(\SUMB[12][14] ), 
        .CO(\CARRYB[13][13] ), .S(\SUMB[13][13] ) );
  FA_X1 S2_13_14 ( .A(\ab[13][14] ), .B(\CARRYB[12][14] ), .CI(\SUMB[12][15] ), 
        .CO(\CARRYB[13][14] ), .S(\SUMB[13][14] ) );
  FA_X1 S2_13_15 ( .A(\ab[13][15] ), .B(\CARRYB[12][15] ), .CI(\SUMB[12][16] ), 
        .CO(\CARRYB[13][15] ), .S(\SUMB[13][15] ) );
  FA_X1 S2_13_16 ( .A(\ab[13][16] ), .B(\CARRYB[12][16] ), .CI(\SUMB[12][17] ), 
        .CO(\CARRYB[13][16] ), .S(\SUMB[13][16] ) );
  FA_X1 S2_13_17 ( .A(\ab[13][17] ), .B(\CARRYB[12][17] ), .CI(\SUMB[12][18] ), 
        .CO(\CARRYB[13][17] ), .S(\SUMB[13][17] ) );
  FA_X1 S2_13_18 ( .A(\ab[13][18] ), .B(\CARRYB[12][18] ), .CI(\SUMB[12][19] ), 
        .S(\SUMB[13][18] ) );
  FA_X1 S1_12_0 ( .A(\ab[12][0] ), .B(\CARRYB[11][0] ), .CI(\SUMB[11][1] ), 
        .CO(\CARRYB[12][0] ), .S(PRODUCT[12]) );
  FA_X1 S2_12_1 ( .A(\ab[12][1] ), .B(\CARRYB[11][1] ), .CI(\SUMB[11][2] ), 
        .CO(\CARRYB[12][1] ), .S(\SUMB[12][1] ) );
  FA_X1 S2_12_2 ( .A(\ab[12][2] ), .B(\CARRYB[11][2] ), .CI(\SUMB[11][3] ), 
        .CO(\CARRYB[12][2] ), .S(\SUMB[12][2] ) );
  FA_X1 S2_12_3 ( .A(\ab[12][3] ), .B(\CARRYB[11][3] ), .CI(\SUMB[11][4] ), 
        .CO(\CARRYB[12][3] ), .S(\SUMB[12][3] ) );
  FA_X1 S2_12_4 ( .A(\ab[12][4] ), .B(\CARRYB[11][4] ), .CI(\SUMB[11][5] ), 
        .CO(\CARRYB[12][4] ), .S(\SUMB[12][4] ) );
  FA_X1 S2_12_5 ( .A(\ab[12][5] ), .B(\CARRYB[11][5] ), .CI(\SUMB[11][6] ), 
        .CO(\CARRYB[12][5] ), .S(\SUMB[12][5] ) );
  FA_X1 S2_12_6 ( .A(\ab[12][6] ), .B(\CARRYB[11][6] ), .CI(\SUMB[11][7] ), 
        .CO(\CARRYB[12][6] ), .S(\SUMB[12][6] ) );
  FA_X1 S2_12_7 ( .A(\ab[12][7] ), .B(\CARRYB[11][7] ), .CI(\SUMB[11][8] ), 
        .CO(\CARRYB[12][7] ), .S(\SUMB[12][7] ) );
  FA_X1 S2_12_8 ( .A(\ab[12][8] ), .B(\CARRYB[11][8] ), .CI(\SUMB[11][9] ), 
        .CO(\CARRYB[12][8] ), .S(\SUMB[12][8] ) );
  FA_X1 S2_12_9 ( .A(\ab[12][9] ), .B(\CARRYB[11][9] ), .CI(\SUMB[11][10] ), 
        .CO(\CARRYB[12][9] ), .S(\SUMB[12][9] ) );
  FA_X1 S2_12_10 ( .A(\ab[12][10] ), .B(\CARRYB[11][10] ), .CI(\SUMB[11][11] ), 
        .CO(\CARRYB[12][10] ), .S(\SUMB[12][10] ) );
  FA_X1 S2_12_11 ( .A(\ab[12][11] ), .B(\CARRYB[11][11] ), .CI(\SUMB[11][12] ), 
        .CO(\CARRYB[12][11] ), .S(\SUMB[12][11] ) );
  FA_X1 S2_12_12 ( .A(\ab[12][12] ), .B(\CARRYB[11][12] ), .CI(\SUMB[11][13] ), 
        .CO(\CARRYB[12][12] ), .S(\SUMB[12][12] ) );
  FA_X1 S2_12_13 ( .A(\ab[12][13] ), .B(\CARRYB[11][13] ), .CI(\SUMB[11][14] ), 
        .CO(\CARRYB[12][13] ), .S(\SUMB[12][13] ) );
  FA_X1 S2_12_14 ( .A(\ab[12][14] ), .B(\CARRYB[11][14] ), .CI(\SUMB[11][15] ), 
        .CO(\CARRYB[12][14] ), .S(\SUMB[12][14] ) );
  FA_X1 S2_12_15 ( .A(\ab[12][15] ), .B(\CARRYB[11][15] ), .CI(\SUMB[11][16] ), 
        .CO(\CARRYB[12][15] ), .S(\SUMB[12][15] ) );
  FA_X1 S2_12_16 ( .A(\ab[12][16] ), .B(\CARRYB[11][16] ), .CI(\SUMB[11][17] ), 
        .CO(\CARRYB[12][16] ), .S(\SUMB[12][16] ) );
  FA_X1 S2_12_17 ( .A(\ab[12][17] ), .B(\CARRYB[11][17] ), .CI(\SUMB[11][18] ), 
        .CO(\CARRYB[12][17] ), .S(\SUMB[12][17] ) );
  FA_X1 S2_12_18 ( .A(\ab[12][18] ), .B(\CARRYB[11][18] ), .CI(\SUMB[11][19] ), 
        .CO(\CARRYB[12][18] ), .S(\SUMB[12][18] ) );
  FA_X1 S2_12_19 ( .A(\ab[12][19] ), .B(\CARRYB[11][19] ), .CI(\SUMB[11][20] ), 
        .S(\SUMB[12][19] ) );
  FA_X1 S1_11_0 ( .A(\ab[11][0] ), .B(\CARRYB[10][0] ), .CI(\SUMB[10][1] ), 
        .CO(\CARRYB[11][0] ), .S(PRODUCT[11]) );
  FA_X1 S2_11_1 ( .A(\ab[11][1] ), .B(\CARRYB[10][1] ), .CI(\SUMB[10][2] ), 
        .CO(\CARRYB[11][1] ), .S(\SUMB[11][1] ) );
  FA_X1 S2_11_2 ( .A(\ab[11][2] ), .B(\CARRYB[10][2] ), .CI(\SUMB[10][3] ), 
        .CO(\CARRYB[11][2] ), .S(\SUMB[11][2] ) );
  FA_X1 S2_11_3 ( .A(\ab[11][3] ), .B(\CARRYB[10][3] ), .CI(\SUMB[10][4] ), 
        .CO(\CARRYB[11][3] ), .S(\SUMB[11][3] ) );
  FA_X1 S2_11_4 ( .A(\ab[11][4] ), .B(\CARRYB[10][4] ), .CI(\SUMB[10][5] ), 
        .CO(\CARRYB[11][4] ), .S(\SUMB[11][4] ) );
  FA_X1 S2_11_5 ( .A(\ab[11][5] ), .B(\CARRYB[10][5] ), .CI(\SUMB[10][6] ), 
        .CO(\CARRYB[11][5] ), .S(\SUMB[11][5] ) );
  FA_X1 S2_11_6 ( .A(\ab[11][6] ), .B(\CARRYB[10][6] ), .CI(\SUMB[10][7] ), 
        .CO(\CARRYB[11][6] ), .S(\SUMB[11][6] ) );
  FA_X1 S2_11_7 ( .A(\ab[11][7] ), .B(\CARRYB[10][7] ), .CI(\SUMB[10][8] ), 
        .CO(\CARRYB[11][7] ), .S(\SUMB[11][7] ) );
  FA_X1 S2_11_8 ( .A(\ab[11][8] ), .B(\CARRYB[10][8] ), .CI(\SUMB[10][9] ), 
        .CO(\CARRYB[11][8] ), .S(\SUMB[11][8] ) );
  FA_X1 S2_11_9 ( .A(\ab[11][9] ), .B(\CARRYB[10][9] ), .CI(\SUMB[10][10] ), 
        .CO(\CARRYB[11][9] ), .S(\SUMB[11][9] ) );
  FA_X1 S2_11_10 ( .A(\ab[11][10] ), .B(\CARRYB[10][10] ), .CI(\SUMB[10][11] ), 
        .CO(\CARRYB[11][10] ), .S(\SUMB[11][10] ) );
  FA_X1 S2_11_11 ( .A(\ab[11][11] ), .B(\CARRYB[10][11] ), .CI(\SUMB[10][12] ), 
        .CO(\CARRYB[11][11] ), .S(\SUMB[11][11] ) );
  FA_X1 S2_11_12 ( .A(\ab[11][12] ), .B(\CARRYB[10][12] ), .CI(\SUMB[10][13] ), 
        .CO(\CARRYB[11][12] ), .S(\SUMB[11][12] ) );
  FA_X1 S2_11_13 ( .A(\ab[11][13] ), .B(\CARRYB[10][13] ), .CI(\SUMB[10][14] ), 
        .CO(\CARRYB[11][13] ), .S(\SUMB[11][13] ) );
  FA_X1 S2_11_14 ( .A(\ab[11][14] ), .B(\CARRYB[10][14] ), .CI(\SUMB[10][15] ), 
        .CO(\CARRYB[11][14] ), .S(\SUMB[11][14] ) );
  FA_X1 S2_11_15 ( .A(\ab[11][15] ), .B(\CARRYB[10][15] ), .CI(\SUMB[10][16] ), 
        .CO(\CARRYB[11][15] ), .S(\SUMB[11][15] ) );
  FA_X1 S2_11_16 ( .A(\ab[11][16] ), .B(\CARRYB[10][16] ), .CI(\SUMB[10][17] ), 
        .CO(\CARRYB[11][16] ), .S(\SUMB[11][16] ) );
  FA_X1 S2_11_17 ( .A(\ab[11][17] ), .B(\CARRYB[10][17] ), .CI(\SUMB[10][18] ), 
        .CO(\CARRYB[11][17] ), .S(\SUMB[11][17] ) );
  FA_X1 S2_11_18 ( .A(\ab[11][18] ), .B(\CARRYB[10][18] ), .CI(\SUMB[10][19] ), 
        .CO(\CARRYB[11][18] ), .S(\SUMB[11][18] ) );
  FA_X1 S2_11_19 ( .A(\ab[11][19] ), .B(\CARRYB[10][19] ), .CI(\SUMB[10][20] ), 
        .CO(\CARRYB[11][19] ), .S(\SUMB[11][19] ) );
  FA_X1 S2_11_20 ( .A(\ab[11][20] ), .B(\CARRYB[10][20] ), .CI(\SUMB[10][21] ), 
        .S(\SUMB[11][20] ) );
  FA_X1 S1_10_0 ( .A(\ab[10][0] ), .B(\CARRYB[9][0] ), .CI(\SUMB[9][1] ), .CO(
        \CARRYB[10][0] ), .S(PRODUCT[10]) );
  FA_X1 S2_10_1 ( .A(\ab[10][1] ), .B(\CARRYB[9][1] ), .CI(\SUMB[9][2] ), .CO(
        \CARRYB[10][1] ), .S(\SUMB[10][1] ) );
  FA_X1 S2_10_2 ( .A(\ab[10][2] ), .B(\CARRYB[9][2] ), .CI(\SUMB[9][3] ), .CO(
        \CARRYB[10][2] ), .S(\SUMB[10][2] ) );
  FA_X1 S2_10_3 ( .A(\ab[10][3] ), .B(\CARRYB[9][3] ), .CI(\SUMB[9][4] ), .CO(
        \CARRYB[10][3] ), .S(\SUMB[10][3] ) );
  FA_X1 S2_10_4 ( .A(\ab[10][4] ), .B(\CARRYB[9][4] ), .CI(\SUMB[9][5] ), .CO(
        \CARRYB[10][4] ), .S(\SUMB[10][4] ) );
  FA_X1 S2_10_5 ( .A(\ab[10][5] ), .B(\CARRYB[9][5] ), .CI(\SUMB[9][6] ), .CO(
        \CARRYB[10][5] ), .S(\SUMB[10][5] ) );
  FA_X1 S2_10_6 ( .A(\ab[10][6] ), .B(\CARRYB[9][6] ), .CI(\SUMB[9][7] ), .CO(
        \CARRYB[10][6] ), .S(\SUMB[10][6] ) );
  FA_X1 S2_10_7 ( .A(\ab[10][7] ), .B(\CARRYB[9][7] ), .CI(\SUMB[9][8] ), .CO(
        \CARRYB[10][7] ), .S(\SUMB[10][7] ) );
  FA_X1 S2_10_8 ( .A(\ab[10][8] ), .B(\CARRYB[9][8] ), .CI(\SUMB[9][9] ), .CO(
        \CARRYB[10][8] ), .S(\SUMB[10][8] ) );
  FA_X1 S2_10_9 ( .A(\ab[10][9] ), .B(\CARRYB[9][9] ), .CI(\SUMB[9][10] ), 
        .CO(\CARRYB[10][9] ), .S(\SUMB[10][9] ) );
  FA_X1 S2_10_10 ( .A(\ab[10][10] ), .B(\CARRYB[9][10] ), .CI(\SUMB[9][11] ), 
        .CO(\CARRYB[10][10] ), .S(\SUMB[10][10] ) );
  FA_X1 S2_10_11 ( .A(\ab[10][11] ), .B(\CARRYB[9][11] ), .CI(\SUMB[9][12] ), 
        .CO(\CARRYB[10][11] ), .S(\SUMB[10][11] ) );
  FA_X1 S2_10_12 ( .A(\ab[10][12] ), .B(\CARRYB[9][12] ), .CI(\SUMB[9][13] ), 
        .CO(\CARRYB[10][12] ), .S(\SUMB[10][12] ) );
  FA_X1 S2_10_13 ( .A(\ab[10][13] ), .B(\CARRYB[9][13] ), .CI(\SUMB[9][14] ), 
        .CO(\CARRYB[10][13] ), .S(\SUMB[10][13] ) );
  FA_X1 S2_10_14 ( .A(\ab[10][14] ), .B(\CARRYB[9][14] ), .CI(\SUMB[9][15] ), 
        .CO(\CARRYB[10][14] ), .S(\SUMB[10][14] ) );
  FA_X1 S2_10_15 ( .A(\ab[10][15] ), .B(\CARRYB[9][15] ), .CI(\SUMB[9][16] ), 
        .CO(\CARRYB[10][15] ), .S(\SUMB[10][15] ) );
  FA_X1 S2_10_16 ( .A(\ab[10][16] ), .B(\CARRYB[9][16] ), .CI(\SUMB[9][17] ), 
        .CO(\CARRYB[10][16] ), .S(\SUMB[10][16] ) );
  FA_X1 S2_10_17 ( .A(\ab[10][17] ), .B(\CARRYB[9][17] ), .CI(\SUMB[9][18] ), 
        .CO(\CARRYB[10][17] ), .S(\SUMB[10][17] ) );
  FA_X1 S2_10_18 ( .A(\ab[10][18] ), .B(\CARRYB[9][18] ), .CI(\SUMB[9][19] ), 
        .CO(\CARRYB[10][18] ), .S(\SUMB[10][18] ) );
  FA_X1 S2_10_19 ( .A(\ab[10][19] ), .B(\CARRYB[9][19] ), .CI(\SUMB[9][20] ), 
        .CO(\CARRYB[10][19] ), .S(\SUMB[10][19] ) );
  FA_X1 S2_10_20 ( .A(\ab[10][20] ), .B(\CARRYB[9][20] ), .CI(\SUMB[9][21] ), 
        .CO(\CARRYB[10][20] ), .S(\SUMB[10][20] ) );
  FA_X1 S2_10_21 ( .A(\ab[10][21] ), .B(\CARRYB[9][21] ), .CI(\SUMB[9][22] ), 
        .S(\SUMB[10][21] ) );
  FA_X1 S1_9_0 ( .A(\ab[9][0] ), .B(\CARRYB[8][0] ), .CI(\SUMB[8][1] ), .CO(
        \CARRYB[9][0] ), .S(PRODUCT[9]) );
  FA_X1 S2_9_1 ( .A(\ab[9][1] ), .B(\CARRYB[8][1] ), .CI(\SUMB[8][2] ), .CO(
        \CARRYB[9][1] ), .S(\SUMB[9][1] ) );
  FA_X1 S2_9_2 ( .A(\ab[9][2] ), .B(\CARRYB[8][2] ), .CI(\SUMB[8][3] ), .CO(
        \CARRYB[9][2] ), .S(\SUMB[9][2] ) );
  FA_X1 S2_9_3 ( .A(\ab[9][3] ), .B(\CARRYB[8][3] ), .CI(\SUMB[8][4] ), .CO(
        \CARRYB[9][3] ), .S(\SUMB[9][3] ) );
  FA_X1 S2_9_4 ( .A(\ab[9][4] ), .B(\CARRYB[8][4] ), .CI(\SUMB[8][5] ), .CO(
        \CARRYB[9][4] ), .S(\SUMB[9][4] ) );
  FA_X1 S2_9_5 ( .A(\ab[9][5] ), .B(\CARRYB[8][5] ), .CI(\SUMB[8][6] ), .CO(
        \CARRYB[9][5] ), .S(\SUMB[9][5] ) );
  FA_X1 S2_9_6 ( .A(\ab[9][6] ), .B(\CARRYB[8][6] ), .CI(\SUMB[8][7] ), .CO(
        \CARRYB[9][6] ), .S(\SUMB[9][6] ) );
  FA_X1 S2_9_7 ( .A(\ab[9][7] ), .B(\CARRYB[8][7] ), .CI(\SUMB[8][8] ), .CO(
        \CARRYB[9][7] ), .S(\SUMB[9][7] ) );
  FA_X1 S2_9_8 ( .A(\ab[9][8] ), .B(\CARRYB[8][8] ), .CI(\SUMB[8][9] ), .CO(
        \CARRYB[9][8] ), .S(\SUMB[9][8] ) );
  FA_X1 S2_9_9 ( .A(\ab[9][9] ), .B(\CARRYB[8][9] ), .CI(\SUMB[8][10] ), .CO(
        \CARRYB[9][9] ), .S(\SUMB[9][9] ) );
  FA_X1 S2_9_10 ( .A(\ab[9][10] ), .B(\CARRYB[8][10] ), .CI(\SUMB[8][11] ), 
        .CO(\CARRYB[9][10] ), .S(\SUMB[9][10] ) );
  FA_X1 S2_9_11 ( .A(\ab[9][11] ), .B(\CARRYB[8][11] ), .CI(\SUMB[8][12] ), 
        .CO(\CARRYB[9][11] ), .S(\SUMB[9][11] ) );
  FA_X1 S2_9_12 ( .A(\ab[9][12] ), .B(\CARRYB[8][12] ), .CI(\SUMB[8][13] ), 
        .CO(\CARRYB[9][12] ), .S(\SUMB[9][12] ) );
  FA_X1 S2_9_13 ( .A(\ab[9][13] ), .B(\CARRYB[8][13] ), .CI(\SUMB[8][14] ), 
        .CO(\CARRYB[9][13] ), .S(\SUMB[9][13] ) );
  FA_X1 S2_9_14 ( .A(\ab[9][14] ), .B(\CARRYB[8][14] ), .CI(\SUMB[8][15] ), 
        .CO(\CARRYB[9][14] ), .S(\SUMB[9][14] ) );
  FA_X1 S2_9_15 ( .A(\ab[9][15] ), .B(\CARRYB[8][15] ), .CI(\SUMB[8][16] ), 
        .CO(\CARRYB[9][15] ), .S(\SUMB[9][15] ) );
  FA_X1 S2_9_16 ( .A(\ab[9][16] ), .B(\CARRYB[8][16] ), .CI(\SUMB[8][17] ), 
        .CO(\CARRYB[9][16] ), .S(\SUMB[9][16] ) );
  FA_X1 S2_9_17 ( .A(\ab[9][17] ), .B(\CARRYB[8][17] ), .CI(\SUMB[8][18] ), 
        .CO(\CARRYB[9][17] ), .S(\SUMB[9][17] ) );
  FA_X1 S2_9_18 ( .A(\ab[9][18] ), .B(\CARRYB[8][18] ), .CI(\SUMB[8][19] ), 
        .CO(\CARRYB[9][18] ), .S(\SUMB[9][18] ) );
  FA_X1 S2_9_19 ( .A(\ab[9][19] ), .B(\CARRYB[8][19] ), .CI(\SUMB[8][20] ), 
        .CO(\CARRYB[9][19] ), .S(\SUMB[9][19] ) );
  FA_X1 S2_9_20 ( .A(\ab[9][20] ), .B(\CARRYB[8][20] ), .CI(\SUMB[8][21] ), 
        .CO(\CARRYB[9][20] ), .S(\SUMB[9][20] ) );
  FA_X1 S2_9_21 ( .A(\ab[9][21] ), .B(\CARRYB[8][21] ), .CI(\SUMB[8][22] ), 
        .CO(\CARRYB[9][21] ), .S(\SUMB[9][21] ) );
  FA_X1 S2_9_22 ( .A(\ab[9][22] ), .B(\CARRYB[8][22] ), .CI(\SUMB[8][23] ), 
        .S(\SUMB[9][22] ) );
  FA_X1 S1_8_0 ( .A(\ab[8][0] ), .B(\CARRYB[7][0] ), .CI(\SUMB[7][1] ), .CO(
        \CARRYB[8][0] ), .S(PRODUCT[8]) );
  FA_X1 S2_8_1 ( .A(\ab[8][1] ), .B(\CARRYB[7][1] ), .CI(\SUMB[7][2] ), .CO(
        \CARRYB[8][1] ), .S(\SUMB[8][1] ) );
  FA_X1 S2_8_2 ( .A(\ab[8][2] ), .B(\CARRYB[7][2] ), .CI(\SUMB[7][3] ), .CO(
        \CARRYB[8][2] ), .S(\SUMB[8][2] ) );
  FA_X1 S2_8_3 ( .A(\ab[8][3] ), .B(\CARRYB[7][3] ), .CI(\SUMB[7][4] ), .CO(
        \CARRYB[8][3] ), .S(\SUMB[8][3] ) );
  FA_X1 S2_8_4 ( .A(\ab[8][4] ), .B(\CARRYB[7][4] ), .CI(\SUMB[7][5] ), .CO(
        \CARRYB[8][4] ), .S(\SUMB[8][4] ) );
  FA_X1 S2_8_5 ( .A(\ab[8][5] ), .B(\CARRYB[7][5] ), .CI(\SUMB[7][6] ), .CO(
        \CARRYB[8][5] ), .S(\SUMB[8][5] ) );
  FA_X1 S2_8_6 ( .A(\ab[8][6] ), .B(\CARRYB[7][6] ), .CI(\SUMB[7][7] ), .CO(
        \CARRYB[8][6] ), .S(\SUMB[8][6] ) );
  FA_X1 S2_8_7 ( .A(\ab[8][7] ), .B(\CARRYB[7][7] ), .CI(\SUMB[7][8] ), .CO(
        \CARRYB[8][7] ), .S(\SUMB[8][7] ) );
  FA_X1 S2_8_8 ( .A(\ab[8][8] ), .B(\CARRYB[7][8] ), .CI(\SUMB[7][9] ), .CO(
        \CARRYB[8][8] ), .S(\SUMB[8][8] ) );
  FA_X1 S2_8_9 ( .A(\ab[8][9] ), .B(\CARRYB[7][9] ), .CI(\SUMB[7][10] ), .CO(
        \CARRYB[8][9] ), .S(\SUMB[8][9] ) );
  FA_X1 S2_8_10 ( .A(\ab[8][10] ), .B(\CARRYB[7][10] ), .CI(\SUMB[7][11] ), 
        .CO(\CARRYB[8][10] ), .S(\SUMB[8][10] ) );
  FA_X1 S2_8_11 ( .A(\ab[8][11] ), .B(\CARRYB[7][11] ), .CI(\SUMB[7][12] ), 
        .CO(\CARRYB[8][11] ), .S(\SUMB[8][11] ) );
  FA_X1 S2_8_12 ( .A(\ab[8][12] ), .B(\CARRYB[7][12] ), .CI(\SUMB[7][13] ), 
        .CO(\CARRYB[8][12] ), .S(\SUMB[8][12] ) );
  FA_X1 S2_8_13 ( .A(\ab[8][13] ), .B(\CARRYB[7][13] ), .CI(\SUMB[7][14] ), 
        .CO(\CARRYB[8][13] ), .S(\SUMB[8][13] ) );
  FA_X1 S2_8_14 ( .A(\ab[8][14] ), .B(\CARRYB[7][14] ), .CI(\SUMB[7][15] ), 
        .CO(\CARRYB[8][14] ), .S(\SUMB[8][14] ) );
  FA_X1 S2_8_15 ( .A(\ab[8][15] ), .B(\CARRYB[7][15] ), .CI(\SUMB[7][16] ), 
        .CO(\CARRYB[8][15] ), .S(\SUMB[8][15] ) );
  FA_X1 S2_8_16 ( .A(\ab[8][16] ), .B(\CARRYB[7][16] ), .CI(\SUMB[7][17] ), 
        .CO(\CARRYB[8][16] ), .S(\SUMB[8][16] ) );
  FA_X1 S2_8_17 ( .A(\ab[8][17] ), .B(\CARRYB[7][17] ), .CI(\SUMB[7][18] ), 
        .CO(\CARRYB[8][17] ), .S(\SUMB[8][17] ) );
  FA_X1 S2_8_18 ( .A(\ab[8][18] ), .B(\CARRYB[7][18] ), .CI(\SUMB[7][19] ), 
        .CO(\CARRYB[8][18] ), .S(\SUMB[8][18] ) );
  FA_X1 S2_8_19 ( .A(\ab[8][19] ), .B(\CARRYB[7][19] ), .CI(\SUMB[7][20] ), 
        .CO(\CARRYB[8][19] ), .S(\SUMB[8][19] ) );
  FA_X1 S2_8_20 ( .A(\ab[8][20] ), .B(\CARRYB[7][20] ), .CI(\SUMB[7][21] ), 
        .CO(\CARRYB[8][20] ), .S(\SUMB[8][20] ) );
  FA_X1 S2_8_21 ( .A(\ab[8][21] ), .B(\CARRYB[7][21] ), .CI(\SUMB[7][22] ), 
        .CO(\CARRYB[8][21] ), .S(\SUMB[8][21] ) );
  FA_X1 S2_8_22 ( .A(\ab[8][22] ), .B(\CARRYB[7][22] ), .CI(\SUMB[7][23] ), 
        .CO(\CARRYB[8][22] ), .S(\SUMB[8][22] ) );
  FA_X1 S2_8_23 ( .A(\ab[8][23] ), .B(\CARRYB[7][23] ), .CI(\SUMB[7][24] ), 
        .S(\SUMB[8][23] ) );
  FA_X1 S1_7_0 ( .A(\ab[7][0] ), .B(\CARRYB[6][0] ), .CI(\SUMB[6][1] ), .CO(
        \CARRYB[7][0] ), .S(PRODUCT[7]) );
  FA_X1 S2_7_1 ( .A(\ab[7][1] ), .B(\CARRYB[6][1] ), .CI(\SUMB[6][2] ), .CO(
        \CARRYB[7][1] ), .S(\SUMB[7][1] ) );
  FA_X1 S2_7_2 ( .A(\ab[7][2] ), .B(\CARRYB[6][2] ), .CI(\SUMB[6][3] ), .CO(
        \CARRYB[7][2] ), .S(\SUMB[7][2] ) );
  FA_X1 S2_7_3 ( .A(\ab[7][3] ), .B(\CARRYB[6][3] ), .CI(\SUMB[6][4] ), .CO(
        \CARRYB[7][3] ), .S(\SUMB[7][3] ) );
  FA_X1 S2_7_4 ( .A(\ab[7][4] ), .B(\CARRYB[6][4] ), .CI(\SUMB[6][5] ), .CO(
        \CARRYB[7][4] ), .S(\SUMB[7][4] ) );
  FA_X1 S2_7_5 ( .A(\ab[7][5] ), .B(\CARRYB[6][5] ), .CI(\SUMB[6][6] ), .CO(
        \CARRYB[7][5] ), .S(\SUMB[7][5] ) );
  FA_X1 S2_7_6 ( .A(\ab[7][6] ), .B(\CARRYB[6][6] ), .CI(\SUMB[6][7] ), .CO(
        \CARRYB[7][6] ), .S(\SUMB[7][6] ) );
  FA_X1 S2_7_7 ( .A(\ab[7][7] ), .B(\CARRYB[6][7] ), .CI(\SUMB[6][8] ), .CO(
        \CARRYB[7][7] ), .S(\SUMB[7][7] ) );
  FA_X1 S2_7_8 ( .A(\ab[7][8] ), .B(\CARRYB[6][8] ), .CI(\SUMB[6][9] ), .CO(
        \CARRYB[7][8] ), .S(\SUMB[7][8] ) );
  FA_X1 S2_7_9 ( .A(\ab[7][9] ), .B(\CARRYB[6][9] ), .CI(\SUMB[6][10] ), .CO(
        \CARRYB[7][9] ), .S(\SUMB[7][9] ) );
  FA_X1 S2_7_10 ( .A(\ab[7][10] ), .B(\CARRYB[6][10] ), .CI(\SUMB[6][11] ), 
        .CO(\CARRYB[7][10] ), .S(\SUMB[7][10] ) );
  FA_X1 S2_7_11 ( .A(\ab[7][11] ), .B(\CARRYB[6][11] ), .CI(\SUMB[6][12] ), 
        .CO(\CARRYB[7][11] ), .S(\SUMB[7][11] ) );
  FA_X1 S2_7_12 ( .A(\ab[7][12] ), .B(\CARRYB[6][12] ), .CI(\SUMB[6][13] ), 
        .CO(\CARRYB[7][12] ), .S(\SUMB[7][12] ) );
  FA_X1 S2_7_13 ( .A(\ab[7][13] ), .B(\CARRYB[6][13] ), .CI(\SUMB[6][14] ), 
        .CO(\CARRYB[7][13] ), .S(\SUMB[7][13] ) );
  FA_X1 S2_7_14 ( .A(\ab[7][14] ), .B(\CARRYB[6][14] ), .CI(\SUMB[6][15] ), 
        .CO(\CARRYB[7][14] ), .S(\SUMB[7][14] ) );
  FA_X1 S2_7_15 ( .A(\ab[7][15] ), .B(\CARRYB[6][15] ), .CI(\SUMB[6][16] ), 
        .CO(\CARRYB[7][15] ), .S(\SUMB[7][15] ) );
  FA_X1 S2_7_16 ( .A(\ab[7][16] ), .B(\CARRYB[6][16] ), .CI(\SUMB[6][17] ), 
        .CO(\CARRYB[7][16] ), .S(\SUMB[7][16] ) );
  FA_X1 S2_7_17 ( .A(\ab[7][17] ), .B(\CARRYB[6][17] ), .CI(\SUMB[6][18] ), 
        .CO(\CARRYB[7][17] ), .S(\SUMB[7][17] ) );
  FA_X1 S2_7_18 ( .A(\ab[7][18] ), .B(\CARRYB[6][18] ), .CI(\SUMB[6][19] ), 
        .CO(\CARRYB[7][18] ), .S(\SUMB[7][18] ) );
  FA_X1 S2_7_19 ( .A(\ab[7][19] ), .B(\CARRYB[6][19] ), .CI(\SUMB[6][20] ), 
        .CO(\CARRYB[7][19] ), .S(\SUMB[7][19] ) );
  FA_X1 S2_7_20 ( .A(\ab[7][20] ), .B(\CARRYB[6][20] ), .CI(\SUMB[6][21] ), 
        .CO(\CARRYB[7][20] ), .S(\SUMB[7][20] ) );
  FA_X1 S2_7_21 ( .A(\ab[7][21] ), .B(\CARRYB[6][21] ), .CI(\SUMB[6][22] ), 
        .CO(\CARRYB[7][21] ), .S(\SUMB[7][21] ) );
  FA_X1 S2_7_22 ( .A(\ab[7][22] ), .B(\CARRYB[6][22] ), .CI(\SUMB[6][23] ), 
        .CO(\CARRYB[7][22] ), .S(\SUMB[7][22] ) );
  FA_X1 S2_7_23 ( .A(\ab[7][23] ), .B(\CARRYB[6][23] ), .CI(\SUMB[6][24] ), 
        .CO(\CARRYB[7][23] ), .S(\SUMB[7][23] ) );
  FA_X1 S2_7_24 ( .A(\ab[7][24] ), .B(\CARRYB[6][24] ), .CI(\SUMB[6][25] ), 
        .S(\SUMB[7][24] ) );
  FA_X1 S1_6_0 ( .A(\ab[6][0] ), .B(\CARRYB[5][0] ), .CI(\SUMB[5][1] ), .CO(
        \CARRYB[6][0] ), .S(PRODUCT[6]) );
  FA_X1 S2_6_1 ( .A(\ab[6][1] ), .B(\CARRYB[5][1] ), .CI(\SUMB[5][2] ), .CO(
        \CARRYB[6][1] ), .S(\SUMB[6][1] ) );
  FA_X1 S2_6_2 ( .A(\ab[6][2] ), .B(\CARRYB[5][2] ), .CI(\SUMB[5][3] ), .CO(
        \CARRYB[6][2] ), .S(\SUMB[6][2] ) );
  FA_X1 S2_6_3 ( .A(\ab[6][3] ), .B(\CARRYB[5][3] ), .CI(\SUMB[5][4] ), .CO(
        \CARRYB[6][3] ), .S(\SUMB[6][3] ) );
  FA_X1 S2_6_4 ( .A(\ab[6][4] ), .B(\CARRYB[5][4] ), .CI(\SUMB[5][5] ), .CO(
        \CARRYB[6][4] ), .S(\SUMB[6][4] ) );
  FA_X1 S2_6_5 ( .A(\ab[6][5] ), .B(\CARRYB[5][5] ), .CI(\SUMB[5][6] ), .CO(
        \CARRYB[6][5] ), .S(\SUMB[6][5] ) );
  FA_X1 S2_6_6 ( .A(\ab[6][6] ), .B(\CARRYB[5][6] ), .CI(\SUMB[5][7] ), .CO(
        \CARRYB[6][6] ), .S(\SUMB[6][6] ) );
  FA_X1 S2_6_7 ( .A(\ab[6][7] ), .B(\CARRYB[5][7] ), .CI(\SUMB[5][8] ), .CO(
        \CARRYB[6][7] ), .S(\SUMB[6][7] ) );
  FA_X1 S2_6_8 ( .A(\ab[6][8] ), .B(\CARRYB[5][8] ), .CI(\SUMB[5][9] ), .CO(
        \CARRYB[6][8] ), .S(\SUMB[6][8] ) );
  FA_X1 S2_6_9 ( .A(\ab[6][9] ), .B(\CARRYB[5][9] ), .CI(\SUMB[5][10] ), .CO(
        \CARRYB[6][9] ), .S(\SUMB[6][9] ) );
  FA_X1 S2_6_10 ( .A(\ab[6][10] ), .B(\CARRYB[5][10] ), .CI(\SUMB[5][11] ), 
        .CO(\CARRYB[6][10] ), .S(\SUMB[6][10] ) );
  FA_X1 S2_6_11 ( .A(\ab[6][11] ), .B(\CARRYB[5][11] ), .CI(\SUMB[5][12] ), 
        .CO(\CARRYB[6][11] ), .S(\SUMB[6][11] ) );
  FA_X1 S2_6_12 ( .A(\ab[6][12] ), .B(\CARRYB[5][12] ), .CI(\SUMB[5][13] ), 
        .CO(\CARRYB[6][12] ), .S(\SUMB[6][12] ) );
  FA_X1 S2_6_13 ( .A(\ab[6][13] ), .B(\CARRYB[5][13] ), .CI(\SUMB[5][14] ), 
        .CO(\CARRYB[6][13] ), .S(\SUMB[6][13] ) );
  FA_X1 S2_6_14 ( .A(\ab[6][14] ), .B(\CARRYB[5][14] ), .CI(\SUMB[5][15] ), 
        .CO(\CARRYB[6][14] ), .S(\SUMB[6][14] ) );
  FA_X1 S2_6_15 ( .A(\ab[6][15] ), .B(\CARRYB[5][15] ), .CI(\SUMB[5][16] ), 
        .CO(\CARRYB[6][15] ), .S(\SUMB[6][15] ) );
  FA_X1 S2_6_16 ( .A(\ab[6][16] ), .B(\CARRYB[5][16] ), .CI(\SUMB[5][17] ), 
        .CO(\CARRYB[6][16] ), .S(\SUMB[6][16] ) );
  FA_X1 S2_6_17 ( .A(\ab[6][17] ), .B(\CARRYB[5][17] ), .CI(\SUMB[5][18] ), 
        .CO(\CARRYB[6][17] ), .S(\SUMB[6][17] ) );
  FA_X1 S2_6_18 ( .A(\ab[6][18] ), .B(\CARRYB[5][18] ), .CI(\SUMB[5][19] ), 
        .CO(\CARRYB[6][18] ), .S(\SUMB[6][18] ) );
  FA_X1 S2_6_19 ( .A(\ab[6][19] ), .B(\CARRYB[5][19] ), .CI(\SUMB[5][20] ), 
        .CO(\CARRYB[6][19] ), .S(\SUMB[6][19] ) );
  FA_X1 S2_6_20 ( .A(\ab[6][20] ), .B(\CARRYB[5][20] ), .CI(\SUMB[5][21] ), 
        .CO(\CARRYB[6][20] ), .S(\SUMB[6][20] ) );
  FA_X1 S2_6_21 ( .A(\ab[6][21] ), .B(\CARRYB[5][21] ), .CI(\SUMB[5][22] ), 
        .CO(\CARRYB[6][21] ), .S(\SUMB[6][21] ) );
  FA_X1 S2_6_22 ( .A(\ab[6][22] ), .B(\CARRYB[5][22] ), .CI(\SUMB[5][23] ), 
        .CO(\CARRYB[6][22] ), .S(\SUMB[6][22] ) );
  FA_X1 S2_6_23 ( .A(\ab[6][23] ), .B(\CARRYB[5][23] ), .CI(\SUMB[5][24] ), 
        .CO(\CARRYB[6][23] ), .S(\SUMB[6][23] ) );
  FA_X1 S2_6_24 ( .A(\ab[6][24] ), .B(\CARRYB[5][24] ), .CI(\SUMB[5][25] ), 
        .CO(\CARRYB[6][24] ), .S(\SUMB[6][24] ) );
  FA_X1 S2_6_25 ( .A(\ab[6][25] ), .B(\CARRYB[5][25] ), .CI(\SUMB[5][26] ), 
        .S(\SUMB[6][25] ) );
  FA_X1 S1_5_0 ( .A(\ab[5][0] ), .B(\CARRYB[4][0] ), .CI(\SUMB[4][1] ), .CO(
        \CARRYB[5][0] ), .S(PRODUCT[5]) );
  FA_X1 S2_5_1 ( .A(\ab[5][1] ), .B(\CARRYB[4][1] ), .CI(\SUMB[4][2] ), .CO(
        \CARRYB[5][1] ), .S(\SUMB[5][1] ) );
  FA_X1 S2_5_2 ( .A(\ab[5][2] ), .B(\CARRYB[4][2] ), .CI(\SUMB[4][3] ), .CO(
        \CARRYB[5][2] ), .S(\SUMB[5][2] ) );
  FA_X1 S2_5_3 ( .A(\ab[5][3] ), .B(\CARRYB[4][3] ), .CI(\SUMB[4][4] ), .CO(
        \CARRYB[5][3] ), .S(\SUMB[5][3] ) );
  FA_X1 S2_5_4 ( .A(\ab[5][4] ), .B(\CARRYB[4][4] ), .CI(\SUMB[4][5] ), .CO(
        \CARRYB[5][4] ), .S(\SUMB[5][4] ) );
  FA_X1 S2_5_5 ( .A(\ab[5][5] ), .B(\CARRYB[4][5] ), .CI(\SUMB[4][6] ), .CO(
        \CARRYB[5][5] ), .S(\SUMB[5][5] ) );
  FA_X1 S2_5_6 ( .A(\ab[5][6] ), .B(\CARRYB[4][6] ), .CI(\SUMB[4][7] ), .CO(
        \CARRYB[5][6] ), .S(\SUMB[5][6] ) );
  FA_X1 S2_5_7 ( .A(\ab[5][7] ), .B(\CARRYB[4][7] ), .CI(\SUMB[4][8] ), .CO(
        \CARRYB[5][7] ), .S(\SUMB[5][7] ) );
  FA_X1 S2_5_8 ( .A(\ab[5][8] ), .B(\CARRYB[4][8] ), .CI(\SUMB[4][9] ), .CO(
        \CARRYB[5][8] ), .S(\SUMB[5][8] ) );
  FA_X1 S2_5_9 ( .A(\ab[5][9] ), .B(\CARRYB[4][9] ), .CI(\SUMB[4][10] ), .CO(
        \CARRYB[5][9] ), .S(\SUMB[5][9] ) );
  FA_X1 S2_5_10 ( .A(\ab[5][10] ), .B(\CARRYB[4][10] ), .CI(\SUMB[4][11] ), 
        .CO(\CARRYB[5][10] ), .S(\SUMB[5][10] ) );
  FA_X1 S2_5_11 ( .A(\ab[5][11] ), .B(\CARRYB[4][11] ), .CI(\SUMB[4][12] ), 
        .CO(\CARRYB[5][11] ), .S(\SUMB[5][11] ) );
  FA_X1 S2_5_12 ( .A(\ab[5][12] ), .B(\CARRYB[4][12] ), .CI(\SUMB[4][13] ), 
        .CO(\CARRYB[5][12] ), .S(\SUMB[5][12] ) );
  FA_X1 S2_5_13 ( .A(\ab[5][13] ), .B(\CARRYB[4][13] ), .CI(\SUMB[4][14] ), 
        .CO(\CARRYB[5][13] ), .S(\SUMB[5][13] ) );
  FA_X1 S2_5_14 ( .A(\ab[5][14] ), .B(\CARRYB[4][14] ), .CI(\SUMB[4][15] ), 
        .CO(\CARRYB[5][14] ), .S(\SUMB[5][14] ) );
  FA_X1 S2_5_15 ( .A(\ab[5][15] ), .B(\CARRYB[4][15] ), .CI(\SUMB[4][16] ), 
        .CO(\CARRYB[5][15] ), .S(\SUMB[5][15] ) );
  FA_X1 S2_5_16 ( .A(\ab[5][16] ), .B(\CARRYB[4][16] ), .CI(\SUMB[4][17] ), 
        .CO(\CARRYB[5][16] ), .S(\SUMB[5][16] ) );
  FA_X1 S2_5_17 ( .A(\ab[5][17] ), .B(\CARRYB[4][17] ), .CI(\SUMB[4][18] ), 
        .CO(\CARRYB[5][17] ), .S(\SUMB[5][17] ) );
  FA_X1 S2_5_18 ( .A(\ab[5][18] ), .B(\CARRYB[4][18] ), .CI(\SUMB[4][19] ), 
        .CO(\CARRYB[5][18] ), .S(\SUMB[5][18] ) );
  FA_X1 S2_5_19 ( .A(\ab[5][19] ), .B(\CARRYB[4][19] ), .CI(\SUMB[4][20] ), 
        .CO(\CARRYB[5][19] ), .S(\SUMB[5][19] ) );
  FA_X1 S2_5_20 ( .A(\ab[5][20] ), .B(\CARRYB[4][20] ), .CI(\SUMB[4][21] ), 
        .CO(\CARRYB[5][20] ), .S(\SUMB[5][20] ) );
  FA_X1 S2_5_21 ( .A(\ab[5][21] ), .B(\CARRYB[4][21] ), .CI(\SUMB[4][22] ), 
        .CO(\CARRYB[5][21] ), .S(\SUMB[5][21] ) );
  FA_X1 S2_5_22 ( .A(\ab[5][22] ), .B(\CARRYB[4][22] ), .CI(\SUMB[4][23] ), 
        .CO(\CARRYB[5][22] ), .S(\SUMB[5][22] ) );
  FA_X1 S2_5_23 ( .A(\ab[5][23] ), .B(\CARRYB[4][23] ), .CI(\SUMB[4][24] ), 
        .CO(\CARRYB[5][23] ), .S(\SUMB[5][23] ) );
  FA_X1 S2_5_24 ( .A(\ab[5][24] ), .B(\CARRYB[4][24] ), .CI(\SUMB[4][25] ), 
        .CO(\CARRYB[5][24] ), .S(\SUMB[5][24] ) );
  FA_X1 S2_5_25 ( .A(\ab[5][25] ), .B(\CARRYB[4][25] ), .CI(\SUMB[4][26] ), 
        .CO(\CARRYB[5][25] ), .S(\SUMB[5][25] ) );
  FA_X1 S2_5_26 ( .A(\ab[5][26] ), .B(\CARRYB[4][26] ), .CI(\SUMB[4][27] ), 
        .S(\SUMB[5][26] ) );
  FA_X1 S1_4_0 ( .A(\ab[4][0] ), .B(\CARRYB[3][0] ), .CI(\SUMB[3][1] ), .CO(
        \CARRYB[4][0] ), .S(PRODUCT[4]) );
  FA_X1 S2_4_1 ( .A(\ab[4][1] ), .B(\CARRYB[3][1] ), .CI(\SUMB[3][2] ), .CO(
        \CARRYB[4][1] ), .S(\SUMB[4][1] ) );
  FA_X1 S2_4_2 ( .A(\ab[4][2] ), .B(\CARRYB[3][2] ), .CI(\SUMB[3][3] ), .CO(
        \CARRYB[4][2] ), .S(\SUMB[4][2] ) );
  FA_X1 S2_4_3 ( .A(\ab[4][3] ), .B(\CARRYB[3][3] ), .CI(\SUMB[3][4] ), .CO(
        \CARRYB[4][3] ), .S(\SUMB[4][3] ) );
  FA_X1 S2_4_4 ( .A(\ab[4][4] ), .B(\CARRYB[3][4] ), .CI(\SUMB[3][5] ), .CO(
        \CARRYB[4][4] ), .S(\SUMB[4][4] ) );
  FA_X1 S2_4_5 ( .A(\ab[4][5] ), .B(\CARRYB[3][5] ), .CI(\SUMB[3][6] ), .CO(
        \CARRYB[4][5] ), .S(\SUMB[4][5] ) );
  FA_X1 S2_4_6 ( .A(\ab[4][6] ), .B(\CARRYB[3][6] ), .CI(\SUMB[3][7] ), .CO(
        \CARRYB[4][6] ), .S(\SUMB[4][6] ) );
  FA_X1 S2_4_7 ( .A(\ab[4][7] ), .B(\CARRYB[3][7] ), .CI(\SUMB[3][8] ), .CO(
        \CARRYB[4][7] ), .S(\SUMB[4][7] ) );
  FA_X1 S2_4_8 ( .A(\ab[4][8] ), .B(\CARRYB[3][8] ), .CI(\SUMB[3][9] ), .CO(
        \CARRYB[4][8] ), .S(\SUMB[4][8] ) );
  FA_X1 S2_4_9 ( .A(\ab[4][9] ), .B(\CARRYB[3][9] ), .CI(\SUMB[3][10] ), .CO(
        \CARRYB[4][9] ), .S(\SUMB[4][9] ) );
  FA_X1 S2_4_10 ( .A(\ab[4][10] ), .B(\CARRYB[3][10] ), .CI(\SUMB[3][11] ), 
        .CO(\CARRYB[4][10] ), .S(\SUMB[4][10] ) );
  FA_X1 S2_4_11 ( .A(\ab[4][11] ), .B(\CARRYB[3][11] ), .CI(\SUMB[3][12] ), 
        .CO(\CARRYB[4][11] ), .S(\SUMB[4][11] ) );
  FA_X1 S2_4_12 ( .A(\ab[4][12] ), .B(\CARRYB[3][12] ), .CI(\SUMB[3][13] ), 
        .CO(\CARRYB[4][12] ), .S(\SUMB[4][12] ) );
  FA_X1 S2_4_13 ( .A(\ab[4][13] ), .B(\CARRYB[3][13] ), .CI(\SUMB[3][14] ), 
        .CO(\CARRYB[4][13] ), .S(\SUMB[4][13] ) );
  FA_X1 S2_4_14 ( .A(\ab[4][14] ), .B(\CARRYB[3][14] ), .CI(\SUMB[3][15] ), 
        .CO(\CARRYB[4][14] ), .S(\SUMB[4][14] ) );
  FA_X1 S2_4_15 ( .A(\ab[4][15] ), .B(\CARRYB[3][15] ), .CI(\SUMB[3][16] ), 
        .CO(\CARRYB[4][15] ), .S(\SUMB[4][15] ) );
  FA_X1 S2_4_16 ( .A(\ab[4][16] ), .B(\CARRYB[3][16] ), .CI(\SUMB[3][17] ), 
        .CO(\CARRYB[4][16] ), .S(\SUMB[4][16] ) );
  FA_X1 S2_4_17 ( .A(\ab[4][17] ), .B(\CARRYB[3][17] ), .CI(\SUMB[3][18] ), 
        .CO(\CARRYB[4][17] ), .S(\SUMB[4][17] ) );
  FA_X1 S2_4_18 ( .A(\ab[4][18] ), .B(\CARRYB[3][18] ), .CI(\SUMB[3][19] ), 
        .CO(\CARRYB[4][18] ), .S(\SUMB[4][18] ) );
  FA_X1 S2_4_19 ( .A(\ab[4][19] ), .B(\CARRYB[3][19] ), .CI(\SUMB[3][20] ), 
        .CO(\CARRYB[4][19] ), .S(\SUMB[4][19] ) );
  FA_X1 S2_4_20 ( .A(\ab[4][20] ), .B(\CARRYB[3][20] ), .CI(\SUMB[3][21] ), 
        .CO(\CARRYB[4][20] ), .S(\SUMB[4][20] ) );
  FA_X1 S2_4_21 ( .A(\ab[4][21] ), .B(\CARRYB[3][21] ), .CI(\SUMB[3][22] ), 
        .CO(\CARRYB[4][21] ), .S(\SUMB[4][21] ) );
  FA_X1 S2_4_22 ( .A(\ab[4][22] ), .B(\CARRYB[3][22] ), .CI(\SUMB[3][23] ), 
        .CO(\CARRYB[4][22] ), .S(\SUMB[4][22] ) );
  FA_X1 S2_4_23 ( .A(\ab[4][23] ), .B(\CARRYB[3][23] ), .CI(\SUMB[3][24] ), 
        .CO(\CARRYB[4][23] ), .S(\SUMB[4][23] ) );
  FA_X1 S2_4_24 ( .A(\ab[4][24] ), .B(\CARRYB[3][24] ), .CI(\SUMB[3][25] ), 
        .CO(\CARRYB[4][24] ), .S(\SUMB[4][24] ) );
  FA_X1 S2_4_25 ( .A(\ab[4][25] ), .B(\CARRYB[3][25] ), .CI(\SUMB[3][26] ), 
        .CO(\CARRYB[4][25] ), .S(\SUMB[4][25] ) );
  FA_X1 S2_4_26 ( .A(\ab[4][26] ), .B(\CARRYB[3][26] ), .CI(\SUMB[3][27] ), 
        .CO(\CARRYB[4][26] ), .S(\SUMB[4][26] ) );
  FA_X1 S2_4_27 ( .A(\ab[4][27] ), .B(\CARRYB[3][27] ), .CI(\SUMB[3][28] ), 
        .S(\SUMB[4][27] ) );
  FA_X1 S1_3_0 ( .A(\ab[3][0] ), .B(\CARRYB[2][0] ), .CI(\SUMB[2][1] ), .CO(
        \CARRYB[3][0] ), .S(PRODUCT[3]) );
  FA_X1 S2_3_1 ( .A(\ab[3][1] ), .B(\CARRYB[2][1] ), .CI(\SUMB[2][2] ), .CO(
        \CARRYB[3][1] ), .S(\SUMB[3][1] ) );
  FA_X1 S2_3_2 ( .A(\ab[3][2] ), .B(\CARRYB[2][2] ), .CI(\SUMB[2][3] ), .CO(
        \CARRYB[3][2] ), .S(\SUMB[3][2] ) );
  FA_X1 S2_3_3 ( .A(\ab[3][3] ), .B(\CARRYB[2][3] ), .CI(\SUMB[2][4] ), .CO(
        \CARRYB[3][3] ), .S(\SUMB[3][3] ) );
  FA_X1 S2_3_4 ( .A(\ab[3][4] ), .B(\CARRYB[2][4] ), .CI(\SUMB[2][5] ), .CO(
        \CARRYB[3][4] ), .S(\SUMB[3][4] ) );
  FA_X1 S2_3_5 ( .A(\ab[3][5] ), .B(\CARRYB[2][5] ), .CI(\SUMB[2][6] ), .CO(
        \CARRYB[3][5] ), .S(\SUMB[3][5] ) );
  FA_X1 S2_3_6 ( .A(\ab[3][6] ), .B(\CARRYB[2][6] ), .CI(\SUMB[2][7] ), .CO(
        \CARRYB[3][6] ), .S(\SUMB[3][6] ) );
  FA_X1 S2_3_7 ( .A(\ab[3][7] ), .B(\CARRYB[2][7] ), .CI(\SUMB[2][8] ), .CO(
        \CARRYB[3][7] ), .S(\SUMB[3][7] ) );
  FA_X1 S2_3_8 ( .A(\ab[3][8] ), .B(\CARRYB[2][8] ), .CI(\SUMB[2][9] ), .CO(
        \CARRYB[3][8] ), .S(\SUMB[3][8] ) );
  FA_X1 S2_3_9 ( .A(\ab[3][9] ), .B(\CARRYB[2][9] ), .CI(\SUMB[2][10] ), .CO(
        \CARRYB[3][9] ), .S(\SUMB[3][9] ) );
  FA_X1 S2_3_10 ( .A(\ab[3][10] ), .B(\CARRYB[2][10] ), .CI(\SUMB[2][11] ), 
        .CO(\CARRYB[3][10] ), .S(\SUMB[3][10] ) );
  FA_X1 S2_3_11 ( .A(\ab[3][11] ), .B(\CARRYB[2][11] ), .CI(\SUMB[2][12] ), 
        .CO(\CARRYB[3][11] ), .S(\SUMB[3][11] ) );
  FA_X1 S2_3_12 ( .A(\ab[3][12] ), .B(\CARRYB[2][12] ), .CI(\SUMB[2][13] ), 
        .CO(\CARRYB[3][12] ), .S(\SUMB[3][12] ) );
  FA_X1 S2_3_13 ( .A(\ab[3][13] ), .B(\CARRYB[2][13] ), .CI(\SUMB[2][14] ), 
        .CO(\CARRYB[3][13] ), .S(\SUMB[3][13] ) );
  FA_X1 S2_3_14 ( .A(\ab[3][14] ), .B(\CARRYB[2][14] ), .CI(\SUMB[2][15] ), 
        .CO(\CARRYB[3][14] ), .S(\SUMB[3][14] ) );
  FA_X1 S2_3_15 ( .A(\ab[3][15] ), .B(\CARRYB[2][15] ), .CI(\SUMB[2][16] ), 
        .CO(\CARRYB[3][15] ), .S(\SUMB[3][15] ) );
  FA_X1 S2_3_16 ( .A(\ab[3][16] ), .B(\CARRYB[2][16] ), .CI(\SUMB[2][17] ), 
        .CO(\CARRYB[3][16] ), .S(\SUMB[3][16] ) );
  FA_X1 S2_3_17 ( .A(\ab[3][17] ), .B(\CARRYB[2][17] ), .CI(\SUMB[2][18] ), 
        .CO(\CARRYB[3][17] ), .S(\SUMB[3][17] ) );
  FA_X1 S2_3_18 ( .A(\ab[3][18] ), .B(\CARRYB[2][18] ), .CI(\SUMB[2][19] ), 
        .CO(\CARRYB[3][18] ), .S(\SUMB[3][18] ) );
  FA_X1 S2_3_19 ( .A(\ab[3][19] ), .B(\CARRYB[2][19] ), .CI(\SUMB[2][20] ), 
        .CO(\CARRYB[3][19] ), .S(\SUMB[3][19] ) );
  FA_X1 S2_3_20 ( .A(\ab[3][20] ), .B(\CARRYB[2][20] ), .CI(\SUMB[2][21] ), 
        .CO(\CARRYB[3][20] ), .S(\SUMB[3][20] ) );
  FA_X1 S2_3_21 ( .A(\ab[3][21] ), .B(\CARRYB[2][21] ), .CI(\SUMB[2][22] ), 
        .CO(\CARRYB[3][21] ), .S(\SUMB[3][21] ) );
  FA_X1 S2_3_22 ( .A(\ab[3][22] ), .B(\CARRYB[2][22] ), .CI(\SUMB[2][23] ), 
        .CO(\CARRYB[3][22] ), .S(\SUMB[3][22] ) );
  FA_X1 S2_3_23 ( .A(\ab[3][23] ), .B(\CARRYB[2][23] ), .CI(\SUMB[2][24] ), 
        .CO(\CARRYB[3][23] ), .S(\SUMB[3][23] ) );
  FA_X1 S2_3_24 ( .A(\ab[3][24] ), .B(\CARRYB[2][24] ), .CI(\SUMB[2][25] ), 
        .CO(\CARRYB[3][24] ), .S(\SUMB[3][24] ) );
  FA_X1 S2_3_25 ( .A(\ab[3][25] ), .B(\CARRYB[2][25] ), .CI(\SUMB[2][26] ), 
        .CO(\CARRYB[3][25] ), .S(\SUMB[3][25] ) );
  FA_X1 S2_3_26 ( .A(\ab[3][26] ), .B(\CARRYB[2][26] ), .CI(\SUMB[2][27] ), 
        .CO(\CARRYB[3][26] ), .S(\SUMB[3][26] ) );
  FA_X1 S2_3_27 ( .A(\ab[3][27] ), .B(\CARRYB[2][27] ), .CI(\SUMB[2][28] ), 
        .CO(\CARRYB[3][27] ), .S(\SUMB[3][27] ) );
  FA_X1 S2_3_28 ( .A(\ab[3][28] ), .B(\CARRYB[2][28] ), .CI(\SUMB[2][29] ), 
        .S(\SUMB[3][28] ) );
  FA_X1 S1_2_0 ( .A(\ab[2][0] ), .B(n27), .CI(n60), .CO(\CARRYB[2][0] ), .S(
        PRODUCT[2]) );
  FA_X1 S2_2_1 ( .A(\ab[2][1] ), .B(n26), .CI(n59), .CO(\CARRYB[2][1] ), .S(
        \SUMB[2][1] ) );
  FA_X1 S2_2_2 ( .A(\ab[2][2] ), .B(n25), .CI(n58), .CO(\CARRYB[2][2] ), .S(
        \SUMB[2][2] ) );
  FA_X1 S2_2_3 ( .A(\ab[2][3] ), .B(n24), .CI(n57), .CO(\CARRYB[2][3] ), .S(
        \SUMB[2][3] ) );
  FA_X1 S2_2_4 ( .A(\ab[2][4] ), .B(n23), .CI(n56), .CO(\CARRYB[2][4] ), .S(
        \SUMB[2][4] ) );
  FA_X1 S2_2_5 ( .A(\ab[2][5] ), .B(n22), .CI(n55), .CO(\CARRYB[2][5] ), .S(
        \SUMB[2][5] ) );
  FA_X1 S2_2_6 ( .A(\ab[2][6] ), .B(n21), .CI(n54), .CO(\CARRYB[2][6] ), .S(
        \SUMB[2][6] ) );
  FA_X1 S2_2_7 ( .A(\ab[2][7] ), .B(n20), .CI(n48), .CO(\CARRYB[2][7] ), .S(
        \SUMB[2][7] ) );
  FA_X1 S2_2_8 ( .A(\ab[2][8] ), .B(n10), .CI(n49), .CO(\CARRYB[2][8] ), .S(
        \SUMB[2][8] ) );
  FA_X1 S2_2_9 ( .A(\ab[2][9] ), .B(n11), .CI(n50), .CO(\CARRYB[2][9] ), .S(
        \SUMB[2][9] ) );
  FA_X1 S2_2_10 ( .A(\ab[2][10] ), .B(n12), .CI(n51), .CO(\CARRYB[2][10] ), 
        .S(\SUMB[2][10] ) );
  FA_X1 S2_2_11 ( .A(\ab[2][11] ), .B(n13), .CI(n52), .CO(\CARRYB[2][11] ), 
        .S(\SUMB[2][11] ) );
  FA_X1 S2_2_12 ( .A(\ab[2][12] ), .B(n14), .CI(n53), .CO(\CARRYB[2][12] ), 
        .S(\SUMB[2][12] ) );
  FA_X1 S2_2_13 ( .A(\ab[2][13] ), .B(n47), .CI(n31), .CO(\CARRYB[2][13] ), 
        .S(\SUMB[2][13] ) );
  FA_X1 S2_2_14 ( .A(\ab[2][14] ), .B(n15), .CI(n32), .CO(\CARRYB[2][14] ), 
        .S(\SUMB[2][14] ) );
  FA_X1 S2_2_15 ( .A(\ab[2][15] ), .B(n16), .CI(n33), .CO(\CARRYB[2][15] ), 
        .S(\SUMB[2][15] ) );
  FA_X1 S2_2_16 ( .A(\ab[2][16] ), .B(n17), .CI(n34), .CO(\CARRYB[2][16] ), 
        .S(\SUMB[2][16] ) );
  FA_X1 S2_2_17 ( .A(\ab[2][17] ), .B(n18), .CI(n35), .CO(\CARRYB[2][17] ), 
        .S(\SUMB[2][17] ) );
  FA_X1 S2_2_18 ( .A(\ab[2][18] ), .B(n19), .CI(n36), .CO(\CARRYB[2][18] ), 
        .S(\SUMB[2][18] ) );
  FA_X1 S2_2_19 ( .A(\ab[2][19] ), .B(n28), .CI(n37), .CO(\CARRYB[2][19] ), 
        .S(\SUMB[2][19] ) );
  FA_X1 S2_2_20 ( .A(\ab[2][20] ), .B(n29), .CI(n38), .CO(\CARRYB[2][20] ), 
        .S(\SUMB[2][20] ) );
  FA_X1 S2_2_21 ( .A(\ab[2][21] ), .B(n30), .CI(n39), .CO(\CARRYB[2][21] ), 
        .S(\SUMB[2][21] ) );
  FA_X1 S2_2_22 ( .A(\ab[2][22] ), .B(n3), .CI(n45), .CO(\CARRYB[2][22] ), .S(
        \SUMB[2][22] ) );
  FA_X1 S2_2_23 ( .A(\ab[2][23] ), .B(n9), .CI(n44), .CO(\CARRYB[2][23] ), .S(
        \SUMB[2][23] ) );
  FA_X1 S2_2_24 ( .A(\ab[2][24] ), .B(n8), .CI(n43), .CO(\CARRYB[2][24] ), .S(
        \SUMB[2][24] ) );
  FA_X1 S2_2_25 ( .A(\ab[2][25] ), .B(n7), .CI(n42), .CO(\CARRYB[2][25] ), .S(
        \SUMB[2][25] ) );
  FA_X1 S2_2_26 ( .A(\ab[2][26] ), .B(n6), .CI(n41), .CO(\CARRYB[2][26] ), .S(
        \SUMB[2][26] ) );
  FA_X1 S2_2_27 ( .A(\ab[2][27] ), .B(n5), .CI(n40), .CO(\CARRYB[2][27] ), .S(
        \SUMB[2][27] ) );
  FA_X1 S2_2_28 ( .A(\ab[2][28] ), .B(n4), .CI(n46), .CO(\CARRYB[2][28] ), .S(
        \SUMB[2][28] ) );
  FA_X1 S2_2_29 ( .A(\ab[2][29] ), .B(n62), .CI(n63), .S(\SUMB[2][29] ) );
  AND2_X1 U2 ( .A1(\ab[0][23] ), .A2(\ab[1][22] ), .ZN(n3) );
  AND2_X1 U3 ( .A1(\ab[0][29] ), .A2(\ab[1][28] ), .ZN(n4) );
  AND2_X1 U4 ( .A1(\ab[0][28] ), .A2(\ab[1][27] ), .ZN(n5) );
  AND2_X1 U5 ( .A1(\ab[0][27] ), .A2(\ab[1][26] ), .ZN(n6) );
  AND2_X1 U6 ( .A1(\ab[0][26] ), .A2(\ab[1][25] ), .ZN(n7) );
  AND2_X1 U7 ( .A1(\ab[0][25] ), .A2(\ab[1][24] ), .ZN(n8) );
  AND2_X1 U8 ( .A1(\ab[0][24] ), .A2(\ab[1][23] ), .ZN(n9) );
  AND2_X1 U9 ( .A1(\ab[0][9] ), .A2(\ab[1][8] ), .ZN(n10) );
  AND2_X1 U10 ( .A1(\ab[0][10] ), .A2(\ab[1][9] ), .ZN(n11) );
  AND2_X1 U11 ( .A1(\ab[0][11] ), .A2(\ab[1][10] ), .ZN(n12) );
  AND2_X1 U12 ( .A1(\ab[0][12] ), .A2(\ab[1][11] ), .ZN(n13) );
  AND2_X1 U13 ( .A1(\ab[0][13] ), .A2(\ab[1][12] ), .ZN(n14) );
  AND2_X1 U14 ( .A1(\ab[0][15] ), .A2(\ab[1][14] ), .ZN(n15) );
  AND2_X1 U15 ( .A1(\ab[0][16] ), .A2(\ab[1][15] ), .ZN(n16) );
  AND2_X1 U16 ( .A1(\ab[0][17] ), .A2(\ab[1][16] ), .ZN(n17) );
  AND2_X1 U17 ( .A1(\ab[0][18] ), .A2(\ab[1][17] ), .ZN(n18) );
  AND2_X1 U18 ( .A1(\ab[0][19] ), .A2(\ab[1][18] ), .ZN(n19) );
  AND2_X1 U19 ( .A1(\ab[0][8] ), .A2(\ab[1][7] ), .ZN(n20) );
  AND2_X1 U20 ( .A1(\ab[0][7] ), .A2(\ab[1][6] ), .ZN(n21) );
  AND2_X1 U21 ( .A1(\ab[0][6] ), .A2(\ab[1][5] ), .ZN(n22) );
  AND2_X1 U22 ( .A1(\ab[0][5] ), .A2(\ab[1][4] ), .ZN(n23) );
  AND2_X1 U23 ( .A1(\ab[0][4] ), .A2(\ab[1][3] ), .ZN(n24) );
  AND2_X1 U24 ( .A1(\ab[0][3] ), .A2(\ab[1][2] ), .ZN(n25) );
  AND2_X1 U25 ( .A1(\ab[0][2] ), .A2(\ab[1][1] ), .ZN(n26) );
  AND2_X1 U26 ( .A1(\ab[0][1] ), .A2(\ab[1][0] ), .ZN(n27) );
  AND2_X1 U27 ( .A1(\ab[0][20] ), .A2(\ab[1][19] ), .ZN(n28) );
  AND2_X1 U28 ( .A1(\ab[0][21] ), .A2(\ab[1][20] ), .ZN(n29) );
  AND2_X1 U29 ( .A1(\ab[0][22] ), .A2(\ab[1][21] ), .ZN(n30) );
  XOR2_X1 U30 ( .A(\ab[1][14] ), .B(\ab[0][15] ), .Z(n31) );
  XOR2_X1 U31 ( .A(\ab[1][15] ), .B(\ab[0][16] ), .Z(n32) );
  XOR2_X1 U32 ( .A(\ab[1][16] ), .B(\ab[0][17] ), .Z(n33) );
  XOR2_X1 U33 ( .A(\ab[1][17] ), .B(\ab[0][18] ), .Z(n34) );
  XOR2_X1 U34 ( .A(\ab[1][18] ), .B(\ab[0][19] ), .Z(n35) );
  XOR2_X1 U35 ( .A(\ab[1][19] ), .B(\ab[0][20] ), .Z(n36) );
  XOR2_X1 U36 ( .A(\ab[1][20] ), .B(\ab[0][21] ), .Z(n37) );
  XOR2_X1 U37 ( .A(\ab[1][21] ), .B(\ab[0][22] ), .Z(n38) );
  XOR2_X1 U38 ( .A(\ab[1][22] ), .B(\ab[0][23] ), .Z(n39) );
  XOR2_X1 U39 ( .A(\ab[1][28] ), .B(\ab[0][29] ), .Z(n40) );
  XOR2_X1 U40 ( .A(\ab[1][27] ), .B(\ab[0][28] ), .Z(n41) );
  XOR2_X1 U41 ( .A(\ab[1][26] ), .B(\ab[0][27] ), .Z(n42) );
  XOR2_X1 U42 ( .A(\ab[1][25] ), .B(\ab[0][26] ), .Z(n43) );
  XOR2_X1 U43 ( .A(\ab[1][24] ), .B(\ab[0][25] ), .Z(n44) );
  XOR2_X1 U44 ( .A(\ab[1][23] ), .B(\ab[0][24] ), .Z(n45) );
  XOR2_X1 U45 ( .A(\ab[1][29] ), .B(\ab[0][30] ), .Z(n46) );
  AND2_X1 U46 ( .A1(\ab[0][14] ), .A2(\ab[1][13] ), .ZN(n47) );
  XOR2_X1 U47 ( .A(\ab[1][8] ), .B(\ab[0][9] ), .Z(n48) );
  XOR2_X1 U48 ( .A(\ab[1][9] ), .B(\ab[0][10] ), .Z(n49) );
  XOR2_X1 U49 ( .A(\ab[1][10] ), .B(\ab[0][11] ), .Z(n50) );
  XOR2_X1 U50 ( .A(\ab[1][11] ), .B(\ab[0][12] ), .Z(n51) );
  XOR2_X1 U51 ( .A(\ab[1][12] ), .B(\ab[0][13] ), .Z(n52) );
  XOR2_X1 U52 ( .A(\ab[1][13] ), .B(\ab[0][14] ), .Z(n53) );
  XOR2_X1 U53 ( .A(\ab[1][7] ), .B(\ab[0][8] ), .Z(n54) );
  XOR2_X1 U54 ( .A(\ab[1][6] ), .B(\ab[0][7] ), .Z(n55) );
  XOR2_X1 U55 ( .A(\ab[1][5] ), .B(\ab[0][6] ), .Z(n56) );
  XOR2_X1 U56 ( .A(\ab[1][4] ), .B(\ab[0][5] ), .Z(n57) );
  XOR2_X1 U57 ( .A(\ab[1][3] ), .B(\ab[0][4] ), .Z(n58) );
  XOR2_X1 U58 ( .A(\ab[1][2] ), .B(\ab[0][3] ), .Z(n59) );
  XOR2_X1 U59 ( .A(\ab[1][1] ), .B(\ab[0][2] ), .Z(n60) );
  XOR2_X1 U60 ( .A(\ab[1][0] ), .B(\ab[0][1] ), .Z(PRODUCT[1]) );
  BUF_X1 U61 ( .A(n133), .Z(n73) );
  BUF_X1 U62 ( .A(n134), .Z(n74) );
  BUF_X1 U63 ( .A(n104), .Z(n66) );
  BUF_X1 U64 ( .A(n103), .Z(n65) );
  BUF_X1 U65 ( .A(n105), .Z(n67) );
  BUF_X1 U66 ( .A(n76), .Z(n64) );
  BUF_X1 U67 ( .A(n106), .Z(n68) );
  INV_X1 U68 ( .A(A[31]), .ZN(n99) );
  AND2_X1 U69 ( .A1(\ab[0][30] ), .A2(\ab[1][29] ), .ZN(n62) );
  BUF_X1 U70 ( .A(n118), .Z(n70) );
  BUF_X1 U71 ( .A(n132), .Z(n72) );
  INV_X1 U72 ( .A(A[0]), .ZN(n104) );
  INV_X1 U73 ( .A(B[6]), .ZN(n135) );
  INV_X1 U74 ( .A(B[5]), .ZN(n134) );
  INV_X1 U75 ( .A(B[4]), .ZN(n133) );
  INV_X1 U76 ( .A(B[1]), .ZN(n118) );
  INV_X1 U77 ( .A(A[1]), .ZN(n103) );
  INV_X1 U78 ( .A(A[3]), .ZN(n105) );
  INV_X1 U79 ( .A(A[4]), .ZN(n76) );
  INV_X1 U80 ( .A(A[5]), .ZN(n75) );
  INV_X1 U81 ( .A(A[2]), .ZN(n106) );
  INV_X1 U82 ( .A(B[7]), .ZN(n136) );
  XOR2_X1 U83 ( .A(\ab[0][31] ), .B(\ab[1][30] ), .Z(n63) );
  INV_X1 U84 ( .A(A[9]), .ZN(n80) );
  INV_X1 U85 ( .A(A[11]), .ZN(n82) );
  INV_X1 U86 ( .A(A[12]), .ZN(n89) );
  INV_X1 U87 ( .A(A[13]), .ZN(n88) );
  INV_X1 U88 ( .A(A[14]), .ZN(n87) );
  BUF_X1 U89 ( .A(n107), .Z(n69) );
  BUF_X1 U90 ( .A(n129), .Z(n71) );
  INV_X1 U91 ( .A(A[10]), .ZN(n81) );
  INV_X1 U92 ( .A(A[6]), .ZN(n77) );
  INV_X1 U93 ( .A(A[7]), .ZN(n78) );
  INV_X1 U94 ( .A(A[8]), .ZN(n79) );
  INV_X1 U95 ( .A(A[15]), .ZN(n90) );
  INV_X1 U96 ( .A(A[16]), .ZN(n85) );
  INV_X1 U97 ( .A(A[17]), .ZN(n84) );
  INV_X1 U98 ( .A(A[18]), .ZN(n83) );
  INV_X1 U99 ( .A(A[19]), .ZN(n86) );
  INV_X1 U100 ( .A(A[20]), .ZN(n97) );
  INV_X1 U101 ( .A(A[21]), .ZN(n96) );
  INV_X1 U102 ( .A(A[22]), .ZN(n95) );
  INV_X1 U103 ( .A(A[23]), .ZN(n98) );
  INV_X1 U104 ( .A(A[24]), .ZN(n91) );
  INV_X1 U105 ( .A(A[25]), .ZN(n92) );
  INV_X1 U106 ( .A(A[26]), .ZN(n93) );
  INV_X1 U107 ( .A(A[27]), .ZN(n94) );
  INV_X1 U108 ( .A(A[28]), .ZN(n102) );
  INV_X1 U109 ( .A(A[29]), .ZN(n101) );
  INV_X1 U110 ( .A(A[30]), .ZN(n100) );
  INV_X1 U111 ( .A(B[9]), .ZN(n138) );
  INV_X1 U112 ( .A(B[11]), .ZN(n109) );
  INV_X1 U113 ( .A(B[12]), .ZN(n110) );
  INV_X1 U114 ( .A(B[13]), .ZN(n111) );
  INV_X1 U115 ( .A(B[14]), .ZN(n112) );
  INV_X1 U116 ( .A(B[15]), .ZN(n113) );
  INV_X1 U117 ( .A(B[17]), .ZN(n115) );
  INV_X1 U118 ( .A(B[18]), .ZN(n116) );
  INV_X1 U119 ( .A(B[19]), .ZN(n117) );
  INV_X1 U120 ( .A(B[20]), .ZN(n119) );
  INV_X1 U121 ( .A(B[21]), .ZN(n120) );
  INV_X1 U122 ( .A(B[23]), .ZN(n122) );
  INV_X1 U123 ( .A(B[25]), .ZN(n124) );
  INV_X1 U124 ( .A(B[26]), .ZN(n125) );
  INV_X1 U125 ( .A(B[27]), .ZN(n126) );
  INV_X1 U126 ( .A(B[16]), .ZN(n114) );
  INV_X1 U127 ( .A(B[10]), .ZN(n108) );
  INV_X1 U128 ( .A(B[24]), .ZN(n123) );
  INV_X1 U129 ( .A(B[22]), .ZN(n121) );
  INV_X1 U130 ( .A(B[28]), .ZN(n127) );
  INV_X1 U131 ( .A(B[29]), .ZN(n128) );
  INV_X1 U132 ( .A(B[3]), .ZN(n132) );
  INV_X1 U133 ( .A(B[2]), .ZN(n129) );
  INV_X1 U134 ( .A(B[8]), .ZN(n137) );
  INV_X1 U135 ( .A(B[30]), .ZN(n130) );
  INV_X1 U136 ( .A(B[31]), .ZN(n131) );
  INV_X1 U137 ( .A(B[0]), .ZN(n107) );
  NOR2_X1 U138 ( .A1(n80), .A2(n138), .ZN(\ab[9][9] ) );
  NOR2_X1 U139 ( .A1(n80), .A2(n137), .ZN(\ab[9][8] ) );
  NOR2_X1 U140 ( .A1(n80), .A2(n136), .ZN(\ab[9][7] ) );
  NOR2_X1 U141 ( .A1(n80), .A2(n135), .ZN(\ab[9][6] ) );
  NOR2_X1 U142 ( .A1(n80), .A2(n134), .ZN(\ab[9][5] ) );
  NOR2_X1 U143 ( .A1(n80), .A2(n133), .ZN(\ab[9][4] ) );
  NOR2_X1 U144 ( .A1(n80), .A2(n132), .ZN(\ab[9][3] ) );
  NOR2_X1 U145 ( .A1(n80), .A2(n71), .ZN(\ab[9][2] ) );
  NOR2_X1 U146 ( .A1(n80), .A2(n121), .ZN(\ab[9][22] ) );
  NOR2_X1 U147 ( .A1(n80), .A2(n120), .ZN(\ab[9][21] ) );
  NOR2_X1 U148 ( .A1(n80), .A2(n119), .ZN(\ab[9][20] ) );
  NOR2_X1 U149 ( .A1(n80), .A2(n118), .ZN(\ab[9][1] ) );
  NOR2_X1 U150 ( .A1(n80), .A2(n117), .ZN(\ab[9][19] ) );
  NOR2_X1 U151 ( .A1(n80), .A2(n116), .ZN(\ab[9][18] ) );
  NOR2_X1 U152 ( .A1(n80), .A2(n115), .ZN(\ab[9][17] ) );
  NOR2_X1 U153 ( .A1(n80), .A2(n114), .ZN(\ab[9][16] ) );
  NOR2_X1 U154 ( .A1(n80), .A2(n113), .ZN(\ab[9][15] ) );
  NOR2_X1 U155 ( .A1(n80), .A2(n112), .ZN(\ab[9][14] ) );
  NOR2_X1 U156 ( .A1(n80), .A2(n111), .ZN(\ab[9][13] ) );
  NOR2_X1 U157 ( .A1(n80), .A2(n110), .ZN(\ab[9][12] ) );
  NOR2_X1 U158 ( .A1(n80), .A2(n109), .ZN(\ab[9][11] ) );
  NOR2_X1 U159 ( .A1(n80), .A2(n108), .ZN(\ab[9][10] ) );
  NOR2_X1 U160 ( .A1(n80), .A2(n69), .ZN(\ab[9][0] ) );
  NOR2_X1 U161 ( .A1(n138), .A2(n79), .ZN(\ab[8][9] ) );
  NOR2_X1 U162 ( .A1(n137), .A2(n79), .ZN(\ab[8][8] ) );
  NOR2_X1 U163 ( .A1(n136), .A2(n79), .ZN(\ab[8][7] ) );
  NOR2_X1 U164 ( .A1(n135), .A2(n79), .ZN(\ab[8][6] ) );
  NOR2_X1 U165 ( .A1(n134), .A2(n79), .ZN(\ab[8][5] ) );
  NOR2_X1 U166 ( .A1(n133), .A2(n79), .ZN(\ab[8][4] ) );
  NOR2_X1 U167 ( .A1(n132), .A2(n79), .ZN(\ab[8][3] ) );
  NOR2_X1 U168 ( .A1(n71), .A2(n79), .ZN(\ab[8][2] ) );
  NOR2_X1 U169 ( .A1(n122), .A2(n79), .ZN(\ab[8][23] ) );
  NOR2_X1 U170 ( .A1(n121), .A2(n79), .ZN(\ab[8][22] ) );
  NOR2_X1 U171 ( .A1(n120), .A2(n79), .ZN(\ab[8][21] ) );
  NOR2_X1 U172 ( .A1(n119), .A2(n79), .ZN(\ab[8][20] ) );
  NOR2_X1 U173 ( .A1(n118), .A2(n79), .ZN(\ab[8][1] ) );
  NOR2_X1 U174 ( .A1(n117), .A2(n79), .ZN(\ab[8][19] ) );
  NOR2_X1 U175 ( .A1(n116), .A2(n79), .ZN(\ab[8][18] ) );
  NOR2_X1 U176 ( .A1(n115), .A2(n79), .ZN(\ab[8][17] ) );
  NOR2_X1 U177 ( .A1(n114), .A2(n79), .ZN(\ab[8][16] ) );
  NOR2_X1 U178 ( .A1(n113), .A2(n79), .ZN(\ab[8][15] ) );
  NOR2_X1 U179 ( .A1(n112), .A2(n79), .ZN(\ab[8][14] ) );
  NOR2_X1 U180 ( .A1(n111), .A2(n79), .ZN(\ab[8][13] ) );
  NOR2_X1 U181 ( .A1(n110), .A2(n79), .ZN(\ab[8][12] ) );
  NOR2_X1 U182 ( .A1(n109), .A2(n79), .ZN(\ab[8][11] ) );
  NOR2_X1 U183 ( .A1(n108), .A2(n79), .ZN(\ab[8][10] ) );
  NOR2_X1 U184 ( .A1(n69), .A2(n79), .ZN(\ab[8][0] ) );
  NOR2_X1 U185 ( .A1(n138), .A2(n78), .ZN(\ab[7][9] ) );
  NOR2_X1 U186 ( .A1(n137), .A2(n78), .ZN(\ab[7][8] ) );
  NOR2_X1 U187 ( .A1(n136), .A2(n78), .ZN(\ab[7][7] ) );
  NOR2_X1 U188 ( .A1(n135), .A2(n78), .ZN(\ab[7][6] ) );
  NOR2_X1 U189 ( .A1(n134), .A2(n78), .ZN(\ab[7][5] ) );
  NOR2_X1 U190 ( .A1(n133), .A2(n78), .ZN(\ab[7][4] ) );
  NOR2_X1 U191 ( .A1(n132), .A2(n78), .ZN(\ab[7][3] ) );
  NOR2_X1 U192 ( .A1(n71), .A2(n78), .ZN(\ab[7][2] ) );
  NOR2_X1 U193 ( .A1(n123), .A2(n78), .ZN(\ab[7][24] ) );
  NOR2_X1 U194 ( .A1(n122), .A2(n78), .ZN(\ab[7][23] ) );
  NOR2_X1 U195 ( .A1(n121), .A2(n78), .ZN(\ab[7][22] ) );
  NOR2_X1 U196 ( .A1(n120), .A2(n78), .ZN(\ab[7][21] ) );
  NOR2_X1 U197 ( .A1(n119), .A2(n78), .ZN(\ab[7][20] ) );
  NOR2_X1 U198 ( .A1(n118), .A2(n78), .ZN(\ab[7][1] ) );
  NOR2_X1 U199 ( .A1(n117), .A2(n78), .ZN(\ab[7][19] ) );
  NOR2_X1 U200 ( .A1(n116), .A2(n78), .ZN(\ab[7][18] ) );
  NOR2_X1 U201 ( .A1(n115), .A2(n78), .ZN(\ab[7][17] ) );
  NOR2_X1 U202 ( .A1(n114), .A2(n78), .ZN(\ab[7][16] ) );
  NOR2_X1 U203 ( .A1(n113), .A2(n78), .ZN(\ab[7][15] ) );
  NOR2_X1 U204 ( .A1(n112), .A2(n78), .ZN(\ab[7][14] ) );
  NOR2_X1 U205 ( .A1(n111), .A2(n78), .ZN(\ab[7][13] ) );
  NOR2_X1 U206 ( .A1(n110), .A2(n78), .ZN(\ab[7][12] ) );
  NOR2_X1 U207 ( .A1(n109), .A2(n78), .ZN(\ab[7][11] ) );
  NOR2_X1 U208 ( .A1(n108), .A2(n78), .ZN(\ab[7][10] ) );
  NOR2_X1 U209 ( .A1(n69), .A2(n78), .ZN(\ab[7][0] ) );
  NOR2_X1 U210 ( .A1(n138), .A2(n77), .ZN(\ab[6][9] ) );
  NOR2_X1 U211 ( .A1(n137), .A2(n77), .ZN(\ab[6][8] ) );
  NOR2_X1 U212 ( .A1(n136), .A2(n77), .ZN(\ab[6][7] ) );
  NOR2_X1 U213 ( .A1(n135), .A2(n77), .ZN(\ab[6][6] ) );
  NOR2_X1 U214 ( .A1(n74), .A2(n77), .ZN(\ab[6][5] ) );
  NOR2_X1 U215 ( .A1(n133), .A2(n77), .ZN(\ab[6][4] ) );
  NOR2_X1 U216 ( .A1(n132), .A2(n77), .ZN(\ab[6][3] ) );
  NOR2_X1 U217 ( .A1(n71), .A2(n77), .ZN(\ab[6][2] ) );
  NOR2_X1 U218 ( .A1(n124), .A2(n77), .ZN(\ab[6][25] ) );
  NOR2_X1 U219 ( .A1(n123), .A2(n77), .ZN(\ab[6][24] ) );
  NOR2_X1 U220 ( .A1(n122), .A2(n77), .ZN(\ab[6][23] ) );
  NOR2_X1 U221 ( .A1(n121), .A2(n77), .ZN(\ab[6][22] ) );
  NOR2_X1 U222 ( .A1(n120), .A2(n77), .ZN(\ab[6][21] ) );
  NOR2_X1 U223 ( .A1(n119), .A2(n77), .ZN(\ab[6][20] ) );
  NOR2_X1 U224 ( .A1(n118), .A2(n77), .ZN(\ab[6][1] ) );
  NOR2_X1 U225 ( .A1(n117), .A2(n77), .ZN(\ab[6][19] ) );
  NOR2_X1 U226 ( .A1(n116), .A2(n77), .ZN(\ab[6][18] ) );
  NOR2_X1 U227 ( .A1(n115), .A2(n77), .ZN(\ab[6][17] ) );
  NOR2_X1 U228 ( .A1(n114), .A2(n77), .ZN(\ab[6][16] ) );
  NOR2_X1 U229 ( .A1(n113), .A2(n77), .ZN(\ab[6][15] ) );
  NOR2_X1 U230 ( .A1(n112), .A2(n77), .ZN(\ab[6][14] ) );
  NOR2_X1 U231 ( .A1(n111), .A2(n77), .ZN(\ab[6][13] ) );
  NOR2_X1 U232 ( .A1(n110), .A2(n77), .ZN(\ab[6][12] ) );
  NOR2_X1 U233 ( .A1(n109), .A2(n77), .ZN(\ab[6][11] ) );
  NOR2_X1 U234 ( .A1(n108), .A2(n77), .ZN(\ab[6][10] ) );
  NOR2_X1 U235 ( .A1(n69), .A2(n77), .ZN(\ab[6][0] ) );
  NOR2_X1 U236 ( .A1(n138), .A2(n75), .ZN(\ab[5][9] ) );
  NOR2_X1 U237 ( .A1(n137), .A2(n75), .ZN(\ab[5][8] ) );
  NOR2_X1 U238 ( .A1(n136), .A2(n75), .ZN(\ab[5][7] ) );
  NOR2_X1 U239 ( .A1(n135), .A2(n75), .ZN(\ab[5][6] ) );
  NOR2_X1 U240 ( .A1(n74), .A2(n75), .ZN(\ab[5][5] ) );
  NOR2_X1 U241 ( .A1(n133), .A2(n75), .ZN(\ab[5][4] ) );
  NOR2_X1 U242 ( .A1(n132), .A2(n75), .ZN(\ab[5][3] ) );
  NOR2_X1 U243 ( .A1(n71), .A2(n75), .ZN(\ab[5][2] ) );
  NOR2_X1 U244 ( .A1(n125), .A2(n75), .ZN(\ab[5][26] ) );
  NOR2_X1 U245 ( .A1(n124), .A2(n75), .ZN(\ab[5][25] ) );
  NOR2_X1 U246 ( .A1(n123), .A2(n75), .ZN(\ab[5][24] ) );
  NOR2_X1 U247 ( .A1(n122), .A2(n75), .ZN(\ab[5][23] ) );
  NOR2_X1 U248 ( .A1(n121), .A2(n75), .ZN(\ab[5][22] ) );
  NOR2_X1 U249 ( .A1(n120), .A2(n75), .ZN(\ab[5][21] ) );
  NOR2_X1 U250 ( .A1(n119), .A2(n75), .ZN(\ab[5][20] ) );
  NOR2_X1 U251 ( .A1(n118), .A2(n75), .ZN(\ab[5][1] ) );
  NOR2_X1 U252 ( .A1(n117), .A2(n75), .ZN(\ab[5][19] ) );
  NOR2_X1 U253 ( .A1(n116), .A2(n75), .ZN(\ab[5][18] ) );
  NOR2_X1 U254 ( .A1(n115), .A2(n75), .ZN(\ab[5][17] ) );
  NOR2_X1 U255 ( .A1(n114), .A2(n75), .ZN(\ab[5][16] ) );
  NOR2_X1 U256 ( .A1(n113), .A2(n75), .ZN(\ab[5][15] ) );
  NOR2_X1 U257 ( .A1(n112), .A2(n75), .ZN(\ab[5][14] ) );
  NOR2_X1 U258 ( .A1(n111), .A2(n75), .ZN(\ab[5][13] ) );
  NOR2_X1 U259 ( .A1(n110), .A2(n75), .ZN(\ab[5][12] ) );
  NOR2_X1 U260 ( .A1(n109), .A2(n75), .ZN(\ab[5][11] ) );
  NOR2_X1 U261 ( .A1(n108), .A2(n75), .ZN(\ab[5][10] ) );
  NOR2_X1 U262 ( .A1(n69), .A2(n75), .ZN(\ab[5][0] ) );
  NOR2_X1 U263 ( .A1(n138), .A2(n64), .ZN(\ab[4][9] ) );
  NOR2_X1 U264 ( .A1(n137), .A2(n64), .ZN(\ab[4][8] ) );
  NOR2_X1 U265 ( .A1(n136), .A2(n64), .ZN(\ab[4][7] ) );
  NOR2_X1 U266 ( .A1(n135), .A2(n64), .ZN(\ab[4][6] ) );
  NOR2_X1 U267 ( .A1(n74), .A2(n76), .ZN(\ab[4][5] ) );
  NOR2_X1 U268 ( .A1(n133), .A2(n76), .ZN(\ab[4][4] ) );
  NOR2_X1 U269 ( .A1(n132), .A2(n76), .ZN(\ab[4][3] ) );
  NOR2_X1 U270 ( .A1(n71), .A2(n76), .ZN(\ab[4][2] ) );
  NOR2_X1 U271 ( .A1(n126), .A2(n76), .ZN(\ab[4][27] ) );
  NOR2_X1 U272 ( .A1(n125), .A2(n76), .ZN(\ab[4][26] ) );
  NOR2_X1 U273 ( .A1(n124), .A2(n76), .ZN(\ab[4][25] ) );
  NOR2_X1 U274 ( .A1(n123), .A2(n76), .ZN(\ab[4][24] ) );
  NOR2_X1 U275 ( .A1(n122), .A2(n76), .ZN(\ab[4][23] ) );
  NOR2_X1 U276 ( .A1(n121), .A2(n76), .ZN(\ab[4][22] ) );
  NOR2_X1 U277 ( .A1(n120), .A2(n76), .ZN(\ab[4][21] ) );
  NOR2_X1 U278 ( .A1(n119), .A2(n76), .ZN(\ab[4][20] ) );
  NOR2_X1 U279 ( .A1(n118), .A2(n64), .ZN(\ab[4][1] ) );
  NOR2_X1 U280 ( .A1(n117), .A2(n64), .ZN(\ab[4][19] ) );
  NOR2_X1 U281 ( .A1(n116), .A2(n64), .ZN(\ab[4][18] ) );
  NOR2_X1 U282 ( .A1(n115), .A2(n64), .ZN(\ab[4][17] ) );
  NOR2_X1 U283 ( .A1(n114), .A2(n64), .ZN(\ab[4][16] ) );
  NOR2_X1 U284 ( .A1(n113), .A2(n64), .ZN(\ab[4][15] ) );
  NOR2_X1 U285 ( .A1(n112), .A2(n64), .ZN(\ab[4][14] ) );
  NOR2_X1 U286 ( .A1(n111), .A2(n64), .ZN(\ab[4][13] ) );
  NOR2_X1 U287 ( .A1(n110), .A2(n64), .ZN(\ab[4][12] ) );
  NOR2_X1 U288 ( .A1(n109), .A2(n64), .ZN(\ab[4][11] ) );
  NOR2_X1 U289 ( .A1(n108), .A2(n64), .ZN(\ab[4][10] ) );
  NOR2_X1 U290 ( .A1(n69), .A2(n64), .ZN(\ab[4][0] ) );
  NOR2_X1 U291 ( .A1(n138), .A2(n105), .ZN(\ab[3][9] ) );
  NOR2_X1 U292 ( .A1(n137), .A2(n105), .ZN(\ab[3][8] ) );
  NOR2_X1 U293 ( .A1(n136), .A2(n105), .ZN(\ab[3][7] ) );
  NOR2_X1 U294 ( .A1(n135), .A2(n105), .ZN(\ab[3][6] ) );
  NOR2_X1 U295 ( .A1(n74), .A2(n105), .ZN(\ab[3][5] ) );
  NOR2_X1 U296 ( .A1(n133), .A2(n67), .ZN(\ab[3][4] ) );
  NOR2_X1 U297 ( .A1(n132), .A2(n67), .ZN(\ab[3][3] ) );
  NOR2_X1 U298 ( .A1(n71), .A2(n67), .ZN(\ab[3][2] ) );
  NOR2_X1 U299 ( .A1(n127), .A2(n67), .ZN(\ab[3][28] ) );
  NOR2_X1 U300 ( .A1(n126), .A2(n67), .ZN(\ab[3][27] ) );
  NOR2_X1 U301 ( .A1(n125), .A2(n67), .ZN(\ab[3][26] ) );
  NOR2_X1 U302 ( .A1(n124), .A2(n67), .ZN(\ab[3][25] ) );
  NOR2_X1 U303 ( .A1(n123), .A2(n67), .ZN(\ab[3][24] ) );
  NOR2_X1 U304 ( .A1(n122), .A2(n67), .ZN(\ab[3][23] ) );
  NOR2_X1 U305 ( .A1(n121), .A2(n67), .ZN(\ab[3][22] ) );
  NOR2_X1 U306 ( .A1(n120), .A2(n67), .ZN(\ab[3][21] ) );
  NOR2_X1 U307 ( .A1(n119), .A2(n67), .ZN(\ab[3][20] ) );
  NOR2_X1 U308 ( .A1(n118), .A2(n105), .ZN(\ab[3][1] ) );
  NOR2_X1 U309 ( .A1(n117), .A2(n67), .ZN(\ab[3][19] ) );
  NOR2_X1 U310 ( .A1(n116), .A2(n105), .ZN(\ab[3][18] ) );
  NOR2_X1 U311 ( .A1(n115), .A2(n105), .ZN(\ab[3][17] ) );
  NOR2_X1 U312 ( .A1(n114), .A2(n105), .ZN(\ab[3][16] ) );
  NOR2_X1 U313 ( .A1(n113), .A2(n105), .ZN(\ab[3][15] ) );
  NOR2_X1 U314 ( .A1(n112), .A2(n105), .ZN(\ab[3][14] ) );
  NOR2_X1 U315 ( .A1(n111), .A2(n105), .ZN(\ab[3][13] ) );
  NOR2_X1 U316 ( .A1(n110), .A2(n105), .ZN(\ab[3][12] ) );
  NOR2_X1 U317 ( .A1(n109), .A2(n105), .ZN(\ab[3][11] ) );
  NOR2_X1 U318 ( .A1(n108), .A2(n105), .ZN(\ab[3][10] ) );
  NOR2_X1 U319 ( .A1(n69), .A2(n105), .ZN(\ab[3][0] ) );
  NOR2_X1 U320 ( .A1(n69), .A2(n99), .ZN(\ab[31][0] ) );
  NOR2_X1 U321 ( .A1(n70), .A2(n100), .ZN(\ab[30][1] ) );
  NOR2_X1 U322 ( .A1(n69), .A2(n100), .ZN(\ab[30][0] ) );
  NOR2_X1 U323 ( .A1(n138), .A2(n106), .ZN(\ab[2][9] ) );
  NOR2_X1 U324 ( .A1(n137), .A2(n106), .ZN(\ab[2][8] ) );
  NOR2_X1 U325 ( .A1(n136), .A2(n106), .ZN(\ab[2][7] ) );
  NOR2_X1 U326 ( .A1(n135), .A2(n106), .ZN(\ab[2][6] ) );
  NOR2_X1 U327 ( .A1(n74), .A2(n106), .ZN(\ab[2][5] ) );
  NOR2_X1 U328 ( .A1(n73), .A2(n106), .ZN(\ab[2][4] ) );
  NOR2_X1 U329 ( .A1(n72), .A2(n68), .ZN(\ab[2][3] ) );
  NOR2_X1 U330 ( .A1(n71), .A2(n68), .ZN(\ab[2][2] ) );
  NOR2_X1 U331 ( .A1(n128), .A2(n68), .ZN(\ab[2][29] ) );
  NOR2_X1 U332 ( .A1(n127), .A2(n68), .ZN(\ab[2][28] ) );
  NOR2_X1 U333 ( .A1(n126), .A2(n68), .ZN(\ab[2][27] ) );
  NOR2_X1 U334 ( .A1(n125), .A2(n68), .ZN(\ab[2][26] ) );
  NOR2_X1 U335 ( .A1(n124), .A2(n68), .ZN(\ab[2][25] ) );
  NOR2_X1 U336 ( .A1(n123), .A2(n68), .ZN(\ab[2][24] ) );
  NOR2_X1 U337 ( .A1(n122), .A2(n68), .ZN(\ab[2][23] ) );
  NOR2_X1 U338 ( .A1(n121), .A2(n68), .ZN(\ab[2][22] ) );
  NOR2_X1 U339 ( .A1(n120), .A2(n68), .ZN(\ab[2][21] ) );
  NOR2_X1 U340 ( .A1(n119), .A2(n68), .ZN(\ab[2][20] ) );
  NOR2_X1 U341 ( .A1(n70), .A2(n106), .ZN(\ab[2][1] ) );
  NOR2_X1 U342 ( .A1(n117), .A2(n68), .ZN(\ab[2][19] ) );
  NOR2_X1 U343 ( .A1(n116), .A2(n106), .ZN(\ab[2][18] ) );
  NOR2_X1 U344 ( .A1(n115), .A2(n106), .ZN(\ab[2][17] ) );
  NOR2_X1 U345 ( .A1(n114), .A2(n106), .ZN(\ab[2][16] ) );
  NOR2_X1 U346 ( .A1(n113), .A2(n106), .ZN(\ab[2][15] ) );
  NOR2_X1 U347 ( .A1(n112), .A2(n106), .ZN(\ab[2][14] ) );
  NOR2_X1 U348 ( .A1(n111), .A2(n106), .ZN(\ab[2][13] ) );
  NOR2_X1 U349 ( .A1(n110), .A2(n106), .ZN(\ab[2][12] ) );
  NOR2_X1 U350 ( .A1(n109), .A2(n106), .ZN(\ab[2][11] ) );
  NOR2_X1 U351 ( .A1(n108), .A2(n106), .ZN(\ab[2][10] ) );
  NOR2_X1 U352 ( .A1(n69), .A2(n106), .ZN(\ab[2][0] ) );
  NOR2_X1 U353 ( .A1(n71), .A2(n101), .ZN(\ab[29][2] ) );
  NOR2_X1 U354 ( .A1(n70), .A2(n101), .ZN(\ab[29][1] ) );
  NOR2_X1 U355 ( .A1(n69), .A2(n101), .ZN(\ab[29][0] ) );
  NOR2_X1 U356 ( .A1(n132), .A2(n102), .ZN(\ab[28][3] ) );
  NOR2_X1 U357 ( .A1(n71), .A2(n102), .ZN(\ab[28][2] ) );
  NOR2_X1 U358 ( .A1(n70), .A2(n102), .ZN(\ab[28][1] ) );
  NOR2_X1 U359 ( .A1(n69), .A2(n102), .ZN(\ab[28][0] ) );
  NOR2_X1 U360 ( .A1(n133), .A2(n94), .ZN(\ab[27][4] ) );
  NOR2_X1 U361 ( .A1(n132), .A2(n94), .ZN(\ab[27][3] ) );
  NOR2_X1 U362 ( .A1(n71), .A2(n94), .ZN(\ab[27][2] ) );
  NOR2_X1 U363 ( .A1(n70), .A2(n94), .ZN(\ab[27][1] ) );
  NOR2_X1 U364 ( .A1(n69), .A2(n94), .ZN(\ab[27][0] ) );
  NOR2_X1 U365 ( .A1(n74), .A2(n93), .ZN(\ab[26][5] ) );
  NOR2_X1 U366 ( .A1(n133), .A2(n93), .ZN(\ab[26][4] ) );
  NOR2_X1 U367 ( .A1(n132), .A2(n93), .ZN(\ab[26][3] ) );
  NOR2_X1 U368 ( .A1(n71), .A2(n93), .ZN(\ab[26][2] ) );
  NOR2_X1 U369 ( .A1(n70), .A2(n93), .ZN(\ab[26][1] ) );
  NOR2_X1 U370 ( .A1(n69), .A2(n93), .ZN(\ab[26][0] ) );
  NOR2_X1 U371 ( .A1(n135), .A2(n92), .ZN(\ab[25][6] ) );
  NOR2_X1 U372 ( .A1(n74), .A2(n92), .ZN(\ab[25][5] ) );
  NOR2_X1 U373 ( .A1(n133), .A2(n92), .ZN(\ab[25][4] ) );
  NOR2_X1 U374 ( .A1(n132), .A2(n92), .ZN(\ab[25][3] ) );
  NOR2_X1 U375 ( .A1(n71), .A2(n92), .ZN(\ab[25][2] ) );
  NOR2_X1 U376 ( .A1(n70), .A2(n92), .ZN(\ab[25][1] ) );
  NOR2_X1 U377 ( .A1(n69), .A2(n92), .ZN(\ab[25][0] ) );
  NOR2_X1 U378 ( .A1(n136), .A2(n91), .ZN(\ab[24][7] ) );
  NOR2_X1 U379 ( .A1(n135), .A2(n91), .ZN(\ab[24][6] ) );
  NOR2_X1 U380 ( .A1(n74), .A2(n91), .ZN(\ab[24][5] ) );
  NOR2_X1 U381 ( .A1(n133), .A2(n91), .ZN(\ab[24][4] ) );
  NOR2_X1 U382 ( .A1(n132), .A2(n91), .ZN(\ab[24][3] ) );
  NOR2_X1 U383 ( .A1(n71), .A2(n91), .ZN(\ab[24][2] ) );
  NOR2_X1 U384 ( .A1(n70), .A2(n91), .ZN(\ab[24][1] ) );
  NOR2_X1 U385 ( .A1(n69), .A2(n91), .ZN(\ab[24][0] ) );
  NOR2_X1 U386 ( .A1(n137), .A2(n98), .ZN(\ab[23][8] ) );
  NOR2_X1 U387 ( .A1(n136), .A2(n98), .ZN(\ab[23][7] ) );
  NOR2_X1 U388 ( .A1(n135), .A2(n98), .ZN(\ab[23][6] ) );
  NOR2_X1 U389 ( .A1(n74), .A2(n98), .ZN(\ab[23][5] ) );
  NOR2_X1 U390 ( .A1(n133), .A2(n98), .ZN(\ab[23][4] ) );
  NOR2_X1 U391 ( .A1(n132), .A2(n98), .ZN(\ab[23][3] ) );
  NOR2_X1 U392 ( .A1(n71), .A2(n98), .ZN(\ab[23][2] ) );
  NOR2_X1 U393 ( .A1(n70), .A2(n98), .ZN(\ab[23][1] ) );
  NOR2_X1 U394 ( .A1(n69), .A2(n98), .ZN(\ab[23][0] ) );
  NOR2_X1 U395 ( .A1(n138), .A2(n95), .ZN(\ab[22][9] ) );
  NOR2_X1 U396 ( .A1(n137), .A2(n95), .ZN(\ab[22][8] ) );
  NOR2_X1 U397 ( .A1(n136), .A2(n95), .ZN(\ab[22][7] ) );
  NOR2_X1 U398 ( .A1(n135), .A2(n95), .ZN(\ab[22][6] ) );
  NOR2_X1 U399 ( .A1(n74), .A2(n95), .ZN(\ab[22][5] ) );
  NOR2_X1 U400 ( .A1(n133), .A2(n95), .ZN(\ab[22][4] ) );
  NOR2_X1 U401 ( .A1(n132), .A2(n95), .ZN(\ab[22][3] ) );
  NOR2_X1 U402 ( .A1(n71), .A2(n95), .ZN(\ab[22][2] ) );
  NOR2_X1 U403 ( .A1(n70), .A2(n95), .ZN(\ab[22][1] ) );
  NOR2_X1 U404 ( .A1(n69), .A2(n95), .ZN(\ab[22][0] ) );
  NOR2_X1 U405 ( .A1(n138), .A2(n96), .ZN(\ab[21][9] ) );
  NOR2_X1 U406 ( .A1(n137), .A2(n96), .ZN(\ab[21][8] ) );
  NOR2_X1 U407 ( .A1(n136), .A2(n96), .ZN(\ab[21][7] ) );
  NOR2_X1 U408 ( .A1(n135), .A2(n96), .ZN(\ab[21][6] ) );
  NOR2_X1 U409 ( .A1(n74), .A2(n96), .ZN(\ab[21][5] ) );
  NOR2_X1 U410 ( .A1(n133), .A2(n96), .ZN(\ab[21][4] ) );
  NOR2_X1 U411 ( .A1(n132), .A2(n96), .ZN(\ab[21][3] ) );
  NOR2_X1 U412 ( .A1(n71), .A2(n96), .ZN(\ab[21][2] ) );
  NOR2_X1 U413 ( .A1(n70), .A2(n96), .ZN(\ab[21][1] ) );
  NOR2_X1 U414 ( .A1(n108), .A2(n96), .ZN(\ab[21][10] ) );
  NOR2_X1 U415 ( .A1(n69), .A2(n96), .ZN(\ab[21][0] ) );
  NOR2_X1 U416 ( .A1(n138), .A2(n97), .ZN(\ab[20][9] ) );
  NOR2_X1 U417 ( .A1(n137), .A2(n97), .ZN(\ab[20][8] ) );
  NOR2_X1 U418 ( .A1(n136), .A2(n97), .ZN(\ab[20][7] ) );
  NOR2_X1 U419 ( .A1(n135), .A2(n97), .ZN(\ab[20][6] ) );
  NOR2_X1 U420 ( .A1(n74), .A2(n97), .ZN(\ab[20][5] ) );
  NOR2_X1 U421 ( .A1(n133), .A2(n97), .ZN(\ab[20][4] ) );
  NOR2_X1 U422 ( .A1(n132), .A2(n97), .ZN(\ab[20][3] ) );
  NOR2_X1 U423 ( .A1(n71), .A2(n97), .ZN(\ab[20][2] ) );
  NOR2_X1 U424 ( .A1(n70), .A2(n97), .ZN(\ab[20][1] ) );
  NOR2_X1 U425 ( .A1(n109), .A2(n97), .ZN(\ab[20][11] ) );
  NOR2_X1 U426 ( .A1(n108), .A2(n97), .ZN(\ab[20][10] ) );
  NOR2_X1 U427 ( .A1(n69), .A2(n97), .ZN(\ab[20][0] ) );
  NOR2_X1 U428 ( .A1(n138), .A2(n65), .ZN(\ab[1][9] ) );
  NOR2_X1 U429 ( .A1(n137), .A2(n65), .ZN(\ab[1][8] ) );
  NOR2_X1 U430 ( .A1(n136), .A2(n65), .ZN(\ab[1][7] ) );
  NOR2_X1 U431 ( .A1(n135), .A2(n65), .ZN(\ab[1][6] ) );
  NOR2_X1 U432 ( .A1(n134), .A2(n65), .ZN(\ab[1][5] ) );
  NOR2_X1 U433 ( .A1(n73), .A2(n65), .ZN(\ab[1][4] ) );
  NOR2_X1 U434 ( .A1(n72), .A2(n65), .ZN(\ab[1][3] ) );
  NOR2_X1 U435 ( .A1(n130), .A2(n103), .ZN(\ab[1][30] ) );
  NOR2_X1 U436 ( .A1(n129), .A2(n65), .ZN(\ab[1][2] ) );
  NOR2_X1 U437 ( .A1(n128), .A2(n103), .ZN(\ab[1][29] ) );
  NOR2_X1 U438 ( .A1(n127), .A2(n103), .ZN(\ab[1][28] ) );
  NOR2_X1 U439 ( .A1(n126), .A2(n103), .ZN(\ab[1][27] ) );
  NOR2_X1 U440 ( .A1(n125), .A2(n103), .ZN(\ab[1][26] ) );
  NOR2_X1 U441 ( .A1(n124), .A2(n103), .ZN(\ab[1][25] ) );
  NOR2_X1 U442 ( .A1(n123), .A2(n103), .ZN(\ab[1][24] ) );
  NOR2_X1 U443 ( .A1(n122), .A2(n103), .ZN(\ab[1][23] ) );
  NOR2_X1 U444 ( .A1(n121), .A2(n103), .ZN(\ab[1][22] ) );
  NOR2_X1 U445 ( .A1(n120), .A2(n103), .ZN(\ab[1][21] ) );
  NOR2_X1 U446 ( .A1(n119), .A2(n65), .ZN(\ab[1][20] ) );
  NOR2_X1 U447 ( .A1(n118), .A2(n65), .ZN(\ab[1][1] ) );
  NOR2_X1 U448 ( .A1(n117), .A2(n65), .ZN(\ab[1][19] ) );
  NOR2_X1 U449 ( .A1(n116), .A2(n65), .ZN(\ab[1][18] ) );
  NOR2_X1 U450 ( .A1(n115), .A2(n65), .ZN(\ab[1][17] ) );
  NOR2_X1 U451 ( .A1(n114), .A2(n65), .ZN(\ab[1][16] ) );
  NOR2_X1 U452 ( .A1(n113), .A2(n65), .ZN(\ab[1][15] ) );
  NOR2_X1 U453 ( .A1(n112), .A2(n65), .ZN(\ab[1][14] ) );
  NOR2_X1 U454 ( .A1(n111), .A2(n65), .ZN(\ab[1][13] ) );
  NOR2_X1 U455 ( .A1(n110), .A2(n65), .ZN(\ab[1][12] ) );
  NOR2_X1 U456 ( .A1(n109), .A2(n65), .ZN(\ab[1][11] ) );
  NOR2_X1 U457 ( .A1(n108), .A2(n65), .ZN(\ab[1][10] ) );
  NOR2_X1 U458 ( .A1(n107), .A2(n65), .ZN(\ab[1][0] ) );
  NOR2_X1 U459 ( .A1(n138), .A2(n86), .ZN(\ab[19][9] ) );
  NOR2_X1 U460 ( .A1(n137), .A2(n86), .ZN(\ab[19][8] ) );
  NOR2_X1 U461 ( .A1(n136), .A2(n86), .ZN(\ab[19][7] ) );
  NOR2_X1 U462 ( .A1(n135), .A2(n86), .ZN(\ab[19][6] ) );
  NOR2_X1 U463 ( .A1(n134), .A2(n86), .ZN(\ab[19][5] ) );
  NOR2_X1 U464 ( .A1(n73), .A2(n86), .ZN(\ab[19][4] ) );
  NOR2_X1 U465 ( .A1(n72), .A2(n86), .ZN(\ab[19][3] ) );
  NOR2_X1 U466 ( .A1(n129), .A2(n86), .ZN(\ab[19][2] ) );
  NOR2_X1 U467 ( .A1(n118), .A2(n86), .ZN(\ab[19][1] ) );
  NOR2_X1 U468 ( .A1(n110), .A2(n86), .ZN(\ab[19][12] ) );
  NOR2_X1 U469 ( .A1(n109), .A2(n86), .ZN(\ab[19][11] ) );
  NOR2_X1 U470 ( .A1(n108), .A2(n86), .ZN(\ab[19][10] ) );
  NOR2_X1 U471 ( .A1(n107), .A2(n86), .ZN(\ab[19][0] ) );
  NOR2_X1 U472 ( .A1(n138), .A2(n83), .ZN(\ab[18][9] ) );
  NOR2_X1 U473 ( .A1(n137), .A2(n83), .ZN(\ab[18][8] ) );
  NOR2_X1 U474 ( .A1(n136), .A2(n83), .ZN(\ab[18][7] ) );
  NOR2_X1 U475 ( .A1(n135), .A2(n83), .ZN(\ab[18][6] ) );
  NOR2_X1 U476 ( .A1(n134), .A2(n83), .ZN(\ab[18][5] ) );
  NOR2_X1 U477 ( .A1(n73), .A2(n83), .ZN(\ab[18][4] ) );
  NOR2_X1 U478 ( .A1(n72), .A2(n83), .ZN(\ab[18][3] ) );
  NOR2_X1 U479 ( .A1(n129), .A2(n83), .ZN(\ab[18][2] ) );
  NOR2_X1 U480 ( .A1(n118), .A2(n83), .ZN(\ab[18][1] ) );
  NOR2_X1 U481 ( .A1(n111), .A2(n83), .ZN(\ab[18][13] ) );
  NOR2_X1 U482 ( .A1(n110), .A2(n83), .ZN(\ab[18][12] ) );
  NOR2_X1 U483 ( .A1(n109), .A2(n83), .ZN(\ab[18][11] ) );
  NOR2_X1 U484 ( .A1(n108), .A2(n83), .ZN(\ab[18][10] ) );
  NOR2_X1 U485 ( .A1(n107), .A2(n83), .ZN(\ab[18][0] ) );
  NOR2_X1 U486 ( .A1(n138), .A2(n84), .ZN(\ab[17][9] ) );
  NOR2_X1 U487 ( .A1(n137), .A2(n84), .ZN(\ab[17][8] ) );
  NOR2_X1 U488 ( .A1(n136), .A2(n84), .ZN(\ab[17][7] ) );
  NOR2_X1 U489 ( .A1(n135), .A2(n84), .ZN(\ab[17][6] ) );
  NOR2_X1 U490 ( .A1(n134), .A2(n84), .ZN(\ab[17][5] ) );
  NOR2_X1 U491 ( .A1(n73), .A2(n84), .ZN(\ab[17][4] ) );
  NOR2_X1 U492 ( .A1(n72), .A2(n84), .ZN(\ab[17][3] ) );
  NOR2_X1 U493 ( .A1(n129), .A2(n84), .ZN(\ab[17][2] ) );
  NOR2_X1 U494 ( .A1(n118), .A2(n84), .ZN(\ab[17][1] ) );
  NOR2_X1 U495 ( .A1(n112), .A2(n84), .ZN(\ab[17][14] ) );
  NOR2_X1 U496 ( .A1(n111), .A2(n84), .ZN(\ab[17][13] ) );
  NOR2_X1 U497 ( .A1(n110), .A2(n84), .ZN(\ab[17][12] ) );
  NOR2_X1 U498 ( .A1(n109), .A2(n84), .ZN(\ab[17][11] ) );
  NOR2_X1 U499 ( .A1(n108), .A2(n84), .ZN(\ab[17][10] ) );
  NOR2_X1 U500 ( .A1(n107), .A2(n84), .ZN(\ab[17][0] ) );
  NOR2_X1 U501 ( .A1(n138), .A2(n85), .ZN(\ab[16][9] ) );
  NOR2_X1 U502 ( .A1(n137), .A2(n85), .ZN(\ab[16][8] ) );
  NOR2_X1 U503 ( .A1(n136), .A2(n85), .ZN(\ab[16][7] ) );
  NOR2_X1 U504 ( .A1(n135), .A2(n85), .ZN(\ab[16][6] ) );
  NOR2_X1 U505 ( .A1(n134), .A2(n85), .ZN(\ab[16][5] ) );
  NOR2_X1 U506 ( .A1(n73), .A2(n85), .ZN(\ab[16][4] ) );
  NOR2_X1 U507 ( .A1(n72), .A2(n85), .ZN(\ab[16][3] ) );
  NOR2_X1 U508 ( .A1(n129), .A2(n85), .ZN(\ab[16][2] ) );
  NOR2_X1 U509 ( .A1(n118), .A2(n85), .ZN(\ab[16][1] ) );
  NOR2_X1 U510 ( .A1(n113), .A2(n85), .ZN(\ab[16][15] ) );
  NOR2_X1 U511 ( .A1(n112), .A2(n85), .ZN(\ab[16][14] ) );
  NOR2_X1 U512 ( .A1(n111), .A2(n85), .ZN(\ab[16][13] ) );
  NOR2_X1 U513 ( .A1(n110), .A2(n85), .ZN(\ab[16][12] ) );
  NOR2_X1 U514 ( .A1(n109), .A2(n85), .ZN(\ab[16][11] ) );
  NOR2_X1 U515 ( .A1(n108), .A2(n85), .ZN(\ab[16][10] ) );
  NOR2_X1 U516 ( .A1(n107), .A2(n85), .ZN(\ab[16][0] ) );
  NOR2_X1 U517 ( .A1(n138), .A2(n90), .ZN(\ab[15][9] ) );
  NOR2_X1 U518 ( .A1(n137), .A2(n90), .ZN(\ab[15][8] ) );
  NOR2_X1 U519 ( .A1(n136), .A2(n90), .ZN(\ab[15][7] ) );
  NOR2_X1 U520 ( .A1(n135), .A2(n90), .ZN(\ab[15][6] ) );
  NOR2_X1 U521 ( .A1(n134), .A2(n90), .ZN(\ab[15][5] ) );
  NOR2_X1 U522 ( .A1(n73), .A2(n90), .ZN(\ab[15][4] ) );
  NOR2_X1 U523 ( .A1(n72), .A2(n90), .ZN(\ab[15][3] ) );
  NOR2_X1 U524 ( .A1(n129), .A2(n90), .ZN(\ab[15][2] ) );
  NOR2_X1 U525 ( .A1(n118), .A2(n90), .ZN(\ab[15][1] ) );
  NOR2_X1 U526 ( .A1(n114), .A2(n90), .ZN(\ab[15][16] ) );
  NOR2_X1 U527 ( .A1(n113), .A2(n90), .ZN(\ab[15][15] ) );
  NOR2_X1 U528 ( .A1(n112), .A2(n90), .ZN(\ab[15][14] ) );
  NOR2_X1 U529 ( .A1(n111), .A2(n90), .ZN(\ab[15][13] ) );
  NOR2_X1 U530 ( .A1(n110), .A2(n90), .ZN(\ab[15][12] ) );
  NOR2_X1 U531 ( .A1(n109), .A2(n90), .ZN(\ab[15][11] ) );
  NOR2_X1 U532 ( .A1(n108), .A2(n90), .ZN(\ab[15][10] ) );
  NOR2_X1 U533 ( .A1(n107), .A2(n90), .ZN(\ab[15][0] ) );
  NOR2_X1 U534 ( .A1(n138), .A2(n87), .ZN(\ab[14][9] ) );
  NOR2_X1 U535 ( .A1(n137), .A2(n87), .ZN(\ab[14][8] ) );
  NOR2_X1 U536 ( .A1(n136), .A2(n87), .ZN(\ab[14][7] ) );
  NOR2_X1 U537 ( .A1(n135), .A2(n87), .ZN(\ab[14][6] ) );
  NOR2_X1 U538 ( .A1(n134), .A2(n87), .ZN(\ab[14][5] ) );
  NOR2_X1 U539 ( .A1(n73), .A2(n87), .ZN(\ab[14][4] ) );
  NOR2_X1 U540 ( .A1(n72), .A2(n87), .ZN(\ab[14][3] ) );
  NOR2_X1 U541 ( .A1(n129), .A2(n87), .ZN(\ab[14][2] ) );
  NOR2_X1 U542 ( .A1(n118), .A2(n87), .ZN(\ab[14][1] ) );
  NOR2_X1 U543 ( .A1(n115), .A2(n87), .ZN(\ab[14][17] ) );
  NOR2_X1 U544 ( .A1(n114), .A2(n87), .ZN(\ab[14][16] ) );
  NOR2_X1 U545 ( .A1(n113), .A2(n87), .ZN(\ab[14][15] ) );
  NOR2_X1 U546 ( .A1(n112), .A2(n87), .ZN(\ab[14][14] ) );
  NOR2_X1 U547 ( .A1(n111), .A2(n87), .ZN(\ab[14][13] ) );
  NOR2_X1 U548 ( .A1(n110), .A2(n87), .ZN(\ab[14][12] ) );
  NOR2_X1 U549 ( .A1(n109), .A2(n87), .ZN(\ab[14][11] ) );
  NOR2_X1 U550 ( .A1(n108), .A2(n87), .ZN(\ab[14][10] ) );
  NOR2_X1 U551 ( .A1(n107), .A2(n87), .ZN(\ab[14][0] ) );
  NOR2_X1 U552 ( .A1(n138), .A2(n88), .ZN(\ab[13][9] ) );
  NOR2_X1 U553 ( .A1(n137), .A2(n88), .ZN(\ab[13][8] ) );
  NOR2_X1 U554 ( .A1(n136), .A2(n88), .ZN(\ab[13][7] ) );
  NOR2_X1 U555 ( .A1(n135), .A2(n88), .ZN(\ab[13][6] ) );
  NOR2_X1 U556 ( .A1(n134), .A2(n88), .ZN(\ab[13][5] ) );
  NOR2_X1 U557 ( .A1(n73), .A2(n88), .ZN(\ab[13][4] ) );
  NOR2_X1 U558 ( .A1(n72), .A2(n88), .ZN(\ab[13][3] ) );
  NOR2_X1 U559 ( .A1(n129), .A2(n88), .ZN(\ab[13][2] ) );
  NOR2_X1 U560 ( .A1(n118), .A2(n88), .ZN(\ab[13][1] ) );
  NOR2_X1 U561 ( .A1(n116), .A2(n88), .ZN(\ab[13][18] ) );
  NOR2_X1 U562 ( .A1(n115), .A2(n88), .ZN(\ab[13][17] ) );
  NOR2_X1 U563 ( .A1(n114), .A2(n88), .ZN(\ab[13][16] ) );
  NOR2_X1 U564 ( .A1(n113), .A2(n88), .ZN(\ab[13][15] ) );
  NOR2_X1 U565 ( .A1(n112), .A2(n88), .ZN(\ab[13][14] ) );
  NOR2_X1 U566 ( .A1(n111), .A2(n88), .ZN(\ab[13][13] ) );
  NOR2_X1 U567 ( .A1(n110), .A2(n88), .ZN(\ab[13][12] ) );
  NOR2_X1 U568 ( .A1(n109), .A2(n88), .ZN(\ab[13][11] ) );
  NOR2_X1 U569 ( .A1(n108), .A2(n88), .ZN(\ab[13][10] ) );
  NOR2_X1 U570 ( .A1(n107), .A2(n88), .ZN(\ab[13][0] ) );
  NOR2_X1 U571 ( .A1(n138), .A2(n89), .ZN(\ab[12][9] ) );
  NOR2_X1 U572 ( .A1(n137), .A2(n89), .ZN(\ab[12][8] ) );
  NOR2_X1 U573 ( .A1(n136), .A2(n89), .ZN(\ab[12][7] ) );
  NOR2_X1 U574 ( .A1(n135), .A2(n89), .ZN(\ab[12][6] ) );
  NOR2_X1 U575 ( .A1(n134), .A2(n89), .ZN(\ab[12][5] ) );
  NOR2_X1 U576 ( .A1(n73), .A2(n89), .ZN(\ab[12][4] ) );
  NOR2_X1 U577 ( .A1(n72), .A2(n89), .ZN(\ab[12][3] ) );
  NOR2_X1 U578 ( .A1(n129), .A2(n89), .ZN(\ab[12][2] ) );
  NOR2_X1 U579 ( .A1(n118), .A2(n89), .ZN(\ab[12][1] ) );
  NOR2_X1 U580 ( .A1(n117), .A2(n89), .ZN(\ab[12][19] ) );
  NOR2_X1 U581 ( .A1(n116), .A2(n89), .ZN(\ab[12][18] ) );
  NOR2_X1 U582 ( .A1(n115), .A2(n89), .ZN(\ab[12][17] ) );
  NOR2_X1 U583 ( .A1(n114), .A2(n89), .ZN(\ab[12][16] ) );
  NOR2_X1 U584 ( .A1(n113), .A2(n89), .ZN(\ab[12][15] ) );
  NOR2_X1 U585 ( .A1(n112), .A2(n89), .ZN(\ab[12][14] ) );
  NOR2_X1 U586 ( .A1(n111), .A2(n89), .ZN(\ab[12][13] ) );
  NOR2_X1 U587 ( .A1(n110), .A2(n89), .ZN(\ab[12][12] ) );
  NOR2_X1 U588 ( .A1(n109), .A2(n89), .ZN(\ab[12][11] ) );
  NOR2_X1 U589 ( .A1(n108), .A2(n89), .ZN(\ab[12][10] ) );
  NOR2_X1 U590 ( .A1(n107), .A2(n89), .ZN(\ab[12][0] ) );
  NOR2_X1 U591 ( .A1(n138), .A2(n82), .ZN(\ab[11][9] ) );
  NOR2_X1 U592 ( .A1(n137), .A2(n82), .ZN(\ab[11][8] ) );
  NOR2_X1 U593 ( .A1(n136), .A2(n82), .ZN(\ab[11][7] ) );
  NOR2_X1 U594 ( .A1(n135), .A2(n82), .ZN(\ab[11][6] ) );
  NOR2_X1 U595 ( .A1(n134), .A2(n82), .ZN(\ab[11][5] ) );
  NOR2_X1 U596 ( .A1(n73), .A2(n82), .ZN(\ab[11][4] ) );
  NOR2_X1 U597 ( .A1(n72), .A2(n82), .ZN(\ab[11][3] ) );
  NOR2_X1 U598 ( .A1(n129), .A2(n82), .ZN(\ab[11][2] ) );
  NOR2_X1 U599 ( .A1(n119), .A2(n82), .ZN(\ab[11][20] ) );
  NOR2_X1 U600 ( .A1(n118), .A2(n82), .ZN(\ab[11][1] ) );
  NOR2_X1 U601 ( .A1(n117), .A2(n82), .ZN(\ab[11][19] ) );
  NOR2_X1 U602 ( .A1(n116), .A2(n82), .ZN(\ab[11][18] ) );
  NOR2_X1 U603 ( .A1(n115), .A2(n82), .ZN(\ab[11][17] ) );
  NOR2_X1 U604 ( .A1(n114), .A2(n82), .ZN(\ab[11][16] ) );
  NOR2_X1 U605 ( .A1(n113), .A2(n82), .ZN(\ab[11][15] ) );
  NOR2_X1 U606 ( .A1(n112), .A2(n82), .ZN(\ab[11][14] ) );
  NOR2_X1 U607 ( .A1(n111), .A2(n82), .ZN(\ab[11][13] ) );
  NOR2_X1 U608 ( .A1(n110), .A2(n82), .ZN(\ab[11][12] ) );
  NOR2_X1 U609 ( .A1(n109), .A2(n82), .ZN(\ab[11][11] ) );
  NOR2_X1 U610 ( .A1(n108), .A2(n82), .ZN(\ab[11][10] ) );
  NOR2_X1 U611 ( .A1(n107), .A2(n82), .ZN(\ab[11][0] ) );
  NOR2_X1 U612 ( .A1(n138), .A2(n81), .ZN(\ab[10][9] ) );
  NOR2_X1 U613 ( .A1(n137), .A2(n81), .ZN(\ab[10][8] ) );
  NOR2_X1 U614 ( .A1(n136), .A2(n81), .ZN(\ab[10][7] ) );
  NOR2_X1 U615 ( .A1(n135), .A2(n81), .ZN(\ab[10][6] ) );
  NOR2_X1 U616 ( .A1(n134), .A2(n81), .ZN(\ab[10][5] ) );
  NOR2_X1 U617 ( .A1(n73), .A2(n81), .ZN(\ab[10][4] ) );
  NOR2_X1 U618 ( .A1(n72), .A2(n81), .ZN(\ab[10][3] ) );
  NOR2_X1 U619 ( .A1(n129), .A2(n81), .ZN(\ab[10][2] ) );
  NOR2_X1 U620 ( .A1(n120), .A2(n81), .ZN(\ab[10][21] ) );
  NOR2_X1 U621 ( .A1(n119), .A2(n81), .ZN(\ab[10][20] ) );
  NOR2_X1 U622 ( .A1(n118), .A2(n81), .ZN(\ab[10][1] ) );
  NOR2_X1 U623 ( .A1(n117), .A2(n81), .ZN(\ab[10][19] ) );
  NOR2_X1 U624 ( .A1(n116), .A2(n81), .ZN(\ab[10][18] ) );
  NOR2_X1 U625 ( .A1(n115), .A2(n81), .ZN(\ab[10][17] ) );
  NOR2_X1 U626 ( .A1(n114), .A2(n81), .ZN(\ab[10][16] ) );
  NOR2_X1 U627 ( .A1(n113), .A2(n81), .ZN(\ab[10][15] ) );
  NOR2_X1 U628 ( .A1(n112), .A2(n81), .ZN(\ab[10][14] ) );
  NOR2_X1 U629 ( .A1(n111), .A2(n81), .ZN(\ab[10][13] ) );
  NOR2_X1 U630 ( .A1(n110), .A2(n81), .ZN(\ab[10][12] ) );
  NOR2_X1 U631 ( .A1(n109), .A2(n81), .ZN(\ab[10][11] ) );
  NOR2_X1 U632 ( .A1(n108), .A2(n81), .ZN(\ab[10][10] ) );
  NOR2_X1 U633 ( .A1(n107), .A2(n81), .ZN(\ab[10][0] ) );
  NOR2_X1 U634 ( .A1(n138), .A2(n104), .ZN(\ab[0][9] ) );
  NOR2_X1 U635 ( .A1(n137), .A2(n104), .ZN(\ab[0][8] ) );
  NOR2_X1 U636 ( .A1(n136), .A2(n104), .ZN(\ab[0][7] ) );
  NOR2_X1 U637 ( .A1(n135), .A2(n104), .ZN(\ab[0][6] ) );
  NOR2_X1 U638 ( .A1(n134), .A2(n104), .ZN(\ab[0][5] ) );
  NOR2_X1 U639 ( .A1(n73), .A2(n104), .ZN(\ab[0][4] ) );
  NOR2_X1 U640 ( .A1(n72), .A2(n104), .ZN(\ab[0][3] ) );
  NOR2_X1 U641 ( .A1(n131), .A2(n104), .ZN(\ab[0][31] ) );
  NOR2_X1 U642 ( .A1(n130), .A2(n66), .ZN(\ab[0][30] ) );
  NOR2_X1 U643 ( .A1(n129), .A2(n66), .ZN(\ab[0][2] ) );
  NOR2_X1 U644 ( .A1(n128), .A2(n66), .ZN(\ab[0][29] ) );
  NOR2_X1 U645 ( .A1(n127), .A2(n66), .ZN(\ab[0][28] ) );
  NOR2_X1 U646 ( .A1(n126), .A2(n66), .ZN(\ab[0][27] ) );
  NOR2_X1 U647 ( .A1(n125), .A2(n66), .ZN(\ab[0][26] ) );
  NOR2_X1 U648 ( .A1(n124), .A2(n66), .ZN(\ab[0][25] ) );
  NOR2_X1 U649 ( .A1(n123), .A2(n66), .ZN(\ab[0][24] ) );
  NOR2_X1 U650 ( .A1(n122), .A2(n66), .ZN(\ab[0][23] ) );
  NOR2_X1 U651 ( .A1(n121), .A2(n66), .ZN(\ab[0][22] ) );
  NOR2_X1 U652 ( .A1(n120), .A2(n66), .ZN(\ab[0][21] ) );
  NOR2_X1 U653 ( .A1(n119), .A2(n66), .ZN(\ab[0][20] ) );
  NOR2_X1 U654 ( .A1(n118), .A2(n104), .ZN(\ab[0][1] ) );
  NOR2_X1 U655 ( .A1(n117), .A2(n104), .ZN(\ab[0][19] ) );
  NOR2_X1 U656 ( .A1(n116), .A2(n104), .ZN(\ab[0][18] ) );
  NOR2_X1 U657 ( .A1(n115), .A2(n104), .ZN(\ab[0][17] ) );
  NOR2_X1 U658 ( .A1(n114), .A2(n104), .ZN(\ab[0][16] ) );
  NOR2_X1 U659 ( .A1(n113), .A2(n104), .ZN(\ab[0][15] ) );
  NOR2_X1 U660 ( .A1(n112), .A2(n104), .ZN(\ab[0][14] ) );
  NOR2_X1 U661 ( .A1(n111), .A2(n104), .ZN(\ab[0][13] ) );
  NOR2_X1 U662 ( .A1(n110), .A2(n104), .ZN(\ab[0][12] ) );
  NOR2_X1 U663 ( .A1(n109), .A2(n104), .ZN(\ab[0][11] ) );
  NOR2_X1 U664 ( .A1(n108), .A2(n104), .ZN(\ab[0][10] ) );
  NOR2_X1 U665 ( .A1(n107), .A2(n104), .ZN(PRODUCT[0]) );
endmodule


module cortexm0ds_logic ( FCLK, SCLK, HCLK, DCLK, PORESETn, DBGRESETn, HRESETn, 
        SWCLKTCK, nTRST, HADDR, HBURST, HMASTLOCK, HPROT, HSIZE, HTRANS, 
        HWDATA, HWRITE, HRDATA, HREADY, HRESP, HMASTER, CODENSEQ, CODEHINTDE, 
        SPECHTRANS, SWDITMS, TDI, SWDO, SWDOEN, TDO, nTDOEN, DBGRESTART, 
        DBGRESTARTED, EDBGRQ, HALTED, NMI, IRQ, TXEV, RXEV, LOCKUP, 
        SYSRESETREQ, STCALIB, STCLKEN, IRQLATENCY, ECOREVNUM, GATEHCLK, 
        SLEEPING, SLEEPDEEP, WAKEUP, WICSENSE, SLEEPHOLDREQn, SLEEPHOLDACKn, 
        WICENREQ, WICENACK, CDBGPWRUPREQ, CDBGPWRUPACK, SE, RSTBYPASS, 
        vis_r0_o, vis_r1_o, vis_r2_o, vis_r3_o, vis_r4_o, vis_r5_o, vis_r6_o, 
        vis_r7_o, vis_r8_o, vis_r9_o, vis_r10_o, vis_r11_o, vis_r12_o, 
        vis_r14_o, vis_msp_o, vis_psp_o, vis_pc_o, vis_apsr_o, vis_tbit_o, 
        vis_ipsr_o, vis_control_o, vis_primask_o );
  output [31:0] HADDR;
  output [2:0] HBURST;
  output [3:0] HPROT;
  output [2:0] HSIZE;
  output [1:0] HTRANS;
  output [31:0] HWDATA;
  input [31:0] HRDATA;
  output [2:0] CODEHINTDE;
  input [31:0] IRQ;
  input [25:0] STCALIB;
  input [7:0] IRQLATENCY;
  input [27:0] ECOREVNUM;
  output [33:0] WICSENSE;
  output [31:0] vis_r0_o;
  output [31:0] vis_r1_o;
  output [31:0] vis_r2_o;
  output [31:0] vis_r3_o;
  output [31:0] vis_r4_o;
  output [31:0] vis_r5_o;
  output [31:0] vis_r6_o;
  output [31:0] vis_r7_o;
  output [31:0] vis_r8_o;
  output [31:0] vis_r9_o;
  output [31:0] vis_r10_o;
  output [31:0] vis_r11_o;
  output [31:0] vis_r12_o;
  output [31:0] vis_r14_o;
  output [29:0] vis_msp_o;
  output [29:0] vis_psp_o;
  output [30:0] vis_pc_o;
  output [3:0] vis_apsr_o;
  output [5:0] vis_ipsr_o;
  input FCLK, SCLK, HCLK, DCLK, PORESETn, DBGRESETn, HRESETn, SWCLKTCK, nTRST,
         HREADY, HRESP, SWDITMS, TDI, DBGRESTART, EDBGRQ, NMI, RXEV, STCLKEN,
         SLEEPHOLDREQn, WICENREQ, CDBGPWRUPACK, SE, RSTBYPASS;
  output HMASTLOCK, HWRITE, HMASTER, CODENSEQ, SPECHTRANS, SWDO, SWDOEN, TDO,
         nTDOEN, DBGRESTARTED, HALTED, TXEV, LOCKUP, SYSRESETREQ, GATEHCLK,
         SLEEPING, SLEEPDEEP, WAKEUP, SLEEPHOLDACKn, WICENACK, CDBGPWRUPREQ,
         vis_tbit_o, vis_control_o, vis_primask_o;
  wire   N427, n8369, n8370, n8371, n8372, n8373, n8374, n8375, n8376, n8377,
         n8378, HPROT_0, n8379, n8380, n8381, n8382, n8383, n8384, n8385,
         n8386, n8387, Qmdhu6, Pndhu6, Oodhu6, O5ohu6, G2ohu6, Q7ohu6, Dtnhu6,
         S3ohu6, \Aphpw6[2] , R9ohu6, Mzihu6, Eyihu6, Wwihu6, Ovihu6, Guihu6,
         Ysihu6, Qrihu6, Iqihu6, Apihu6, Snihu6, Kmihu6, Clihu6, Ujihu6,
         Miihu6, Ehihu6, Wfihu6, Oeihu6, Gdihu6, Ybihu6, Qaihu6, I9ihu6,
         A8ihu6, S6ihu6, K5ihu6, C4ihu6, U2ihu6, M1ihu6, E0ihu6, Wyhhu6,
         Oxhhu6, Gwhhu6, Edkhu6, Wbkhu6, N438, Oakhu6, G9khu6, Y7khu6, Q6khu6,
         I5khu6, M9ohu6, Uilhu6, Nhlhu6, Gglhu6, Zelhu6, Sdlhu6, Lclhu6,
         Eblhu6, W9lhu6, O8lhu6, G7lhu6, Y5lhu6, Q4lhu6, I3lhu6, A2lhu6,
         S0lhu6, Kzkhu6, Cykhu6, Uwkhu6, Mvkhu6, Eukhu6, Wskhu6, Orkhu6,
         Gqkhu6, Yokhu6, Qnkhu6, Imkhu6, Alkhu6, Sjkhu6, Kikhu6, Chkhu6,
         Ufkhu6, Avmhu6, Ttmhu6, N439, Msmhu6, Frmhu6, Ypmhu6, Romhu6, Knmhu6,
         Dqfhu6, Qbfpw6_10, Qbfpw6_5, Qbfpw6_4, Qbfpw6_3, Qbfpw6_2, Qbfpw6_1,
         Qbfpw6_0, D5epw6, I4epw6, B4epw6, U3epw6, N3epw6, G3epw6, Z2epw6,
         L2epw6, X1epw6, Q1epw6, J1epw6, C1epw6, Q5phu6, W4epw6, S2epw6,
         E2epw6, X3yhu6, O2yhu6, Hvxhu6, Avxhu6, Ytxhu6, Isxhu6, Sqxhu6,
         Xpxhu6, Qixhu6, Tgxhu6, Mgxhu6, Fgxhu6, Kfxhu6, Dfxhu6, Wexhu6,
         Pexhu6, Iexhu6, Bexhu6, Udxhu6, Ndxhu6, Gdxhu6, Zcxhu6, Scxhu6,
         Lcxhu6, Ecxhu6, Xbxhu6, Qbxhu6, Jbxhu6, Cbxhu6, Vaxhu6, Oaxhu6,
         Haxhu6, Aaxhu6, T9xhu6, M9xhu6, F9xhu6, Z5xhu6, L5xhu6, E5xhu6,
         Q4xhu6, J4xhu6, Cyohu6, Jyohu6, Qyohu6, Ezohu6, Lzohu6, Zzohu6,
         R2phu6, D2phu6, K2phu6, Y2phu6, F3phu6, A4phu6, H4phu6, V4phu6,
         Uwdpw6, Nwdpw6, Npghu6, W0xhu6, P0xhu6, I0xhu6, Mivhu6, Fivhu6,
         Yhvhu6, Pgvhu6, Igvhu6, Bgvhu6, Nfvhu6, Zevhu6, Sevhu6, Levhu6,
         Eevhu6, Xdvhu6, Jdvhu6, Cdvhu6, Vcvhu6, Ocvhu6, Davhu6, W9vhu6,
         P9vhu6, I9vhu6, B9vhu6, L7vhu6, Q6vhu6, J6vhu6, L0vhu6, Hyuhu6,
         Pvuhu6, Uuuhu6, Ztuhu6, Ltuhu6, Xsuhu6, Jsuhu6, Vruhu6, Vsthu6,
         Osthu6, Hsthu6, Asthu6, Trthu6, Kqthu6, Wpthu6, Ppthu6, Bpthu6,
         Uothu6, Nothu6, Gothu6, Znthu6, Snthu6, Lnthu6, Enthu6, Jmthu6,
         Cmthu6, Zgthu6, Sgthu6, Xfthu6, Cfthu6, Vethu6, Oethu6, Hethu6,
         Aethu6, Tdthu6, Mdthu6, Fdthu6, Ycthu6, Rcthu6, Kcthu6, Dcthu6,
         Wbthu6, Pbthu6, Ibthu6, Bbthu6, Uathu6, Nathu6, Gathu6, Z9thu6,
         S9thu6, L9thu6, E9thu6, X8thu6, Q8thu6, J8thu6, C8thu6, V7thu6,
         O7thu6, H7thu6, A7thu6, T6thu6, M6thu6, F6thu6, Y5thu6, R5thu6,
         K5thu6, D5thu6, W4thu6, P4thu6, I4thu6, B4thu6, U3thu6, N3thu6,
         G3thu6, Z2thu6, S2thu6, L2thu6, E2thu6, X1thu6, Q1thu6, J1thu6,
         C1thu6, V0thu6, O0thu6, H0thu6, A0thu6, Tzshu6, Mzshu6, Fzshu6,
         Yyshu6, Ryshu6, Kyshu6, Dyshu6, Wxshu6, Pxshu6, Ixshu6, Bxshu6,
         Uwshu6, Nwshu6, Gwshu6, Zvshu6, Svshu6, Lvshu6, Evshu6, Xushu6,
         Qushu6, Jushu6, Cushu6, Vtshu6, Otshu6, Atshu6, Tsshu6, Msshu6,
         Fsshu6, Yrshu6, Rrshu6, Krshu6, Drshu6, Wqshu6, Pqshu6, Iqshu6,
         Bqshu6, Upshu6, Npshu6, Gpshu6, Zoshu6, Soshu6, Eoshu6, Xnshu6,
         Qnshu6, Jnshu6, Cnshu6, Vmshu6, Omshu6, Hmshu6, Amshu6, Tlshu6,
         Mlshu6, Flshu6, Ykshu6, Rkshu6, Kkshu6, Dkshu6, Pjshu6, Ijshu6,
         Bjshu6, Uishu6, Nishu6, Gishu6, Zhshu6, Shshu6, Lhshu6, Ehshu6,
         Xgshu6, Qgshu6, Jgshu6, Cgshu6, Vfshu6, Ofshu6, Afshu6, Teshu6,
         Meshu6, Feshu6, Ydshu6, Rdshu6, Kdshu6, Ddshu6, Wcshu6, Pcshu6,
         Icshu6, Bcshu6, Ubshu6, Nbshu6, Gbshu6, Zashu6, Sashu6, Eashu6,
         X9shu6, Q9shu6, J9shu6, C9shu6, V8shu6, O8shu6, H8shu6, A8shu6,
         T7shu6, M7shu6, F7shu6, Y6shu6, R6shu6, K6shu6, D6shu6, P5shu6,
         I5shu6, B5shu6, U4shu6, N4shu6, G4shu6, Z3shu6, S3shu6, L3shu6,
         E3shu6, X2shu6, Q2shu6, J2shu6, C2shu6, V1shu6, O1shu6, A1shu6,
         T0shu6, M0shu6, F0shu6, Yzrhu6, Rzrhu6, Kzrhu6, Dzrhu6, Wyrhu6,
         Pyrhu6, Iyrhu6, Byrhu6, Uxrhu6, Nxrhu6, Gxrhu6, Zwrhu6, Swrhu6,
         Lwrhu6, Ewrhu6, Xvrhu6, Qvrhu6, Jvrhu6, Cvrhu6, Vurhu6, Ourhu6,
         Hurhu6, Aurhu6, Ttrhu6, Mtrhu6, Ftrhu6, Ysrhu6, Rsrhu6, Ksrhu6,
         Wrrhu6, Prrhu6, Brrhu6, Uqrhu6, Nqrhu6, Gqrhu6, Zprhu6, Sprhu6,
         Lprhu6, Eprhu6, Xorhu6, Qorhu6, Jorhu6, Corhu6, Vnrhu6, Onrhu6,
         Hnrhu6, Tmrhu6, Mmrhu6, Fmrhu6, Ylrhu6, Rlrhu6, Klrhu6, Dlrhu6,
         Wkrhu6, Pkrhu6, Ikrhu6, Bkrhu6, Ujrhu6, Njrhu6, Gjrhu6, Zirhu6,
         Sirhu6, Lirhu6, Xhrhu6, Qhrhu6, Jhrhu6, Chrhu6, Vgrhu6, Ogrhu6,
         Hgrhu6, Agrhu6, Tfrhu6, Mfrhu6, Ffrhu6, Yerhu6, Rerhu6, Kerhu6,
         Derhu6, Wdrhu6, Idrhu6, Bdrhu6, Ucrhu6, Ncrhu6, Gcrhu6, Zbrhu6,
         Sbrhu6, Lbrhu6, Ebrhu6, Xarhu6, Qarhu6, Jarhu6, Carhu6, V9rhu6,
         O9rhu6, H9rhu6, T8rhu6, M8rhu6, F8rhu6, Y7rhu6, R7rhu6, K7rhu6,
         D7rhu6, W6rhu6, P6rhu6, I6rhu6, B6rhu6, U5rhu6, N5rhu6, G5rhu6,
         Z4rhu6, S4rhu6, E4rhu6, X3rhu6, Q3rhu6, J3rhu6, C3rhu6, V2rhu6,
         O2rhu6, H2rhu6, A2rhu6, T1rhu6, M1rhu6, F1rhu6, Y0rhu6, R0rhu6,
         K0rhu6, D0rhu6, Pzqhu6, Izqhu6, Bzqhu6, Uyqhu6, Nyqhu6, Gyqhu6,
         Zxqhu6, Sxqhu6, Lxqhu6, Exqhu6, Xwqhu6, Qwqhu6, Jwqhu6, Cwqhu6,
         Vvqhu6, Ovqhu6, Avqhu6, Tuqhu6, Muqhu6, Fuqhu6, Ytqhu6, Rtqhu6,
         Ktqhu6, Dtqhu6, Wsqhu6, Psqhu6, Isqhu6, Bsqhu6, Urqhu6, Nrqhu6,
         Grqhu6, Zqqhu6, Lqqhu6, Eqqhu6, Xpqhu6, Qpqhu6, Jpqhu6, Cpqhu6,
         Voqhu6, Ooqhu6, Hoqhu6, Aoqhu6, Tnqhu6, Mnqhu6, Fnqhu6, Ymqhu6,
         Rmqhu6, Kmqhu6, Wlqhu6, Plqhu6, Ilqhu6, Blqhu6, Ukqhu6, Nkqhu6,
         Gkqhu6, Zjqhu6, Sjqhu6, Ljqhu6, Ejqhu6, Xiqhu6, Qiqhu6, Jiqhu6,
         Ciqhu6, Vhqhu6, Hhqhu6, Ahqhu6, Tgqhu6, Mgqhu6, Fgqhu6, Yfqhu6,
         Rfqhu6, Kfqhu6, Dfqhu6, Weqhu6, Peqhu6, Ieqhu6, Beqhu6, Udqhu6,
         Ndqhu6, Gdqhu6, Scqhu6, Lcqhu6, Ecqhu6, Xbqhu6, Qbqhu6, Jbqhu6,
         Cbqhu6, Vaqhu6, Oaqhu6, Haqhu6, Aaqhu6, T9qhu6, M9qhu6, F9qhu6,
         Y8qhu6, R8qhu6, D8qhu6, W7qhu6, P7qhu6, I7qhu6, B7qhu6, U6qhu6,
         N6qhu6, G6qhu6, Z5qhu6, S5qhu6, L5qhu6, E5qhu6, X4qhu6, Q4qhu6,
         J4qhu6, C4qhu6, O3qhu6, H3qhu6, A3qhu6, T2qhu6, M2qhu6, F2qhu6,
         Y1qhu6, R1qhu6, K1qhu6, D1qhu6, W0qhu6, P0qhu6, I0qhu6, B0qhu6,
         Uzphu6, Nzphu6, Zyphu6, Syphu6, Lyphu6, Eyphu6, Xxphu6, Qxphu6,
         Jxphu6, Cxphu6, Vwphu6, Owphu6, Hwphu6, Awphu6, Tvphu6, Mvphu6,
         Fvphu6, Yuphu6, Ruphu6, Duphu6, Wtphu6, Ptphu6, Itphu6, Btphu6,
         Usphu6, Nsphu6, Gsphu6, Zrphu6, Srphu6, Lrphu6, Erphu6, Xqphu6,
         Qqphu6, Jqphu6, Cqphu6, Opphu6, Hpphu6, Apphu6, Tophu6, Mophu6,
         Fophu6, Ynphu6, Rnphu6, Knphu6, Dnphu6, Wmphu6, Pmphu6, Imphu6,
         Bmphu6, Ulphu6, Nlphu6, Skphu6, Lkphu6, Ekphu6, Xjphu6, Qjphu6,
         Jjphu6, Cjphu6, Viphu6, Oiphu6, Hiphu6, Aiphu6, Thphu6, Mhphu6,
         Fhphu6, Ygphu6, Rgphu6, Kgphu6, Wfphu6, Pfphu6, Vxohu6, Oxohu6,
         Twohu6, Mwohu6, Fwohu6, Yvohu6, Rvohu6, Wuohu6, Ntohu6, Ssohu6,
         Lsohu6, Qrohu6, Jrohu6, Crohu6, Aqohu6, Miohu6, Gfohu6, Leohu6,
         Fmdhu6, N701, n25, n27, n28, n30, n31, n33, n36, n37, n38, n40, n41,
         n42, n47, n49, n51, n52, n53, n55, n56, n57, n61, n62, n63, n65, n66,
         n67, n68, n69, n70, n72, n73, n77, n79, n80, n81, n82, n84, n85, n87,
         n88, n89, n90, n93, n94, n95, n97, n98, n99, n100, n101, n102, n103,
         n104, n109, n110, n111, n113, n114, n115, n117, n118, n119, n122,
         n123, n124, n125, n127, n128, n129, n130, n131, n132, n133, n134,
         n135, n136, n137, n138, n139, n140, n141, n149, n150, n151, n152,
         n154, n155, n158, n159, n161, n162, n163, n164, n165, n167, n170,
         n171, n172, n173, n175, n176, n180, n181, n182, n183, n186, n187,
         n188, n189, n194, n197, n198, n199, n200, n201, n202, n203, n204,
         n205, n209, n210, n211, n212, n213, n216, n220, n223, n224, n227,
         n231, n232, n235, n238, n240, n241, n245, n246, n248, n251, n252,
         n255, n257, n258, n259, n262, n263, n264, n268, n269, n271, n273,
         n274, n275, n276, n278, n280, n282, n284, n286, n289, n291, n292,
         n294, n296, n297, n299, n301, n302, n304, n306, n307, n309, n311,
         n312, n315, n318, n319, n321, n324, n325, n327, n330, n331, n333,
         n336, n337, n340, n341, n342, n346, n347, n348, n351, n353, n354,
         n357, n358, n361, n362, n363, n367, n368, n369, n372, n374, n375,
         n378, n379, n381, n385, n386, n388, n392, n393, n395, n397, n401,
         n402, n404, n405, n406, n407, n409, n410, n411, n412, n413, n414,
         n415, n416, n417, n418, n419, n426, n427, n428, n429, n433, n434,
         n435, n440, n441, n443, n444, n445, n446, n447, n449, n452, n453,
         n454, n455, n457, n461, n462, n465, n466, n467, n469, n471, n472,
         n473, n474, n478, n480, n481, n483, n484, n487, n488, n489, n490,
         n493, n494, n495, n496, n497, n498, n499, n500, n501, n504, n506,
         n507, n509, n510, n511, n512, n513, n514, n515, n518, n519, n520,
         n525, n527, n528, n530, n531, n532, n533, n534, n535, n537, n539,
         n542, n543, n544, n545, n546, n548, n549, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n562, n566, n570, n571, n573,
         n574, n579, n580, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n600, n601, n603,
         n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
         n616, n618, n619, n620, n621, n622, n624, n626, n630, n633, n634,
         n636, n637, n638, n639, n641, n642, n643, n644, n645, n647, n648,
         n649, n651, n652, n653, n655, n656, n657, n658, n662, n663, n665,
         n666, n668, n673, n675, n676, n677, n689, n692, n693, n698, n699,
         n700, n702, n703, n705, n707, n708, n710, n711, n715, n716, n717,
         n718, n719, n720, n721, n723, n724, n725, n726, n727, n728, n730,
         n732, n735, n741, n742, n745, n746, n750, n752, n754, n756, n758,
         n759, n763, n765, n766, n769, n770, n773, n774, n777, n778, n781,
         n782, n785, n786, n789, n790, n792, n793, n795, n796, n797, n798,
         n801, n802, n804, n805, n806, n808, n810, n811, n812, n813, n814,
         n816, n817, n819, n820, n821, n822, n823, n825, n826, n827, n829,
         n831, n832, n834, n835, n837, n838, n839, n840, n842, n843, n844,
         n845, n846, n849, n851, n852, n853, n856, n858, n859, n860, n861,
         n862, n864, n865, n867, n868, n869, n870, n871, n873, n874, n876,
         n877, n879, n880, n882, n884, n886, n887, n888, n889, n893, n895,
         n896, n898, n899, n900, n901, n902, n903, n904, n905, n907, n909,
         n910, n911, n912, n914, n915, n916, n918, n919, n920, n921, n922,
         n923, n924, n925, n926, n927, n929, n930, n932, n933, n935, n936,
         n937, n938, n939, n940, n942, n943, n944, n945, n947, n948, n949,
         n951, n953, n954, n957, n958, n959, n960, n962, n965, n966, n967,
         n968, n969, n970, n971, n973, n978, n979, n980, n981, n982, n983,
         n984, n985, n987, n988, n989, n990, n991, n992, n993, n994, n996,
         n997, n998, n999, n1000, n1002, n1003, n1004, n1005, n1006, n1007,
         n1008, n1009, n1011, n1012, n1015, n1016, n1017, n1018, n1020, n1021,
         n1022, n1023, n1026, n1027, n1028, n1029, n1030, n1032, n1034, n1035,
         n1036, n1037, n1039, n1042, n1043, n1044, n1045, n1047, n1050, n1051,
         n1052, n1053, n1054, n1055, n1056, n1058, n1059, n1062, n1064, n1065,
         n1066, n1069, n1070, n1073, n1074, n1075, n1076, n1077, n1079, n1080,
         n1082, n1083, n1085, n1086, n1087, n1089, n1090, n1091, n1093, n1094,
         n1097, n1098, n1101, n1102, n1104, n1106, n1107, n1108, n1109, n1110,
         n1111, n1116, n1118, n1120, n1121, n1123, n1124, n1125, n1127, n1129,
         n1131, n1133, n1135, n1136, n1137, n1139, n1140, n1142, n1144, n1146,
         n1147, n1148, n1149, n1151, n1152, n1153, n1154, n1156, n1158, n1160,
         n1162, n1164, n1165, n1166, n1167, n1169, n1171, n1172, n1173, n1174,
         n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1186, n1189,
         n1191, n1192, n1193, n1194, n1195, n1196, n1199, n1200, n1201, n1202,
         n1203, n1204, n1206, n1207, n1208, n1209, n1211, n1213, n1214, n1215,
         n1216, n1217, n1218, n1219, n1220, n1222, n1223, n1224, n1225, n1227,
         n1228, n1229, n1230, n1232, n1234, n1235, n1237, n1238, n1239, n1240,
         n1241, n1242, n1244, n1245, n1246, n1247, n1248, n1249, n1251, n1253,
         n1255, n1258, n1260, n1262, n1263, n1264, n1265, n1266, n1267, n1269,
         n1270, n1271, n1272, n1273, n1274, n1275, n1277, n1278, n1280, n1281,
         n1282, n1283, n1284, n1287, n1290, n1291, n1292, n1293, n1294, n1295,
         n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1309,
         n1310, n1311, n1313, n1315, n1316, n1318, n1319, n1320, n1321, n1323,
         n1324, n1325, n1327, n1328, n1329, n1330, n1332, n1333, n1334, n1335,
         n1337, n1338, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348,
         n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360,
         n1361, n1362, n1363, n1364, n1365, n1366, n1369, n1371, n1373, n1374,
         n1376, n1377, n1378, n1379, n1383, n1385, n1387, n1389, n1390, n1391,
         n1392, n1394, n1396, n1398, n1400, n1403, n1404, n1407, n1408, n1410,
         n1411, n1412, n1413, n1414, n1417, n1418, n1419, n1422, n1424, n1425,
         n1426, n1428, n1430, n1431, n1433, n1435, n1436, n1437, n1438, n1439,
         n1440, n1441, n1442, n1443, n1444, n1445, n1451, n1452, n1453, n1454,
         n1455, n1456, n1457, n1458, n1459, n1461, n1462, n1463, n1464, n1465,
         n1466, n1468, n1470, n1471, n1473, n1474, n1475, n1477, n1478, n1479,
         n1480, n1482, n1483, n1486, n1487, n1488, n1489, n1493, n1494, n1495,
         n1496, n1497, n1498, n1499, n1501, n1502, n1503, n1504, n1505, n1511,
         n1512, n1513, n1518, n1519, n1520, n1521, n1522, n1524, n1528, n1531,
         n1532, n1533, n1534, n1535, n1536, n1538, n1539, n1540, n1541, n1546,
         n1547, n1548, n1549, n1550, n1554, n1555, n1556, n1557, n1558, n1559,
         n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569,
         n1570, n1571, n1572, n1576, n1577, n1578, n1579, n1583, n1584, n1585,
         n1586, n1587, n1588, n1589, n1591, n1592, n1593, n1594, n1595, n1598,
         n1599, n1600, n1601, n1602, n1605, n1607, n1609, n1611, n1612, n1613,
         n1615, n1617, n1619, n1620, n1621, n1622, n1623, n1624, n1625, n1626,
         n1627, n1628, n1629, n1630, n1634, n1635, n1636, n1638, n1640, n1641,
         n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1651, n1653,
         n1654, n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665, n1666,
         n1667, n1668, n1670, n1672, n1673, n1674, n1675, n1676, n1678, n1679,
         n1682, n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691,
         n1694, n1695, n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704,
         n1705, n1706, n1707, n1708, n1710, n1711, n1712, n1713, n1714, n1715,
         n1720, n1721, n1722, n1723, n1724, n1725, n1727, n1728, n1729, n1730,
         n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1739, n1740, n1741,
         n1742, n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751,
         n1752, n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761,
         n1762, n1763, n1765, n1768, n1771, n1773, n1776, n1777, n1778, n1781,
         n1784, n1787, n1789, n1792, n1794, n1796, n1797, n1800, n1803, n1806,
         n1807, n1810, n1813, n1816, n1818, n1821, n1824, n1827, n1830, n1833,
         n1835, n1836, n1839, n1842, n1845, n1848, n1850, n1853, n1854, n1856,
         n1857, n1858, n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867,
         n1868, n1869, n1870, n1871, n1872, n1873, n1874, n1875, n1876, n1877,
         n1878, n1879, n1880, n1881, n1882, n1883, n1884, n1886, n1887, n1890,
         n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1901,
         n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1911, n1912,
         n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922, n1924,
         n1928, n1929, n1930, n1931, n1932, n1933, n1935, n1937, n1938, n1940,
         n1941, n1942, n1943, n1944, n1946, n1948, n1949, n1950, n1951, n1952,
         n1953, n1954, n1955, n1956, n1957, n1959, n1960, n1961, n1962, n1963,
         n1965, n1966, n1968, n1969, n1971, n1972, n1973, n1976, n1977, n1978,
         n1980, n1981, n1982, n1983, n1984, n1985, n1987, n1988, n1990, n1991,
         n1992, n1993, n1995, n1996, n1997, n2005, n2006, n2007, n2008, n2010,
         n2011, n2013, n2014, n2015, n2017, n2019, n2021, n2023, n2025, n2027,
         n2029, n2030, n2032, n2034, n2036, n2038, n2039, n2040, n2042, n2043,
         n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053,
         n2054, n2056, n2057, n2058, n2059, n2060, n2061, n2063, n2064, n2065,
         n2066, n2067, n2068, n2071, n2072, n2073, n2074, n2077, n2079, n2081,
         n2083, n2085, n2087, n2089, n2091, n2093, n2095, n2097, n2099, n2101,
         n2103, n2105, n2106, n2108, n2109, n2112, n2113, n2114, n2115, n2116,
         n2117, n2120, n2123, n2127, n2129, n2132, n2134, n2137, n2141, n2144,
         n2147, n2149, n2151, n2152, n2153, n2154, n2155, n2156, n2157, n2159,
         n2160, n2162, n2165, n2166, n2168, n2169, n2170, n2171, n2172, n2174,
         n2177, n2178, n2179, n2180, n2182, n2183, n2184, n2186, n2187, n2188,
         n2192, n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201,
         n2202, n2205, n2209, n2210, n2213, n2214, n2217, n2218, n2221, n2223,
         n2225, n2228, n2229, n2230, n2231, n2236, n2237, n2239, n2240, n2241,
         n2245, n2248, n2249, n2252, n2253, n2255, n2257, n2259, n2261, n2263,
         n2264, n2269, n2271, n2274, n2276, n2278, n2284, n2285, n2288, n2289,
         n2292, n2295, n2297, n2299, n2300, n2302, n2303, n2305, n2306, n2307,
         n2308, n2311, n2314, n2315, n2318, n2319, n2321, n2323, n2325, n2327,
         n2329, n2331, n2333, n2335, n2337, n2340, n2343, n2344, n2348, n2352,
         n2354, n2356, n2357, n2359, n2362, n2369, n2371, n2372, n2373, n2374,
         n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382, n2386, n2393,
         n2394, n2395, n2399, n2401, n2404, n2405, n2407, n2408, n2409, n2410,
         n2412, n2414, n2417, n2421, n2422, n2424, n2426, n2430, n2431, n2434,
         n2439, n2441, n2446, n2448, n2450, n2452, n2453, n2454, n2455, n2461,
         n2463, n2465, n2467, n2469, n2471, n2472, n2480, n2482, n2483, n2484,
         n2487, n2488, n2489, n2491, n2492, n2493, n2494, n2495, n2496, n2497,
         n2498, n2499, n2501, n2503, n2504, n2505, n2518, n2520, n2521, n2523,
         n2525, n2526, n2531, n2532, n2534, n2536, n2540, n2542, n2552, n2554,
         n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562, n2563, n2564,
         n2565, n2566, n2567, n2568, n2570, n2571, n2573, n2574, n2576, n2577,
         n2578, n2579, n2580, n2581, n2583, n2585, n2586, n2587, n2588, n2589,
         n2592, n2593, n2600, n2602, n2604, n2611, n2612, n2613, n2618, n2619,
         n2620, n2621, n2622, n2623, n2624, n2625, n2626, n2627, n2628, n2629,
         n2630, n2631, n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640,
         n2641, n2642, n2643, n2658, n2659, n2661, n2662, n2665, n2668, n2669,
         n2672, n2673, n2677, n2680, n2681, n2683, n2685, n2687, n2695, n2701,
         n2704, n2705, n2706, n2707, n2709, n2733, n2734, n2735, n2736, n2737,
         n2738, n2739, n2740, n2741, n2742, n2743, n2744, n2746, n2747, n2748,
         n2749, n2750, n2751, n2752, n2753, n2754, n2755, n2756, n2760, n2761,
         n2762, n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2771, n2772,
         n2773, n2774, n2775, n2780, n2784, n2785, n2791, n2795, n2796, n2798,
         n2800, n2801, n2802, n2803, n2804, n2805, n2806, n2807, n2808, n2810,
         n2819, n2821, n2823, n2824, n2829, n2830, n2831, n2837, n2838, n2839,
         n2841, n2842, n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850,
         n2851, n2853, n2854, n2859, n2860, n2861, n2862, n2863, n2864, n2867,
         n2868, n2870, n2871, n2872, n2873, n2874, n2875, n2876, n2877, n2878,
         n2879, n2880, n2881, n2887, n2888, n2889, n2890, n2891, n2892, n2893,
         n2894, n2895, n2896, n2898, n2899, n2900, n2902, n2903, n2904, n2905,
         n2907, n2908, n2909, n2910, n2911, n2912, n2913, n2914, n2915, n2916,
         n2917, n2918, n2919, n2920, n2921, n2922, n2923, n2924, n2925, n2926,
         n2927, n2928, n2929, n2930, n2931, n2932, n2933, n2934, n2935, n2936,
         n2939, n2940, n2941, n2945, n2946, n2947, n2948, n2950, n2951, n2952,
         n2953, n2954, n2956, n2957, n2958, n2959, n2962, n2966, n2968, n2970,
         n2971, n2979, n2980, n2981, n2982, n2984, n2990, n2991, n2993, n2994,
         n2995, n2996, n2997, n2999, n3000, n3001, n3003, n3005, n3011, n3022,
         n3023, n3025, n3026, n3027, n3028, n3029, n3034, n3035, n3038, n3043,
         n3044, n3046, n3049, n3050, n3051, n3052, n3053, n3054, n3055, n3057,
         n3058, n3059, n3069, n3070, n3071, n3073, n3074, n3075, n3076, n3077,
         n3079, n3088, n3090, n3092, n3093, n3094, n3095, n3097, n3098, n3099,
         n3100, n3134, n3148, n3155, n3157, n3159, n3160, n3161, n3162, n3163,
         n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173,
         n3174, n3175, n3176, n3177, n3178, n3179, n3181, n3182, n3183, n3184,
         n3185, n3186, n3187, n3188, n3189, n3193, n3194, n3196, n3198, n3199,
         n3206, n3207, n3209, n3210, n3211, n3213, n3214, n3217, n3218, n3220,
         n3221, n3222, n3224, n3227, n3228, n3229, n3230, n3231, n3232, n3234,
         n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3243, n3244, n3245,
         n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3253, n3254, n3255,
         n3256, n3257, n3260, n3261, n3262, n3263, n3264, n3265, n3266, n3267,
         n3269, n3270, n3271, n3273, n3275, n3277, n3281, n3282, n3283, n3284,
         n3285, n3286, n3288, n3289, n3291, n3294, n3295, n3297, n3298, n3299,
         n3301, n3302, n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3311,
         n3312, n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321,
         n3322, n3323, n3325, n3326, n3327, n3328, n3330, n3331, n3332, n3333,
         n3334, n3336, n3338, n3339, n3340, n3342, n3344, n3345, n3346, n3348,
         n3349, n3350, n3352, n3353, n3354, n3355, n3356, n3357, n3359, n3360,
         n3361, n3362, n3363, n3364, n3365, n3366, n3367, n3368, n3370, n3371,
         n3372, n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381,
         n3382, n3383, n3384, n3385, n3386, n3387, n3390, n3391, n3392, n3393,
         n3394, n3395, n3396, n3398, n3399, n3400, n3401, n3402, n3403, n3406,
         n3407, n3408, n3409, n3410, n3411, n3412, n3413, n3414, n3415, n3416,
         n3417, n3418, n3420, n3421, n3422, n3423, n3424, n3425, n3426, n3427,
         n3428, n3429, n3430, n3431, n3432, n3433, n3434, n3435, n3436, n3437,
         n3438, n3440, n3442, n3445, n3447, n3448, n3449, n3452, n3455, n3457,
         n3458, n3459, n3461, n3462, n3463, n3464, n3465, n3466, n3469, n3477,
         n3485, n3487, n3489, n3490, n3491, n3492, n3493, n3494, n3495, n3496,
         n3497, n3498, n3499, n3500, n3501, n3502, n3504, n3506, n3507, n3508,
         n3509, n3510, n3511, n3512, n3513, n3514, n3515, n3516, n3517, n3518,
         n3519, n3521, n3522, n3523, n3524, n3525, n3526, n3527, n3528, n3529,
         n3530, n3531, n3536, n3537, n3539, n3541, n3542, n3552, n3553, n3555,
         n3557, n3558, n3559, n3560, n3561, n3562, n3563, n3564, n3565, n3567,
         n3568, n3569, n3570, n3572, n3573, n3574, n3575, n3577, n3578, n3579,
         n3580, n3582, n3584, n3585, n3589, n3590, n3594, n3595, n3597, n3599,
         n3600, n3603, n3605, n3606, n3609, n3610, n3612, n3613, n3615, n3616,
         n3619, n3621, n3622, n3624, n3626, n3627, n3629, n3632, n3633, n3636,
         n3637, n3639, n3641, n3642, n3644, n3646, n3647, n3649, n3651, n3652,
         n3655, n3657, n3658, n3660, n3662, n3663, n3665, n3667, n3670, n3671,
         n3674, n3675, n3677, n3678, n3679, n3680, n3681, n3683, n3685, n3687,
         n3688, n3689, n3691, n3692, n3693, n3694, n3695, n3696, n3700, n3704,
         n3708, n3711, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722,
         n3723, n3724, n3728, n3729, n3731, n3734, n3735, n3736, n3738, n3739,
         n3741, n3742, n3743, n3745, n3747, n3748, n3750, n3751, n3752, n3753,
         n3754, n3755, n3756, n3758, n3759, n3770, n3771, n3772, n3776, n3777,
         n3778, n3779, n3782, n3789, n3791, n3792, n3793, n3794, n3795, n3796,
         n3797, n3798, n3799, n3801, n3802, n3806, n3807, n3808, n3809, n3810,
         n3811, n3812, n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820,
         n3821, n3822, n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3834,
         n3839, n3842, n3844, n3847, n3848, n3850, n3852, n3853, n3854, n3856,
         n3857, n3859, n3861, n3862, n3872, n3873, n3874, n3876, n3878, n3881,
         n3885, n3887, n3888, n3889, n3891, n3892, n3893, n3896, n3897, n3898,
         n3900, n3901, n3902, n3903, n3905, n3906, n3907, n3908, n3909, n3910,
         n3912, n3914, n3916, n3917, n3918, n3919, n3920, n3921, n3923, n3927,
         n3929, n3932, n3933, n3941, n3942, n3943, n3944, n3945, n3949, n3950,
         n3953, n3956, n3958, n3962, n3963, n3964, n3965, n3966, n3969, n3970,
         n3974, n3976, n3982, n3991, n3992, n3993, n3994, n3995, n3996, n3997,
         n3998, n3999, n4000, n4012, n4013, n4014, n4019, n4020, n4021, n4023,
         n4025, n4026, n4030, n4031, n4037, n4039, n4043, n4045, n4047, n4050,
         n4051, n4056, n4057, n4058, n4059, n4060, n4062, n4064, n4065, n4067,
         n4068, n4069, n4071, n4073, n4074, n4075, n4076, n4077, n4079, n4080,
         n4081, n4082, n4083, n4084, n4085, n4087, n4088, n4089, n4090, n4091,
         n4092, n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101,
         n4102, n4103, n4104, n4105, n4106, n4107, n4108, n4113, n4114, n4120,
         n4121, n4122, n4124, n4125, n4127, n4128, n4129, n4130, n4131, n4132,
         n4133, n4137, n4143, n4147, n4148, n4150, n4153, n4154, n4155, n4156,
         n4159, n4162, n4165, n4166, n4168, n4169, n4171, n4173, n4174, n4175,
         n4176, n4177, n4183, n4191, n4192, n4197, n4198, n4200, n4201, n4206,
         n4207, n4208, n4209, n4210, n4211, n4212, n4213, n4214, n4216, n4217,
         n4218, n4219, n4220, n4221, n4223, n4224, n4225, n4226, n4227, n4228,
         n4230, n4231, n4233, n4234, n4235, n4236, n4238, n4239, n4241, n4242,
         n4243, n4247, n4248, n4249, n4251, n4252, n4253, n4254, n4255, n4256,
         n4257, n4258, n4259, n4260, n4261, n4262, n4264, n4266, n4267, n4268,
         n4269, n4270, n4274, n4276, n4277, n4279, n4283, n4284, n4286, n4287,
         n4288, n4289, n4290, n4291, n4292, n4294, n4295, n4296, n4298, n4299,
         n4300, n4302, n4303, n4304, n4305, n4307, n4308, n4309, n4310, n4311,
         n4312, n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321,
         n4322, n4323, n4325, n4326, n4327, n4328, n4331, n4332, n4334, n4337,
         n4338, n4339, n4340, n4342, n4343, n4344, n4345, n4346, n4347, n4349,
         n4350, n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361,
         n4362, n4363, n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372,
         n4373, n4374, n4375, n4377, n4380, n4381, n4382, n4383, n4384, n4385,
         n4386, n4387, n4388, n4389, n4390, n4391, n4392, n4393, n4396, n4397,
         n4398, n4399, n4400, n4401, n4403, n4404, n4407, n4411, n4412, n4413,
         n4414, n4415, n4416, n4417, n4418, n4419, n4421, n4422, n4423, n4424,
         n4425, n4426, n4427, n4428, n4429, n4430, n4438, n4439, n4440, n4443,
         n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4455,
         n4456, n4457, n4458, n4461, n4462, n4463, n4464, n4469, n4471, n4472,
         n4475, n4476, n4477, n4479, n4480, n4481, n4483, n4484, n4485, n4486,
         n4488, n4489, n4490, n4492, n4493, n4494, n4495, n4496, n4497, n4498,
         n4499, n4500, n4501, n4502, n4503, n4504, n4505, n4508, n4509, n4510,
         n4511, n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4522,
         n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532,
         n4533, n4534, n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543,
         n4544, n4547, n4549, n4550, n4551, n4552, n4553, n4556, n4557, n4558,
         n4559, n4560, n4561, n4562, n4563, n4565, n4567, n4568, n4569, n4570,
         n4571, n4573, n4574, n4575, n4576, n4577, n4578, n4580, n4581, n4582,
         n4583, n4584, n4585, n4586, n4589, n4590, n4592, n4593, n4594, n4595,
         n4596, n4597, n4599, n4600, n4601, n4603, n4604, n4605, n4606, n4607,
         n4609, n4612, n4613, n4614, n4615, n4617, n4618, n4619, n4620, n4621,
         n4622, n4623, n4624, n4625, n4626, n4627, n4629, n4630, n4632, n4634,
         n4636, n4638, n4639, n4640, n4641, n4643, n4644, n4645, n4646, n4647,
         n4648, n4649, n4652, n4653, n4654, n4655, n4656, n4657, n4659, n4660,
         n4661, n4662, n4663, n4664, n4665, n4666, n4671, n4675, n4676, n4677,
         n4678, n4679, n4680, n4681, n4682, n4683, n4684, n4686, n4689, n4690,
         n4691, n4692, n4696, n4697, n4698, n4705, n4706, n4709, n4710, n4711,
         n4712, n4714, n4715, n4716, n4717, n4718, n4719, n4722, n4723, n4726,
         n4727, n4728, n4729, n4730, n4731, n4733, n4734, n4735, n4736, n4737,
         n4739, n4740, n4741, n4742, n4743, n4744, n4745, n4746, n4747, n4748,
         n4750, n4751, n4752, n4754, n4755, n4757, n4758, n4759, n4760, n4762,
         n4763, n4767, n4768, n4769, n4770, n4771, n4775, n4778, n4779, n4780,
         n4781, n4784, n4785, n4786, n4788, n4789, n4790, n4791, n4792, n4793,
         n4794, n4796, n4798, n4800, n4803, n4804, n4808, n4809, n4812, n4813,
         n4814, n4815, n4817, n4819, n4820, n4821, n4822, n4823, n4824, n4825,
         n4827, n4828, n4829, n4830, n4831, n4832, n4833, n4834, n4835, n4836,
         n4837, n4838, n4840, n4842, n4843, n4844, n4845, n4846, n4847, n4848,
         n4849, n4850, n4851, n4852, n4853, n4854, n4856, n4857, n4858, n4859,
         n4860, n4861, n4862, n4863, n4864, n4865, n4866, n4867, n4868, n4869,
         n4870, n4871, n4872, n4873, n4874, n4875, n4876, n4877, n4878, n4879,
         n4880, n4881, n4882, n4883, n4884, n4885, n4886, n4887, n4888, n4889,
         n4890, n4891, n4892, n4893, n4894, n4895, n4896, n4897, n4898, n4899,
         n4900, n4901, n4902, n4903, n4904, n4905, n4906, n4909, n4911, n4912,
         n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922,
         n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4933,
         n4934, n4935, n4936, n4937, n4938, n4939, n4941, n4942, n4943, n4944,
         n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952, n4953, n4954,
         n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962, n4963, n4964,
         n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972, n4973, n4974,
         n4975, n4976, n4977, n4979, n4980, n4981, n4982, n4983, n4984, n4985,
         n4986, n4988, n4989, n4990, n4991, n4992, n4994, n4995, n4996, n4997,
         n4998, n4999, n5000, n5001, n5003, n5004, n5005, n5006, n5007, n5008,
         n5009, n5010, n5011, n5012, n5013, n5014, n5015, n5016, n5017, n5018,
         n5019, n5020, n5021, n5022, n5023, n5024, n5025, n5026, n5027, n5028,
         n5029, n5030, n5031, n5032, n5033, n5034, n5035, n5036, n5038, n5039,
         n5040, n5041, n5043, n5044, n5045, n5046, n5048, n5049, n5050, n5051,
         n5052, n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061,
         n5062, n5064, n5066, n5067, n5068, n5069, n5071, n5072, n5073, n5075,
         n5076, n5077, n5078, n5079, n5080, n5081, n5082, n5083, n5084, n5085,
         n5086, n5087, n5089, n5090, n5091, n5092, n5093, n5094, n5095, n5096,
         n5097, n5098, n5099, n5100, n5101, n5102, n5103, n5104, n5106, n5107,
         n5108, n5109, n5110, n5113, n5114, n5115, n5116, n5117, n5118, n5119,
         n5120, n5121, n5122, n5123, n5124, n5125, n5127, n5130, n5131, n5132,
         n5133, n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142, n5143,
         n5144, n5145, n5146, n5147, n5149, n5150, n5151, n5152, n5153, n5155,
         n5156, n5157, n5158, n5159, n5160, n5161, n5162, n5163, n5164, n5165,
         n5166, n5167, n5168, n5169, n5170, n5171, n5172, n5173, n5174, n5176,
         n5177, n5178, n5179, n5181, n5182, n5183, n5184, n5185, n5186, n5187,
         n5188, n5189, n5190, n5191, n5194, n5195, n5196, n5199, n5200, n5201,
         n5202, n5203, n5204, n5205, n5206, n5207, n5208, n5211, n5212, n5213,
         n5214, n5215, n5217, n5218, n5219, n5220, n5221, n5222, n5223, n5224,
         n5226, n5227, n5228, n5229, n5230, n5231, n5232, n5233, n5234, n5235,
         n5238, n5239, n5240, n5241, n5242, n5243, n5244, n5245, n5246, n5247,
         n5248, n5249, n5250, n5251, n5252, n5253, n5254, n5255, n5259, n5260,
         n5261, n5262, n5263, n5264, n5265, n5267, n5268, n5269, n5271, n5274,
         n5275, n5276, n5279, n5280, n5281, n5283, n5285, n5286, n5287, n5288,
         n5289, n5290, n5292, n5295, n5296, n5297, n5298, n5300, n5301, n5303,
         n5305, n5306, n5308, n5309, n5310, n5311, n5314, n5315, n5316, n5318,
         n5320, n5321, n5322, n5323, n5324, n5325, n5327, n5328, n5329, n5330,
         n5331, n5332, n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342,
         n5343, n5344, n5345, n5346, n5347, n5349, n5350, n5351, n5353, n5354,
         n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362, n5363, n5364,
         n5365, n5367, n5368, n5371, n5373, n5374, n5375, n5376, n5377, n5378,
         n5379, n5380, n5381, n5382, n5383, n5384, n5385, n5387, n5388, n5389,
         n5390, n5391, n5392, n5393, n5395, n5396, n5397, n5398, n5399, n5400,
         n5401, n5402, n5404, n5405, n5406, n5407, n5408, n5412, n5413, n5414,
         n5415, n5416, n5417, n5418, n5420, n5421, n5422, n5423, n5424, n5425,
         n5426, n5429, n5430, n5431, n5432, n5434, n5435, n5436, n5437, n5438,
         n5439, n5440, n5441, n5442, n5443, n5444, n5445, n5446, n5447, n5448,
         n5450, n5452, n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5466,
         n5469, n5471, n5472, n5473, n5474, n5475, n5476, n5477, n5478, n5479,
         n5480, n5481, n5482, n5483, n5486, n5487, n5488, n5489, n5490, n5491,
         n5492, n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502,
         n5503, n5504, n5505, n5508, n5509, n5510, n5511, n5512, n5513, n5514,
         n5515, n5516, n5517, n5518, n5519, n5524, n5525, n5527, n5528, n5529,
         n5530, n5531, n5533, n5535, n5536, n5537, n5538, n5539, n5542, n5543,
         n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5553, n5554, n5557,
         n5558, n5559, n5560, n5561, n5563, n5564, n5565, n5566, n5567, n5568,
         n5569, n5570, n5571, n5572, n5573, n5574, n5575, n5576, n5577, n5578,
         n5581, n5582, n5583, n5585, n5586, n5587, n5588, n5589, n5590, n5591,
         n5592, n5593, n5594, n5595, n5596, n5597, n5599, n5600, n5601, n5602,
         n5603, n5604, n5605, n5607, n5608, n5609, n5610, n5611, n5612, n5613,
         n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622, n5623,
         n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632, n5633, n5634,
         n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5643, n5644, n5645,
         n5646, n5647, n5648, n5649, n5650, n5651, n5652, n5653, n5655, n5656,
         n5657, n5658, n5659, n5660, n5661, n5664, n5665, n5666, n5667, n5668,
         n5670, n5671, n5672, n5674, n5675, n5677, n5678, n5679, n5680, n5681,
         n5685, n5686, n5687, n5688, n5690, n5691, n5692, n5693, n5694, n5695,
         n5696, n5697, n5698, n5699, n5700, n5701, n5702, n5703, n5704, n5705,
         n5706, n5707, n5708, n5712, n5713, n5714, n5715, n5716, n5717, n5719,
         n5720, n5721, n5722, n5723, n5724, n5727, n5728, n5731, n5732, n5733,
         n5734, n5735, n5737, n5738, n5740, n5741, n5742, n5743, n5744, n5745,
         n5746, n5747, n5748, n5749, n5750, n5751, n5753, n5754, n5755, n5756,
         n5757, n5758, n5759, n5760, n5761, n5762, n5763, n5764, n5765, n5766,
         n5767, n5768, n5769, n5770, n5771, n5772, n5773, n5774, n5775, n5776,
         n5777, n5778, n5779, n5780, n5781, n5782, n5783, n5784, n5785, n5786,
         n5787, n5788, n5790, n5791, n5792, n5795, n5796, n5797, n5798, n5800,
         n5801, n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5812, n5813,
         n5815, n5816, n5817, n5818, n5819, n5821, n5823, n5824, n5826, n5827,
         n5828, n5830, n5831, n5833, n5835, n5836, n5837, n5838, n5840, n5841,
         n5842, n5843, n5844, n5845, n5847, n5850, n5852, n5853, n5854, n5855,
         n5856, n5857, n5858, n5861, n5862, n5863, n5864, n5866, n5867, n5868,
         n5869, n5870, n5871, n5874, n5878, n5879, n5880, n5881, n5882, n5883,
         n5884, n5885, n5888, n5889, n5890, n5893, n5896, n5900, n5902, n5903,
         n5904, n5906, n5907, n5908, n5909, n5910, n5911, n5912, n5913, n5916,
         n5917, n5918, n5919, n5920, n5921, n5922, n5923, n5925, n5926, n5927,
         n5929, n5930, n5931, n5932, n5933, n5934, n5936, n5942, n5943, n5944,
         n5945, n5946, n5947, n5949, n5950, n5951, n5952, n5953, n5954, n5957,
         n5958, n5962, n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972,
         n5973, n5974, n5975, n5977, n5978, n5979, n5980, n5981, n5982, n5983,
         n5984, n5985, n5986, n5987, n5988, n5991, n5992, n5994, n5995, n5996,
         n5997, n5998, n5999, n6000, n6001, n6002, n6003, n6004, n6005, n6006,
         n6007, n6008, n6009, n6010, n6011, n6012, n6013, n6014, n6015, n6016,
         n6017, n6018, n6019, n6020, n6021, n6022, n6023, n6024, n6025, n6026,
         n6027, n6028, n6029, n6030, n6031, n6032, n6033, n6034, n6035, n6036,
         n6037, n6038, n6040, n6041, n6042, n6043, n6044, n6045, n6046, n6047,
         n6048, n6049, n6050, n6051, n6052, n6053, n6054, n6055, n6056, n6057,
         n6058, n6059, n6060, n6061, n6062, n6063, n6064, n6065, n6066, n6067,
         n6068, n6069, n6070, n6071, n6072, n6073, n6074, n6075, n6076, n6077,
         n6078, n6079, n6081, n6082, n6083, n6084, n6085, n6086, n6087, n6088,
         n6089, n6090, n6091, n6092, n6093, n6094, n6095, n6096, n6097, n6098,
         n6099, n6100, n6101, n6102, n6103, n6106, n6107, n6108, n6109, n6110,
         n6111, n6112, n6113, n6114, n6115, n6116, n6117, n6118, n6123, n6125,
         n6126, n6127, n6130, n6131, n6132, n6133, n6134, n6135, n6137, n6139,
         n6140, n6141, n6143, n6145, n6147, n6149, n6154, n6155, n6157, n6158,
         n6159, n6160, n6161, n6162, n6163, n6164, n6165, n6166, n6169, n6170,
         n6171, n6172, n6173, n6174, n6179, n6180, n6181, n6182, n6184, n6185,
         n6186, n6187, n6189, n6190, n6191, n6192, n6193, n6194, n6195, n6196,
         n6197, n6198, n6199, n6200, n6201, n6203, n6204, n6205, n6206, n6208,
         n6209, n6211, n6213, n6214, n6215, n6216, n6217, n6222, n6223, n6224,
         n6226, n6227, n6228, n6230, n6231, n6232, n6233, n6235, n6236, n6237,
         n6238, n6240, n6243, n6244, n6245, n6246, n6247, n6248, n6250, n6251,
         n6252, n6254, n6255, n6256, n6258, n6259, n6261, n6262, n6263, n6265,
         n6268, n6269, n6270, n6272, n6273, n6274, n6275, n6276, n6277, n6278,
         n6279, n6282, n6283, n6284, n6285, n6286, n6287, n6288, n6293, n6295,
         n6296, n6297, n6298, n6299, n6300, n6301, n6302, n6303, n6304, n6305,
         n6307, n6308, n6309, n6310, n6311, n6312, n6314, n6315, n6316, n6318,
         n6319, n6320, n6321, n6322, n6323, n6325, n6326, n6327, n6332, n6333,
         n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6342, n6343, n6344,
         n6345, n6346, n6347, n6348, n6350, n6353, n6354, n6356, n6357, n6358,
         n6359, n6360, n6361, n6362, n6363, n6364, n6366, n6367, n6368, n6369,
         n6370, n6371, n6373, n6374, n6375, n6376, n6379, n6381, n6382, n6383,
         n6384, n6385, n6388, n6389, n6390, n6391, n6392, n6393, n6396, n6397,
         n6398, n6400, n6401, n6402, n6403, n6404, n6405, n6406, n6407, n6408,
         n6409, n6410, n6411, n6412, n6413, n6414, n6415, n6416, n6417, n6418,
         n6419, n6420, n6421, n6422, n6423, n6424, n6426, n6427, n6428, n6429,
         n6430, n6431, n6432, n6433, n6434, n6435, n6436, n6437, n6438, n6439,
         n6440, n6441, n6442, n6443, n6444, n6445, n6446, n6447, n6448, n6449,
         n6450, n6451, n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460,
         n6461, n6462, n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470,
         n6471, n6472, n6473, n6474, n6475, n6476, n6477, n6481, n6482, n6483,
         n6485, n6488, n6489, n6490, n6491, n6492, n6493, n6494, n6495, n6496,
         n6497, n6498, n6499, n6500, n6501, n6502, n6503, n6505, n6506, n6507,
         n6508, n6509, n6510, n6511, n6512, n6513, n6514, n6515, n6516, n6517,
         n6519, n6520, n6521, n6522, n6523, n6525, n6527, n6528, n6529, n6530,
         n6531, n6532, n6533, n6534, n6535, n6536, n6538, n6539, n6540, n6541,
         n6542, n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551,
         n6552, n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6561, n6562,
         n6563, n6565, n6566, n6567, n6568, n6569, n6572, n6573, n6575, n6576,
         n6578, n6579, n6580, n6581, n6582, n6584, n6587, n6589, n6591, n6592,
         n6593, n6594, n6596, n6597, n6598, n6601, n6602, n6604, n6606, n6608,
         n6609, n6610, n6611, n6612, n6613, n6614, n6615, n6616, n6617, n6618,
         n6619, n6620, n6621, n6622, n6623, n6624, n6625, n6627, n6629, n6630,
         n6631, n6632, n6633, n6634, n6635, n6637, n6640, n6641, n6643, n6644,
         n6645, n6647, n6648, n6649, n6651, n6652, n6653, n6654, n6655, n6656,
         n6658, n6659, n6660, n6661, n6662, n6664, n6665, n6666, n6667, n6670,
         n6671, n6672, n6673, n6675, n6676, n6679, n6680, n6681, n6682, n6683,
         n6684, n6685, n6687, n6688, n6689, n6690, n6691, n6692, n6693, n6694,
         n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702, n6703, n6704,
         n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712, n6713, n6714,
         n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722, n6723, n6724,
         n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732, n6733, n6734,
         n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742, n6743, n6744,
         n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752, n6753, n6754,
         n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762, n6763, n6764,
         n6765, n6766, n6767, n6768, n6769, n6770, n6772, n6773, n6774, n6775,
         n6776, n6777, n6778, n6779, n6780, n6781, n6782, n6783, n6784, n6785,
         n6786, n6787, n6788, n6789, n6790, n6791, n6792, n6793, n6794, n6795,
         n6796, n6797, n6798, n6799, n6800, n6801, n6802, n6803, n6804, n6805,
         n6806, n6807, n6808, n6809, n6811, n6812, n6813, n6814, n6815, n6816,
         n6817, n6818, n6820, n6821, n6822, n6823, n6824, n6825, n6827, n6828,
         n6829, n6830, n6831, n6832, n6833, n6834, n6836, n6837, n6838, n6839,
         n6840, n6841, n6842, n6843, n6844, n6845, n6846, n6847, n6848, n6849,
         n6850, n6851, n6852, n6853, n6854, n6855, n6856, n6857, n6858, n6859,
         n6860, n6861, n6862, n6864, n6865, n6866, n6867, n6868, n6869, n6870,
         n6872, n6873, n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881,
         n6882, n6883, n6884, n6885, n6887, n6888, n6889, n6890, n6891, n6892,
         n6893, n6894, n6895, n6896, n6897, n6898, n6900, n6901, n6902, n6903,
         n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912, n6913,
         n6914, n6915, n6916, n6917, n6919, n6920, n6921, n6922, n6923, n6924,
         n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932, n6933, n6934,
         n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942, n6943, n6944,
         n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952, n6953, n6954,
         n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962, n6963, n6964,
         n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972, n6973, n6974,
         n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982, n6983, n6984,
         n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992, n6993, n6994,
         n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002, n7003, n7004,
         n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012, n7013, n7014,
         n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022, n7023, n7024,
         n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7032, n7033, n7034,
         n7035, n7036, n7037, n7038, n7039, n7040, n7041, n7042, n7043, n7044,
         n7045, n7046, n7047, n7048, n7049, n7050, n7051, n7052, n7053, n7054,
         n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062, n7063, n7064,
         n7065, n7066, n7067, n7068, n7069, n7070, n7071, n7072, n7073, n7074,
         n7075, n7076, n7077, n7078, n7079, n7080, n7081, n7082, n7083, n7084,
         n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092, n7093, n7094,
         n7095, n7096, n7097, n7098, n7099, n7100, n7101, n7102, n7103, n7104,
         n7105, n7106, n7107, n7108, n7109, n7110, n7111, n7112, n7113, n7114,
         n7115, n7116, n7117, n7118, n7119, n7120, n7121, n7122, n7123, n7124,
         n7125, n7126, n7127, n7128, n7129, n7130, n7131, n7132, n7133, n7134,
         n7135, n7136, n7137, n7138, n7139, n7140, n7141, n7142, n7143, n7144,
         n7145, n7146, n7147, n7148, n7149, n7150, n7151, n7152, n7153, n7154,
         n7155, n7156, n7157, n7158, n7159, n7160, n7161, n7162, n7163, n7164,
         n7165, n7166, n7167, n7168, n7169, n7170, n7171, n7172, n7173, n7174,
         n7175, n7176, n7177, n7178, n7179, n7180, n7181, n7182, n7183, n7184,
         n7185, n7186, n7187, n7188, n7189, n7190, n7191, n7192, n7193, n7194,
         n7195, n7196, n7197, n7198, n7199, n7200, n7201, n7202, n7203, n7204,
         n7205, n7206, n7207, n7208, n7209, n7210, n7211, n7212, n7213, n7214,
         n7215, n7216, n7217, n7218, n7219, n7220, n7221, n7222, n7223, n7224,
         n7225, n7226, n7227, n7228, n7229, n7230, n7231, n7232, n7233, n7234,
         n7235, n7236, n7237, n7238, n7239, n7240, n7241, n7242, n7243, n7244,
         n7245, n7246, n7247, n7248, n7249, n7250, n7251, n7252, n7253, n7254,
         n7255, n7256, n7257, n7258, n7259, n7260, n7262, n7263, n7264, n7265,
         n7266, n7267, n7268, n7269, n7270, n7271, n7272, n7273, n7274, n7275,
         n7276, n7277, n7278, n7279, n7280, n7281, n7282, n7283, n7284, n7285,
         n7286, n7287, n7288, n7289, n7290, n7291, n7292, n7293, n7294, n7295,
         n7296, n7297, n7298, n7299, n7300, n7301, n7302, n7303, n7304, n7305,
         n7306, n7308, n7309, n7310, n7311, n7312, n7313, n7314, n7315, n7316,
         n7317, n7318, n7319, n7320, n7321, n7322, n7323, n7324, n7325, n7326,
         n7327, n7328, n7329, n7330, n7331, n7332, n7333, n7334, n7335, n7336,
         n7337, n7338, n7339, n7340, n7343, n7344, n7345, n7346, n7347, n7348,
         n7349, n7350, n7351, n7352, n7353, n7354, n7355, n7356, n7357, n7358,
         n7359, n7360, n7361, n7362, n7363, n7364, n7365, n7366, n7367, n7368,
         n7369, n7371, n7373, n7374, n7375, n7378, n7379, n7380, n7381, n7382,
         n7383, n7384, n7385, n7386, n7387, n7388, n7389, n7390, n7391, n7392,
         n7393, n7394, n7395, n7396, n7397, n7398, n7399, n7400, n7401, n7402,
         n7403, n7404, n7405, n7406, n7407, n7408, n7409, n7410, n7411, n7412,
         n7413, n7414, n7415, n7416, n7417, n7418, n7419, n7420, n7421, n7422,
         n7423, n7424, n7425, n7426, n7427, n7428, n7429, n7430, n7431, n7432,
         n7433, n7434, n7435, n7436, n7437, n7438, n7439, n7440, n7441, n7442,
         n7443, n7444, n7445, n7446, n7447, n7448, n7449, n7450, n7451, n7452,
         n7453, n7454, n7455, n7456, n7457, n7458, n7459, n7460, n7461, n7462,
         n7463, n7464, n7465, n7466, n7467, n7468, n7469, n7470, n7471, n7472,
         n7473, n7474, n7475, n7476, n7477, n7478, n7479, n7480, n7481, n7482,
         n7483, n7484, n7485, n7486, n7487, n7488, n7489, n7490, n7491, n7492,
         n7493, n7494, n7495, n7496, n7497, n7498, n7499, n7500, n7501, n7502,
         n7503, n7504, n7505, n7506, n7507, n7508, n7509, n7510, n7511, n7513,
         n7514, n7515, n7516, n7517, n7518, n7519, n7520, n7521, n7522, n7523,
         n7524, n7525, n7526, n7527, n7528, n7529, n7530, n7531, n7532, n7533,
         n7534, n7535, n7536, n7537, n7538, n7539, n7540, n7541, n7542, n7543,
         n7544, n7545, n7546, n7547, n7548, n7549, n7550, n7551, n7552, n7553,
         n7554, n7555, n7556, n7557, n7558, n7559, n7560, n7561, n7562, n7563,
         n7564, n7565, n7566, n7567, n7568, n7569, n7570, n7572, n7574, n7576,
         n7581, n7582, n7583, n7584, n7585, n7586, n7587, n7588, n7589, n7590,
         n7591, n7592, n7593, n7594, n7595, n7596, n7597, n7598, n7599, n7601,
         n7602, n7604, n7605, n7606, n7607, n7608, n7609, n7610, n7611, n7612,
         n7613, n7614, n7615, n7616, n7617, n7618, n7619, n7620, n7621, n7622,
         n7623, n7624, n7625, n7626, n7627, n7628, n7629, n7630, n7631, n7632,
         n7633, n7634, n7635, n7636, n7637, n7638, n7639, n7640, n7641, n7642,
         n7645, n7646, n7647, n7648, n7649, n7650, n7651, n7652, n7653, n7654,
         n7655, n7656, n7657, n7658, n7659, n7660, n7661, n7662, n7663, n7664,
         n7665, n7666, n7667, n7669, n7670, n7671, n7672, n7673, n7674, n7675,
         n7676, n7677, n7678, n7679, n7680, n7681, n7682, n7683, n7684, n7685,
         n7686, n7687, n7688, n7689, n7690, n7691, n7692, n7693, n7694, n7696,
         n7697, n7698, n7699, n7700, n7701, n7702, n7703, n7705, n7706, n7707,
         n7708, n7709, n7710, n7711, n7712, n7713, n7714, n7715, n7716, n7717,
         n7718, n7719, n7720, n7721, n7722, n7723, n7724, n7725, n7726, n7727,
         n7728, n7729, n7730, n7731, n7732, n7733, n7734, n7735, n7736, n7737,
         n7738, n7739, n7740, n7741, n7742, n7743, n7744, n7746, n7747, n7749,
         n7750, n7752, n7753, n7755, n7756, n7758, n7759, n7761, n7762, n7764,
         n7765, n7767, n7768, n7770, n7771, n7773, n7774, n7776, n7777, n7779,
         n7780, n7782, n7783, n7785, n7786, n7788, n7789, n7791, n7792, n7794,
         n7795, n7796, n7798, n7799, n7801, n7803, n7804, n7805, n7807, n7808,
         n7810, n7812, n7813, n7814, n7816, n7817, n7819, n7820, n7822, n7823,
         n7825, n7826, n7827, n7828, n7829, n7830, n7831, n7832, n7833, n7834,
         n7835, n7836, n7837, n7838, n7839, n7840, n7841, n7842, n7843, n7844,
         n7845, n7846, n7847, n7848, n7849, n7850, n7851, n7852, n7853, n7854,
         n7855, n7856, n7857, n7858, n7859, n7860, n7861, n7862, n7863, n7864,
         n7865, n7866, n7867, n7868, n7869, n7870, n7871, n7872, n7873, n7874,
         n7875, n7876, n7877, n7878, n7879, n7880, n7881, n7882, n7883, n7884,
         n7885, n7886, n7887, n7888, n7889, n7890, n7891, n7892, n7893, n7894,
         n7895, n7896, n7897, n7898, n7899, n7900, n7901, n7902, n7903, n7904,
         n7905, n7906, n7907, n7908, n7909, n7910, n7911, n7912, n7913, n7914,
         n7915, n7916, n7917, n7918, n7919, n7920, n7921, n7923, n7924, n7925,
         n7926, n7927, n7928, n7929, n7930, n7931, n7932, n7933, n7934, n7935,
         n7936, n7937, n7938, n7939, n7940, n7941, n7942, n7943, n7944, n7945,
         n7946, n7947, n7948, n7949, n7950, n7951, n7952, n7953, n7954, n7955,
         n7956, n7957, n7958, n7959, n7960, n7961, n7962, n7963, n7964, n7965,
         n7966, n7967, n7968, n7969, n7970, n7971, n7972, n7973, n7974, n7975,
         n7976, n7977, n7978, n7979, n7980, n7981, n7982, n7983, n7984, n7985,
         n7986, n7987, n7988, n7989, n7990, n7991, n7992, n7993, n7994, n7995,
         n7996, n7997, n7998, n7999, n8000, n8001, n8002, n8003, n8004, n8005,
         n8006, n8007, n8009, n8010, n8011, n8012, n8013, n8014, n8015, n8016,
         n8017, n8020, n8021, n8022, n8023, n8024, n8025, n8026, n8027, n8028,
         n8029, n8030, n8031, n8032, n8033, n8034, n8035, n8037, n8039, n8041,
         n8042, n8043, n8044, n8045, n8046, n8047, n8048, n8049, n8050, n8051,
         n8052, n8053, n8054, \Ozkbx6[9] , \Ozkbx6[8] , \Ozkbx6[7] ,
         \Ozkbx6[6] , \Ozkbx6[5] , \Ozkbx6[4] , \Ozkbx6[3] , \Ozkbx6[33] ,
         \Ozkbx6[32] , \Ozkbx6[31] , \Ozkbx6[30] , \Ozkbx6[2] , \Ozkbx6[29] ,
         \Ozkbx6[28] , \Ozkbx6[27] , \Ozkbx6[26] , \Ozkbx6[25] , \Ozkbx6[24] ,
         \Ozkbx6[23] , \Ozkbx6[22] , \Ozkbx6[21] , \Ozkbx6[20] , \Ozkbx6[1] ,
         \Ozkbx6[19] , \Ozkbx6[18] , \Ozkbx6[17] , \Ozkbx6[16] , \Ozkbx6[15] ,
         \Ozkbx6[14] , \Ozkbx6[13] , \Ozkbx6[12] , \Ozkbx6[11] , \Ozkbx6[10] ,
         \eq_3147/A[0] , \eq_3147/A[1] , \eq_3147/A[2] , \eq_3147/A[3] ,
         \eq_3147/A[4] , \eq_3147/A[5] , \eq_3147/A[6] , \eq_3147/A[7] ,
         \eq_3147/A[8] , \eq_3147/A[9] , \eq_3147/A[10] , \eq_3147/A[11] ,
         \eq_3147/A[12] , \eq_3147/A[13] , \eq_3147/A[14] , \eq_3147/A[15] ,
         \eq_3147/A[16] , \eq_3147/A[17] , \eq_3147/A[18] , \eq_3147/A[19] ,
         \eq_3147/A[20] , \eq_3147/A[21] , \eq_3147/A[22] , \eq_3147/A[23] ,
         \eq_3147/A[24] , \eq_3147/A[25] , \eq_3147/A[26] , \sub_3151/A[0] ,
         \add_3107/carry[4] , \add_3107/carry[3] , \add_3107/B[1] , n221, n222,
         n225, n226, n228, n229, n230, n233, n234, n236, n237, n239, n242,
         n243, n244, n247, n249, n250, n253, n254, n265, n266, n267, n270,
         n272, n277, n279, n281, n283, n285, n287, n288, n290, n293, n298,
         n303, n308, n313, n316, n320, n323, n328, n332, n335, n339, n344,
         n349, n352, n356, n360, n365, n370, n371, n373, n376, n377, n380,
         n382, n384, n387, n389, n390, n391, n394, n396, n398, n399, n400,
         n403, n408, n420, n421, n422, n423, n424, n425, n430, n431, n432,
         n436, n437, n438, n439, n442, n448, n450, n451, n456, n458, n459,
         n460, n463, n464, n468, n470, n475, n476, n477, n479, n482, n485,
         n486, n491, n492, n502, n503, n505, n508, n516, n517, n521, n522,
         n523, n524, n526, n529, n536, n538, n540, n541, n547, n550, n561,
         n563, n564, n565, n567, n568, n569, n572, n575, n576, n577, n578,
         n581, n582, n599, n602, n615, n617, n623, n625, n627, n628, n629,
         n631, n632, n635, n640, n646, n650, n654, n659, n660, n661, n664,
         n667, n669, n670, n671, n672, n674, n678, n679, n680, n681, n682,
         n683, n684, n685, n686, n687, n688, n690, n691, n694, n695, n696,
         n697, n701, n704, n706, n709, n712, n713, n714, n722, n729, n731,
         n733, n734, n736, n737, n738, n739, n740, n743, n744, n747, n748,
         n749, n751, n753, n755, n757, n760, n761, n762, n764, n767, n768,
         n771, n772, n775, n776, n779, n780, n783, n784, n787, n788, n791,
         n794, n799, n800, n803, n807, n809, n815, n818, n824, n828, n830,
         n833, n836, n841, n847, n848, n850, n854, n855, n857, n863, n866,
         n872, n875, n878, n881, n883, n885, n890, n891, n892, n894, n897,
         n906, n908, n913, n917, n928, n931, n934, n941, n946, n950, n952,
         n955, n956, n961, n963, n964, n972, n974, n975, n976, n977, n986,
         n995, n1001, n1010, n1013, n1014, n1019, n1024, n1025, n1031, n1033,
         n1038, n1040, n1041, n1046, n1048, n1049, n1057, n1060, n1061, n1063,
         n1067, n1068, n1071, n1072, n1078, n1081, n1084, n1088, n1092, n1095,
         n1096, n1099, n1100, n1103, n1105, n1112, n1113, n1114, n1115, n1117,
         n1119, n1122, n1126, n1128, n1130, n1132, n1134, n1138, n1141, n1143,
         n1145, n1150, n1155, n1157, n1159, n1161, n1163, n1168, n1170, n1175,
         n1184, n1185, n1187, n1188, n1190, n1197, n1198, n1205, n1210, n1212,
         n1221, n1226, n1231, n1233, n1236, n1243, n1250, n1252, n1254, n1256,
         n1257, n1259, n1261, n1268, n1276, n1279, n1285, n1286, n1288, n1289,
         n1305, n1306, n1307, n1308, n1312, n1314, n1317, n1322, n1326, n1331,
         n1336, n1339, n1340, n1349, n1350, n1367, n1368, n1370, n1372, n1375,
         n1380, n1381, n1382, n1384, n1386, n1388, n1393, n1395, n1397, n1399,
         n1401, n1402, n1405, n1406, n1409, n1415, n1416, n1420, n1421, n1423,
         n1427, n1429, n1432, n1434, n1446, n1447, n1448, n1449, n1450, n1460,
         n1467, n1469, n1472, n1476, n1481, n1484, n1485, n1490, n1491, n1492,
         n1500, n1506, n1507, n1508, n1509, n1510, n1514, n1515, n1516, n1517,
         n1523, n1525, n1526, n1527, n1529, n1530, n1537, n1542, n1543, n1544,
         n1545, n1551, n1552, n1553, n1573, n1574, n1575, n1580, n1581, n1582,
         n1590, n1596, n1597, n1603, n1604, n1606, n1608, n1610, n1614, n1616,
         n1618, n1631, n1632, n1633, n1637, n1639, n1650, n1652, n1655, n1656,
         n1657, n1669, n1671, n1677, n1680, n1681, n1692, n1693, n1696, n1709,
         n1716, n1717, n1718, n1719, n1726, n1738, n1764, n1766, n1767, n1769,
         n1770, n1772, n1774, n1775, n1779, n1780, n1782, n1783, n1785, n1786,
         n1788, n1790, n1791, n1793, n1795, n1798, n1799, n1801, n1802, n1804,
         n1805, n1808, n1809, n1811, n1812, n1814, n1815, n1817, n1819, n1820,
         n1822, n1823, n1825, n1826, n1828, n1829, n1831, n1832, n1834, n1837,
         n1838, n1840, n1841, n1843, n1844, n1846, n1847, n1849, n1851, n1852,
         n1855, n1859, n1885, n1888, n1889, n1900, n1910, n1913, n1923, n1925,
         n1926, n1927, n1934, n1936, n1939, n1945, n1947, n1958, n1964, n1967,
         n1970, n1974, n1975, n1979, n1986, n1989, n1994, n1998, n1999, n2000,
         n2001, n2002, n2003, n2004, n2009, n2012, n2016, n2018, n2020, n2022,
         n2024, n2026, n2028, n2031, n2033, n2035, n2037, n2041, n2055, n2062,
         n2069, n2070, n2075, n2076, n2078, n2080, n2082, n2084, n2086, n2088,
         n2090, n2092, n2094, n2096, n2098, n2100, n2102, n2104, n2107, n2110,
         n2111, n2118, n2119, n2121, n2122, n2124, n2125, n2126, n2128, n2130,
         n2131, n2133, n2135, n2136, n2138, n2139, n2140, n2142, n2143, n2145,
         n2146, n2148, n2150, n2158, n2161, n2163, n2164, n2167, n2173, n2175,
         n2176, n2181, n2185, n2189, n2190, n2191, n2203, n2204, n2206, n2207,
         n2208, n2211, n2212, n2215, n2216, n2219, n2220, n2222, n2224, n2226,
         n2227, n2232, n2233, n2234, n2235, n2238, n2242, n2243, n2244, n2246,
         n2247, n2250, n2251, n2254, n2256, n2258, n2260, n2262, n2265, n2266,
         n2267, n2268, n2270, n2272, n2273, n2275, n2277, n2279, n2280, n2281,
         n2282, n2283, n2286, n2287, n2290, n2291, n2293, n2294, n2296, n2298,
         n2301, n2304, n2309, n2310, n2312, n2313, n2316, n2317, n2320, n2322,
         n2324, n2326, n2328, n2330, n2332, n2334, n2336, n2338, n2339, n2341,
         n2342, n2345, n2346, n2347, n2349, n2350, n2351, n2353, n2355, n2358,
         n2360, n2361, n2363, n2364, n2365, n2366, n2367, n2368, n2370, n2383,
         n2384, n2385, n2387, n2388, n2389, n2390, n2391, n2392, n2396, n2397,
         n2398, n2400, n2402, n2403, n2406, n2411, n2413, n2415, n2416, n2418,
         n2419, n2420, n2423, n2425, n2427, n2428, n2429, n2432, n2433, n2435,
         n2436, n2437, n2438, n2440, n2442, n2443, n2444, n2445, n2447, n2449,
         n2451, n2456, n2457, n2458, n2459, n2460, n2462, n2464, n2466, n2468,
         n2470, n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2481, n2485,
         n2486, n2490, n2500, n2502, n2506, n2507, n2508, n2509, n2510, n2511,
         n2512, n2513, n2514, n2515, n2516, n2517, n2519, n2522, n2524, n2527,
         n2528, n2529, n2530, n2533, n2535, n2537, n2538, n2539, n2541, n2543,
         n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2553, n2569,
         n2572, n2575, n2582, n2584, n2590, n2591, n2594, n2595, n2596, n2597,
         n2598, n2599, n2601, n2603, n2605, n2606, n2607, n2608, n2609, n2610,
         n2614, n2615, n2616, n2617, n2632, n2644, n2645, n2646, n2647, n2648,
         n2649, n2650, n2651, n2652, n2653, n2654, n2655, n2656, n2657, n2660,
         n2663, n2664, n2666, n2667, n2670, n2671, n2674, n2675, n2676, n2678,
         n2679, n2682, n2684, n2686, n2688, n2689, n2690, n2691, n2692, n2693,
         n2694, n2696, n2697, n2698, n2699, n2700, n2702, n2703, n2708, n2710,
         n2711, n2712, n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720,
         n2721, n2722, n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730,
         n2731, n2732, n2745, n2757, n2758, n2759, n2770, n2776, n2777, n2778,
         n2779, n2781, n2782, n2783, n2786, n2787, n2788, n2789, n2790, n2792,
         n2793, n2794, n2797, n2799, n2809, n2811, n2812, n2813, n2814, n2815,
         n2816, n2817, n2818, n2820, n2822, n2825, n2826, n2827, n2828, n2832,
         n2833, n2834, n2835, n2836, n2840, n2852, n2855, n2856, n2857, n2858,
         n2865, n2866, n2869, n2882, n2883, n2884, n2885, n2886, n2897, n2901,
         n2906, n2937, n2938, n2942, n2943, n2944, n2949, n2955, n2960, n2961,
         n2963, n2964, n2965, n2967, n2969, n2972, n2973, n2974, n2975, n2976,
         n2977, n2978, n2983, n2985, n2986, n2987, n2988, n2989, n2992, n2998,
         n3002, n3004, n3006, n3007, n3008, n3009, n3010, n3012, n3013, n3014,
         n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3024, n3030, n3031,
         n3032, n3033, n3036, n3037, n3039, n3040, n3041, n3042, n3045, n3047,
         n3048, n3056, n3060, n3061, n3062, n3063, n3064, n3065, n3066, n3067,
         n3068, n3072, n3078, n3080, n3081, n3082, n3083, n3084, n3085, n3086,
         n3087, n3089, n3091, n3096, n3101, n3102, n3103, n3104, n3105, n3106,
         n3107, n3108, n3109, n3110, n3111, n3112, n3113, n3114, n3115, n3116,
         n3117, n3118, n3119, n3120, n3121, n3122, n3123, n3124, n3125, n3126,
         n3127, n3128, n3129, n3130, n3131, n3132, n3133, n3135, n3136, n3137,
         n3138, n3139, n3140, n3141, n3142, n3143, n3144, n3145, n3146, n3147,
         n3149, n3150, n3151, n3152, n3153, n3154, n3156, n3158, n3180, n3190,
         n3191, n3192, n3195, n3197, n3200, n3201, n3202, n3203, n3204, n3205,
         n3208, n3212, n3215, n3216, n3219, n3223, n3225, n3226, n3233, n3242,
         n3258, n3259, n3268, n3272, n3274, n3276, n3278, n3279, n3280, n3287,
         n3290, n3292, n3293, n3296, n3300, n3310, n3324, n3329, n3335, n3337,
         n3341, n3343, n3347, n3351, n3358, n3369, n3388, n3389, n3397, n3404,
         n3405, n3419, n3439, n3441, n3443, n3444, n3446, n3450, n3451, n3453,
         n3454, n3456, n3460, n3467, n3468, n3470, n3471, n3472, n3473, n3474,
         n3475, n3476, n3478, n3479, n3480, n3481, n3482, n3483, n3484, n3486,
         n3488, n3503, n3505, n3520, n3532, n3533, n3534, n3535, n3538, n3540,
         n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3554,
         n3556, n3566, n3571, n3576, n3581, n3583, n3586, n3587, n3588, n3591,
         n3592, n3593, n3596, n3598, n3601, n3602, n3604, n3607, n3608, n3611,
         n3614, n3617, n3618, n3620, n3623, n3625, n3628, n3630, n3631, n3634,
         n3635, n3638, n3640, n3643, n3645, n3648, n3650, n3653, n3654, n3656,
         n3659, n3661, n3664, n3666, n3668, n3669, n3672, n3673, n3676, n3682,
         n3684, n3686, n3690, n3697, n3698, n3699, n3701, n3702, n3703, n3705,
         n3706, n3707, n3709, n3710, n3712, n3713, n3714, n3725, n3726, n3727,
         n3730, n3732, n3733, n3737, n3740, n3744, n3746, n3749, n3757, n3760,
         n3761, n3762, n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3773,
         n3774, n3775, n3780, n3781, n3783, n3784, n3785, n3786, n3787, n3788,
         n3790, n3800, n3803, n3804, n3805, n3830, n3831, n3832, n3833, n3835,
         n3836, n3837, n3838, n3840, n3841, n3843, n3845, n3846, n3849, n3851,
         n3855, n3858, n3860, n3863, n3864, n3865, n3866, n3867, n3868, n3869,
         n3870, n3871, n3875, n3877, n3879, n3880, n3882, n3883, n3884, n3886,
         n3890, n3894, n3895, n3899, n3904, n3911, n3913, n3915, n3922, n3924,
         n3925, n3926, n3928, n3930, n3931, n3934, n3935, n3936, n3937, n3938,
         n3939, n3940, n3946, n3947, n3948, n3951, n3952, n3954, n3955, n3957,
         n3959, n3960, n3961, n3967, n3968, n3971, n3972, n3973, n3975, n3977,
         n3978, n3979, n3980, n3981, n3983, n3984, n3985, n3986, n3987, n3988,
         n3989, n3990, n4001, n4002, n4003, n4004, n4005, n4006, n4007, n4008,
         n4009, n4010, n4011, n4015, n4016, n4017, n4018, n4022, n4024, n4027,
         n4028, n4029, n4032, n4033, n4034, n4035, n4036, n4038, n4040, n4041,
         n4042, n4044, n4046, n4048, n4049, n4052, n4053, n4054, n4055, n4061,
         n4063, n4066, n4070, n4072, n4078, n4086, n4109, n4110, n4111, n4112,
         n4115, n4116, n4117, n4118, n4119, n4123, n4126, n4134, n4135, n4136,
         n4138, n4139, n4140, n4141, n4142, n4144, n4145, n4146, n4149, n4151,
         n4152, n4157, n4158, n4160, n4161, n4163, n4164, n4167, n4170, n4172,
         n4178, n4179, n4180, n4181, n4182, n4184, n4185, n4186, n4187, n4188,
         n4189, n4190, n4193, n4194, n4195, n4196, n4199, n4202, n4203, n4204,
         n4205, n4215, n4222, n4229, n4232, n4237, n4240, n4244, n4245, n4246,
         n4250, n4263, n4265, n4271, n4272, n4273, n4275, n4278, n4280, n4281,
         n4282, n4285, n4293, n4297, n4301, n4306, n4324, n4329, n4330, n4333,
         n4335, n4336, n4341, n4348, n4351, n4352, n4364, n4376, n4378, n4379,
         n4394, n4395, n4402, n4405, n4406, n4408, n4409, n4410, n4420, n4431,
         n4432, n4433, n4434, n4435, n4436, n4437, n4441, n4442, n4453, n4454,
         n4459, n4460, n4465, n4466, n4467, n4468, n4470, n4473, n4474, n4478,
         n4482, n4487, n4491, n4506, n4507, n4512, n4521, n4535, n4545, n4546,
         n4548, n4554, n4555, n4564, n4566, n4572, n4579, n4587, n4588, n4591,
         n4598, n4602, n4608, n4610, n4611, n4616, n4628, n4631, n4633, n4635,
         n4637, n4642, n4650, n4651, n4658, n4667, n4668, n4669, n4670, n4672,
         n4673, n4674, n4685, n4687, n4688, n4693, n4694, n4695, n4699, n4700,
         n4701, n4702, n4703, n4704, n4707, n4708, n4713, n4720, n4721, n4724,
         n4725, n4732, n4738, n4749, n4753, n4756, n4761, n4764, n4765, n4766,
         n4772, n4773, n4774, n4776, n4777, n4782, n4783, n4787, n4795, n4797,
         n4799, n4801, n4802, n4805, n4806, n4807, n4810, n4811, n4816, n4818,
         n4826, n4839, n4841, n4855, n4908, n4910, n4932, n4940, n4978, n4987,
         n4993, n5002, n5037, n5042, n5047, n5063, n5065, n5070, n5074, n5088,
         n5105, n5111, n5112, n5126, n5128, n5129, n5134, n5148, n5154, n5175,
         n5180, n5192, n5193, n5197, n5198, n5209, n5210, n5216, n5225, n5236,
         n5237, n5256, n5257, n5258, n5266, n5270, n5272, n5273, n5277, n5278,
         n5282, n5284, n5291, n5293, n5294, n5299, n5302, n5304, n5307, n5312,
         n5313, n5317, n5319, n5326, n5333, n5334, n5348, n5352, n5366, n5369,
         n5370, n5372, n5386, n5394, n5403, n5409, n5410, n5411, n5419, n5427,
         n5428, n5433, n5449, n5451, n5460, n5461, n5462, n5463, n5464, n5465,
         n5467, n5468, n5470, n5484, n5485, n5493, n5506, n5507, n5520, n5521,
         n5522, n5523, n5526, n5532, n5534, n5540, n5541, n5551, n5552, n5555,
         n5556, n5562, n5579, n5580, n5584, n5598, n5606, n5624, n5642, n5654,
         n5662, n5663, n5669, n5673, n5676, n5682, n5683, n5684, n5689, n5709,
         n5710, n5711, n5718, n5725, n5726, n5729, n5730, n5736, n5739, n5752,
         n5789, n5793, n5794, n5799, n5802, n5810, n5811, n5814, n5820, n5822,
         n5825, n5829, n5832, n5834, n5839, n5846, n5848, n5849, n5851, n5859,
         n5860, n5865, n5872, n5873, n5875, n5876, n5877, n5886, n5887, n5891,
         n5892, n5894, n5895, n5897, n5898, n5899, n5901, n5905, n5914, n5915,
         n5924, n5928, n5935, n5937, n5938, n5939, n5940, n5941, n5948, n5955,
         n5956, n5959, n5960, n5961, n5963, n5964, n5976, n5989, n5990, n5993,
         n6039, n6080, n6104, n6105, n6119, n6120, n6121, n6122, n6124, n6128,
         n6129, n6136, n6138, n6142, n6144, n6146, n6148, n6150, n6151, n6152,
         n6153, n6156, n6167, n6168, n6175, n6176, n6177, n6178, n6183, n6188,
         n6202, n6207, n6210, n6212, n6218, n6219, n6220, n6221, n6225, n6229,
         n6234, n6239, n6241, n6242, n6249, n6253, n6257, n6260, n6264, n6266,
         n6267, n6271, n6280, n6281, n6289, n6290, n6291, n6292, n6294, n6306,
         n6313, n6317, n6324, n6328, n6329, n6330, n6331, n6341, n6349, n6351,
         n6352, n6355, n6365, n6372, n6377, n6378, n6380, n6386, n6387, n6394,
         n6395, n6399, n6425, n6452, n6478, n6479, n6480, n6484, n6486, n6487,
         n6504, n6518, n6524, n6526, n6537, n6560, n6564, n6570, n6571, n6574,
         n6577, n6583, n6585, n6586, n6588, n6590, n6595, n6599, n6600, n6603,
         n6605, n6607, n6626, n6628, n6636, n6638, n6639, n6642, n6646, n6650,
         n6657, n6663, n6668, n6669, n6674, n6677, n6678, n6686, n6771, n6810,
         n6819, n6826, n6835, n6863, n6871, n6886, n6899, n6918, n7261, n7307,
         n7341, n7342, n7370, n7372, n7376, n7377, n7512, n7571, n7573, n7575,
         n7577, n7578, n7579, n7580, n7600, n7603, n7643, n7644, n7668, n7695,
         n7704, n7745, n7748, n7751, n7754, n7757, n7760, n7763, n7766, n7769,
         n7772, n7775, n7778, n7781, n7784, n7787, n7790, n7793, n7797, n7800,
         n7802, n7806, n7809, n7811, n7815, n7818, n7821, n7824, n7922, n8008,
         n8018, n8019, n8036, n8038, n8040, n8055, n8056, n8057, n8058, n8059,
         n8060, n8061, n8062, n8063, n8064, n8065, n8066, n8067, n8068, n8069,
         n8070, n8071, n8072, n8073, n8074, n8075, n8076, n8077, n8078, n8079,
         n8080, n8081, n8082, n8083, n8084, n8085, n8086, n8087, n8088, n8089,
         n8090, n8091, n8092, n8093, n8094, n8095, n8096, n8097, n8098, n8099,
         n8100, n8101, n8102, n8103, n8104, n8105, n8106, n8107, n8108, n8109,
         n8110, n8111, n8112, n8113, n8114, n8115, n8116, n8117, n8118, n8119,
         n8120, n8121, n8122, n8123, n8124, n8125, n8126, n8127, n8128, n8129,
         n8130, n8131, n8132, n8133, n8134, n8135, n8136, n8137, n8138, n8139,
         n8140, n8141, n8142, n8143, n8144, n8145, n8146, n8147, n8148, n8149,
         n8150, n8151, n8152, n8153, n8154, n8155, n8156, n8157, n8158, n8159,
         n8160, n8161, n8162, n8163, n8164, n8165, n8166, n8167, n8168, n8169,
         n8170, n8171, n8172, n8173, n8174, n8175, n8176, n8177, n8178, n8179,
         n8180, n8181, n8182, n8183, n8184, n8185, n8186, n8187, n8188, n8189,
         n8190, n8191, n8192, n8193, n8194, n8195, n8196, n8197, n8198, n8199,
         n8200, n8201, n8202, n8203, n8204, n8205, n8206, n8207, n8208, n8209,
         n8210, n8211, n8212, n8213, n8214, n8215, n8216, n8217, n8218, n8219,
         n8220, n8221, n8222, n8223, n8224, n8225, n8226, n8227, n8228, n8229,
         n8230, n8231, n8232, n8233, n8234, n8235, n8236, n8237, n8238, n8239,
         n8240, n8241, n8242, n8243, n8244, n8245, n8246, n8247, n8248, n8249,
         n8250, n8251, n8252, n8253, n8254, n8255, n8256, n8257, n8258, n8259,
         n8260, n8261, n8262, n8263, n8264, n8265, n8266, n8267, n8268, n8269,
         n8270, n8271, n8272, n8273, n8274, n8275, n8276, n8277, n8278, n8279,
         n8280, n8281, n8282, n8283, n8284, n8285, n8286, n8287, n8288, n8289,
         n8290, n8291, n8292, n8293, n8294, n8295, n8296, n8297, n8298, n8299,
         n8300, n8301, n8302, n8303, n8304, n8305, n8306, n8307, n8308, n8309,
         n8310, n8311, n8312, n8313, n8314, n8315, n8316, n8317, n8318, n8319,
         n8320, n8321, n8322, n8323, n8324, n8325, n8326, n8327, n8328, n8329,
         n8330, n8331, n8332, n8333, n8334, n8335, n8336, n8337, n8338, n8339,
         n8340, n8341, n8342, n8343, n8344, n8345, n8346, n8347, n8348, n8349,
         n8350, n8351, n8352, n8353, n8354, n8355, n8356, n8357, n8358, n8359,
         n8360, n8361;
  wire   [23:0] Tzfpw6;
  wire   [31:4] Jshpw6;
  wire   [3:0] Tnhpw6;
  wire   [31:2] K7hpw6;
  wire   [31:2] E1hpw6;
  wire   [28:2] Gtgpw6;
  wire   [28:2] Togpw6;
  wire   [28:2] Gqgpw6;
  wire   [28:2] Trgpw6;
  wire   [10:1] Vrkbx6;
  wire   [30:0] Ntkbx6;
  wire   [30:0] Nvkbx6;
  wire   [23:0] L6gpw6;
  wire   [7:0] Vnfpw6;
  wire   [8:1] Xlfpw6;
  wire   [30:0] Zsfpw6;
  wire   [30:2] N5fpw6;
  wire   [31:0] Mifpw6;
  wire   [31:0] Tgfpw6;
  wire   [31:0] Affpw6;
  wire   [33:1] Nxkbx6;
  wire   [30:23] Qbfpw6;
  wire   [31:0] Idfpw6;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15, 
        SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17, 
        SYNOPSYS_UNCONNECTED__18, SYNOPSYS_UNCONNECTED__19, 
        SYNOPSYS_UNCONNECTED__20, SYNOPSYS_UNCONNECTED__21, 
        SYNOPSYS_UNCONNECTED__22, SYNOPSYS_UNCONNECTED__23, 
        SYNOPSYS_UNCONNECTED__24, SYNOPSYS_UNCONNECTED__25, 
        SYNOPSYS_UNCONNECTED__26, SYNOPSYS_UNCONNECTED__27, 
        SYNOPSYS_UNCONNECTED__28, SYNOPSYS_UNCONNECTED__29, 
        SYNOPSYS_UNCONNECTED__30, SYNOPSYS_UNCONNECTED__31, 
        SYNOPSYS_UNCONNECTED__32, SYNOPSYS_UNCONNECTED__33, 
        SYNOPSYS_UNCONNECTED__34;
  assign N427 = RSTBYPASS;
  assign HPROT[0] = HPROT_0;
  assign N701 = HREADY;

  DFFR_X1 Evhpw6_reg ( .D(1'b1), .CK(SWCLKTCK), .RN(PORESETn), .Q(Qmdhu6) );
  DFFR_X1 Hwhpw6_reg ( .D(Qmdhu6), .CK(SWCLKTCK), .RN(PORESETn), .Q(Pndhu6) );
  DFFR_X1 Kxhpw6_reg ( .D(Pndhu6), .CK(SWCLKTCK), .RN(PORESETn), .Q(Oodhu6) );
  DFFR_X1 Nyhpw6_reg ( .D(CDBGPWRUPACK), .CK(SWCLKTCK), .RN(Fmdhu6), .Q(O5ohu6) );
  DFFR_X1 Isjpw6_reg ( .D(E5xhu6), .CK(DCLK), .RN(DBGRESETn), .Q(n6683), .QN(
        n3008) );
  DFF_X1 Hg7ax6_reg ( .D(n7912), .CK(DCLK), .Q(n6644) );
  DFF_X1 Nrkpw6_reg ( .D(n7903), .CK(DCLK), .Q(n6654) );
  DFF_X1 E6iax6_reg ( .D(n7870), .CK(SCLK), .QN(n3620) );
  DFFR_X1 Mk3bx6_reg ( .D(A4phu6), .CK(SCLK), .RN(HRESETn), .Q(n6576), .QN(
        n3645) );
  DFF_X1 V53qw6_reg ( .D(n7910), .CK(DCLK), .Q(n6648), .QN(n3883) );
  DFF_X1 Pifax6_reg ( .D(Avxhu6), .CK(SWCLKTCK), .Q(n6596), .QN(n4044) );
  DFF_X1 Xu2qw6_reg ( .D(n7911), .CK(DCLK), .QN(n4048) );
  DFFR_X1 Qufax6_reg ( .D(Dtnhu6), .CK(SWCLKTCK), .RN(n956), .Q(S3ohu6) );
  DFFR_X1 Utqpw6_reg ( .D(n7830), .CK(SWCLKTCK), .RN(Fmdhu6), .Q(G2ohu6), .QN(
        n6675) );
  DFFR_X1 Xvqpw6_reg ( .D(G2ohu6), .CK(DCLK), .RN(DBGRESETn), .Q(Q7ohu6) );
  DFFR_X1 Xkqpw6_reg ( .D(Ytxhu6), .CK(SWCLKTCK), .RN(Fmdhu6), .Q(CDBGPWRUPREQ), .QN(n7349) );
  DFFR_X1 Rekbx6_reg ( .D(n7880), .CK(HCLK), .RN(HRESETn), .Q(SYSRESETREQ), 
        .QN(n6661) );
  DFFS_X1 K7vpw6_reg ( .D(n8010), .CK(DCLK), .SN(DBGRESETn), .Q(DBGRESTARTED)
         );
  DFFR_X1 Bciax6_reg ( .D(n7871), .CK(SCLK), .RN(HRESETn), .QN(n5236) );
  DFF_X1 Nckbx6_reg ( .D(n7908), .CK(DCLK), .QN(n8284) );
  DFFR_X1 Dqkbx6_reg ( .D(n7841), .CK(SWCLKTCK), .RN(Fmdhu6), .Q(SWDOEN), .QN(
        n6670) );
  OAI33_X1 U40 ( .A1(n2281), .A2(Nxkbx6[32]), .A3(n2537), .B1(n1544), .B2(
        Idfpw6[31]), .B3(D5epw6), .ZN(n104) );
  OAI33_X1 U62 ( .A1(n136), .A2(n137), .A3(n138), .B1(n139), .B2(n140), .B3(
        n141), .ZN(n135) );
  OAI33_X1 U79 ( .A1(HADDR[11]), .A2(n164), .A3(HADDR[8]), .B1(n167), .B2(
        n1772), .B3(n328), .ZN(n165) );
  OAI33_X1 U102 ( .A1(n394), .A2(n7468), .A3(n7469), .B1(n390), .B2(n7474), 
        .B3(n7475), .ZN(n189) );
  OAI33_X1 U103 ( .A1(n396), .A2(n7472), .A3(n7473), .B1(n391), .B2(n7470), 
        .B3(n7471), .ZN(n188) );
  OAI33_X1 U110 ( .A1(n394), .A2(n7469), .A3(n7483), .B1(n390), .B2(n7475), 
        .B3(n7484), .ZN(n205) );
  OAI33_X1 U113 ( .A1(n396), .A2(n7473), .A3(n7485), .B1(n391), .B2(n7471), 
        .B3(n7486), .ZN(n204) );
  OAI33_X1 U580 ( .A1(Jshpw6[8]), .A2(n951), .A3(n8172), .B1(n953), .B2(n947), 
        .B3(n954), .ZN(n949) );
  OAI33_X1 U881 ( .A1(n1283), .A2(n4405), .A3(n4333), .B1(n3915), .B2(n3478), 
        .B3(n1309), .ZN(n998) );
  OAI33_X1 U1058 ( .A1(n3705), .A2(n3123), .A3(n2529), .B1(n2266), .B2(n475), 
        .B3(n1939), .ZN(n1445) );
  OAI33_X1 U1085 ( .A1(n2243), .A2(n878), .A3(n1958), .B1(n1936), .B2(n524), 
        .B3(n7516), .ZN(n1513) );
  OAI33_X1 U1148 ( .A1(n3709), .A2(n7497), .A3(n4608), .B1(n2243), .B2(n476), 
        .B3(n1958), .ZN(n1648) );
  OAI33_X1 U1160 ( .A1(n2607), .A2(n3550), .A3(n3714), .B1(n1670), .B2(n2697), 
        .B3(n4186), .ZN(n1667) );
  OAI33_X1 U1184 ( .A1(n4195), .A2(n2524), .A3(n4246), .B1(n2603), .B2(n3556), 
        .B3(n3714), .ZN(n1715) );
  OAI33_X1 U1189 ( .A1(n508), .A2(n1721), .A3(n516), .B1(n1722), .B2(n4610), 
        .B3(n1572), .ZN(n1713) );
  OAI33_X1 U1201 ( .A1(n3835), .A2(n7373), .A3(n2572), .B1(n1739), .B2(n270), 
        .B3(n2277), .ZN(n1736) );
  OAI33_X1 U1344 ( .A1(n1891), .A2(n7352), .A3(n1890), .B1(n1892), .B2(n7702), 
        .B3(n1886), .ZN(n8003) );
  OAI33_X1 U1377 ( .A1(n3746), .A2(n266), .A3(n3803), .B1(n5002), .B2(n1946), 
        .B3(n1934), .ZN(n1944) );
  OAI33_X1 U2332 ( .A1(n3803), .A2(n536), .A3(n2572), .B1(n1572), .B2(n2561), 
        .B3(n523), .ZN(n2559) );
  OAI33_X1 U2482 ( .A1(n3142), .A2(n2704), .A3(n4024), .B1(n2705), .B2(n548), 
        .B3(n3208), .ZN(n2184) );
  OAI33_X1 U2525 ( .A1(n516), .A2(n2737), .A3(n4693), .B1(n2738), .B2(n4195), 
        .B3(n2594), .ZN(n2736) );
  OAI33_X1 U2537 ( .A1(n2756), .A2(n270), .A3(n2124), .B1(n4199), .B2(n3713), 
        .B3(n2524), .ZN(n2748) );
  OAI33_X1 U2639 ( .A1(n3628), .A2(n2698), .A3(n2262), .B1(n2529), .B2(n267), 
        .B3(n265), .ZN(n2847) );
  OAI33_X1 U2655 ( .A1(n522), .A2(n7359), .A3(n4688), .B1(n2864), .B2(n7259), 
        .B3(n7325), .ZN(n2863) );
  XOR2_X1 U2704 ( .A(n2925), .B(n4572), .Z(n65) );
  XOR2_X1 U2706 ( .A(n2930), .B(n2931), .Z(n2929) );
  OAI33_X1 U2711 ( .A1(n4245), .A2(n524), .A3(n4237), .B1(n4196), .B2(n7374), 
        .B3(n3804), .ZN(n2936) );
  XOR2_X1 U2769 ( .A(n2504), .B(n2505), .Z(n2503) );
  OAI33_X1 U2952 ( .A1(n4608), .A2(n7373), .A3(n522), .B1(n2524), .B2(n517), 
        .B3(n4237), .ZN(n3171) );
  OAI33_X1 U3014 ( .A1(n4188), .A2(n7514), .A3(n2273), .B1(n444), .B2(n7399), 
        .B3(n3628), .ZN(n2846) );
  XOR2_X1 U3037 ( .A(n7329), .B(n3241), .Z(n3247) );
  OAI33_X1 U3124 ( .A1(n3308), .A2(n3309), .A3(n3072), .B1(n3311), .B2(n3312), 
        .B3(n3313), .ZN(n3307) );
  OAI33_X1 U3126 ( .A1(n3317), .A2(n3318), .A3(n3319), .B1(n3320), .B2(n3321), 
        .B3(n3322), .ZN(n3316) );
  OAI33_X1 U3145 ( .A1(n3080), .A2(n3309), .A3(n3078), .B1(n3370), .B2(n3371), 
        .B3(n3372), .ZN(n3350) );
  OAI33_X1 U3147 ( .A1(n3376), .A2(n3366), .A3(n3365), .B1(n3377), .B2(n3378), 
        .B3(n3379), .ZN(n3375) );
  OAI33_X1 U3235 ( .A1(n4265), .A2(n2572), .A3(n4650), .B1(n3705), .B2(n3123), 
        .B3(n2608), .ZN(n3501) );
  OAI33_X1 U3253 ( .A1(n4232), .A2(n2572), .A3(n516), .B1(n5037), .B2(n7381), 
        .B3(n2256), .ZN(n3519) );
  OAI33_X1 U3256 ( .A1(n3625), .A2(n1595), .A3(n4187), .B1(n4188), .B2(n7381), 
        .B3(n4572), .ZN(n3525) );
  OAI33_X1 U3295 ( .A1(n3838), .A2(n265), .A3(n2524), .B1(n3232), .B2(n878), 
        .B3(n4263), .ZN(n3563) );
  OAI33_X1 U3482 ( .A1(n3722), .A2(n7374), .A3(n3723), .B1(n3724), .B2(n4265), 
        .B3(n4591), .ZN(n3719) );
  OAI33_X1 U3697 ( .A1(n950), .A2(n7489), .A3(n2395), .B1(n3896), .B2(n669), 
        .B3(n3897), .ZN(n8379) );
  XOR2_X1 U3735 ( .A(n3908), .B(n1981), .Z(n3907) );
  XOR2_X1 U3905 ( .A(n754), .B(n7494), .Z(n4000) );
  XOR2_X1 U3906 ( .A(n756), .B(n7495), .Z(n3999) );
  OAI33_X1 U4032 ( .A1(n4598), .A2(n4693), .A3(n4263), .B1(n4688), .B2(n4081), 
        .B3(n4512), .ZN(n4076) );
  XOR2_X1 U4136 ( .A(n2545), .B(n4165), .Z(n4162) );
  OAI33_X1 U4181 ( .A1(n1934), .A2(n7381), .A3(n4212), .B1(n2572), .B2(n4213), 
        .B3(n4693), .ZN(n4211) );
  OAI33_X1 U4192 ( .A1(n1958), .A2(n878), .A3(n4217), .B1(n1925), .B2(n4218), 
        .B3(n4507), .ZN(n4210) );
  OAI33_X1 U4197 ( .A1(n4220), .A2(n1947), .A3(n4987), .B1(n4221), .B2(n2260), 
        .B3(n1936), .ZN(n4209) );
  OAI33_X1 U4229 ( .A1(n2509), .A2(n878), .A3(n3737), .B1(n4230), .B2(n2524), 
        .B3(n3727), .ZN(n4228) );
  XOR2_X1 U4259 ( .A(n4257), .B(n4258), .Z(n4255) );
  OAI33_X1 U4391 ( .A1(n2275), .A2(n4369), .A3(n4188), .B1(n2694), .B2(n7510), 
        .B3(n4370), .ZN(n4368) );
  XOR2_X1 U4451 ( .A(n4392), .B(n4258), .Z(n4386) );
  XOR2_X1 U4481 ( .A(n2545), .B(n4423), .Z(n4422) );
  XOR2_X1 U4536 ( .A(n2545), .B(n4481), .Z(n4480) );
  XOR2_X1 U4590 ( .A(n2545), .B(n4518), .Z(n4511) );
  XOR2_X1 U4662 ( .A(n2545), .B(n4601), .Z(n4600) );
  XOR2_X1 U4697 ( .A(n4624), .B(n4258), .Z(n4617) );
  XOR2_X1 U4779 ( .A(n2545), .B(n4686), .Z(n4660) );
  XOR2_X1 U4829 ( .A(n4742), .B(n4258), .Z(n4741) );
  XOR2_X1 U4930 ( .A(n2545), .B(n4798), .Z(G3epw6) );
  XOR2_X1 U4971 ( .A(n4831), .B(n4258), .Z(n4824) );
  OAI33_X1 U5374 ( .A1(n1925), .A2(n470), .A3(n4572), .B1(n3757), .B2(n5036), 
        .B3(n449), .ZN(n5035) );
  XOR2_X1 U5470 ( .A(n2545), .B(n5073), .Z(n5072) );
  XOR2_X1 U5514 ( .A(n5099), .B(n4258), .Z(n5094) );
  XOR2_X1 U5623 ( .A(n2545), .B(n5157), .Z(n5156) );
  OAI33_X1 U5741 ( .A1(n4265), .A2(n4512), .A3(n4611), .B1(n4687), .B2(n1539), 
        .B3(n5211), .ZN(n5208) );
  OAI33_X1 U5755 ( .A1(n3828), .A2(n265), .A3(n3858), .B1(n4195), .B2(n7373), 
        .B3(n3804), .ZN(n5212) );
  OAI33_X1 U5829 ( .A1(n3729), .A2(n3113), .A3(n485), .B1(n1524), .B2(n4243), 
        .B3(n2572), .ZN(n5252) );
  OAI33_X1 U6111 ( .A1(n4790), .A2(n5314), .A3(n5320), .B1(n5458), .B2(n5459), 
        .B3(n2783), .ZN(n5455) );
  XOR2_X1 U6307 ( .A(n2545), .B(n5609), .Z(n5608) );
  OAI33_X1 U6348 ( .A1(n3831), .A2(n516), .A3(n3730), .B1(n3055), .B2(n479), 
        .B3(n522), .ZN(n5628) );
  OAI33_X1 U6410 ( .A1(n2607), .A2(n7373), .A3(n4507), .B1(n4608), .B2(n878), 
        .B3(n3714), .ZN(n5636) );
  OAI33_X1 U6571 ( .A1(n4642), .A2(n4237), .A3(n522), .B1(n2470), .B2(n7284), 
        .B3(n7343), .ZN(n5732) );
  OAI33_X1 U6582 ( .A1(n3804), .A2(n265), .A3(n272), .B1(n2572), .B2(n7282), 
        .B3(n7374), .ZN(n5735) );
  XOR2_X1 U6586 ( .A(n5740), .B(n4258), .Z(n5715) );
  OAI33_X1 U6590 ( .A1(n3730), .A2(n517), .A3(n7373), .B1(n4196), .B2(n7283), 
        .B3(n524), .ZN(n5744) );
  OAI33_X1 U6605 ( .A1(n2591), .A2(n4237), .A3(n3764), .B1(n3788), .B2(n228), 
        .B3(n4199), .ZN(n5748) );
  OAI33_X1 U7284 ( .A1(n3015), .A2(n6114), .A3(n6115), .B1(n6116), .B2(n5316), 
        .B3(n6117), .ZN(n6113) );
  OAI33_X1 U7294 ( .A1(n6141), .A2(n3036), .A3(n2792), .B1(n6143), .B2(n3120), 
        .B3(n6145), .ZN(n6140) );
  OAI33_X1 U7434 ( .A1(n6258), .A2(n6194), .A3(n6259), .B1(n3292), .B2(n3866), 
        .B3(n3869), .ZN(n6193) );
  OAI33_X1 U8112 ( .A1(n3723), .A2(n517), .A3(n3764), .B1(n3855), .B2(n7282), 
        .B3(n4651), .ZN(n6551) );
  OAI33_X1 U8143 ( .A1(n4232), .A2(n479), .A3(n3804), .B1(n4246), .B2(n272), 
        .B3(n3858), .ZN(n6561) );
  NOR3_X2 U275 ( .A1(n2130), .A2(n1851), .A3(n258), .ZN(n182) );
  OAI21_X2 U2464 ( .B1(n4158), .B2(n4111), .A(HMASTER), .ZN(SPECHTRANS) );
  NOR2_X2 U2467 ( .A1(n7560), .A2(n5237), .ZN(SLEEPDEEP) );
  OAI21_X2 U3701 ( .B1(HADDR[31]), .B2(n1553), .A(HPROT[2]), .ZN(HPROT[3]) );
  OAI21_X2 U3788 ( .B1(n952), .B2(n3920), .A(n3921), .ZN(HADDR[0]) );
  AOI21_X2 U3870 ( .B1(SLEEPHOLDACKn), .B2(n5237), .A(CDBGPWRUPACK), .ZN(
        GATEHCLK) );
  NOR2_X2 U4420 ( .A1(n7519), .A2(n33), .ZN(CODEHINTDE[1]) );
  NOR2_X2 U4421 ( .A1(n4670), .A2(n33), .ZN(CODEHINTDE[0]) );
  NOR3_X2 U5210 ( .A1(n4047), .A2(n3897), .A3(n3878), .ZN(n4850) );
  NOR2_X2 U6496 ( .A1(n632), .A2(n4253), .ZN(n4446) );
  NOR3_X2 U6585 ( .A1(n4244), .A2(n7279), .A3(n4190), .ZN(n4253) );
  NOR3_X2 U6990 ( .A1(n3913), .A2(n7448), .A3(n3470), .ZN(n844) );
  NOR2_X2 U7872 ( .A1(n5387), .A2(n3327), .ZN(n4717) );
  AOI211_X2 U7877 ( .C1(n524), .C2(n433), .A(n479), .B(n6473), .ZN(n5786) );
  NOR2_X2 U7918 ( .A1(n5387), .A2(n3105), .ZN(n4690) );
  OAI21_X2 U7920 ( .B1(n254), .B2(n6481), .A(n6482), .ZN(n3327) );
  NOR2_X2 U8118 ( .A1(n7373), .A2(n521), .ZN(n493) );
  cortexm0ds_logic_DW01_inc_0 add_3152 ( .A(vis_pc_o), .SUM(Zsfpw6) );
  cortexm0ds_logic_DW01_dec_1 sub_3150 ( .A(Tzfpw6), .SUM(L6gpw6) );
  cortexm0ds_logic_DW01_cmp6_4 eq_3124 ( .A({M9ohu6, Uilhu6, Nhlhu6, Gglhu6, 
        Zelhu6, Sdlhu6, Lclhu6, Eblhu6, W9lhu6, O8lhu6, G7lhu6, Y5lhu6, Q4lhu6, 
        I3lhu6, A2lhu6, S0lhu6, Kzkhu6, Cykhu6, Uwkhu6, Mvkhu6, Eukhu6, Wskhu6, 
        Orkhu6, Gqkhu6, Yokhu6, Qnkhu6, Imkhu6, Alkhu6, Sjkhu6, Kikhu6, Chkhu6, 
        Ufkhu6}), .B({K7hpw6, Avmhu6, Ttmhu6}), .TC(1'b0), .EQ(N439) );
  cortexm0ds_logic_DW01_ash_0 sll_3129 ( .A({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1}), .DATA_TC(1'b0), .SH({Msmhu6, Frmhu6, Ypmhu6, Romhu6, 
        Knmhu6}), .SH_TC(1'b0), .B(Nvkbx6) );
  cortexm0ds_logic_DW01_cmp6_5 eq_3110 ( .A({R9ohu6, Mzihu6, Eyihu6, Wwihu6, 
        Ovihu6, Guihu6, Ysihu6, Qrihu6, Iqihu6, Apihu6, Snihu6, Kmihu6, Clihu6, 
        Ujihu6, Miihu6, Ehihu6, Wfihu6, Oeihu6, Gdihu6, Ybihu6, Qaihu6, I9ihu6, 
        A8ihu6, S6ihu6, K5ihu6, C4ihu6, U2ihu6, M1ihu6, E0ihu6, Wyhhu6, Oxhhu6, 
        Gwhhu6}), .B({E1hpw6, Edkhu6, Wbkhu6}), .TC(1'b0), .EQ(N438) );
  cortexm0ds_logic_DW01_ash_1 sll_3115 ( .A({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1}), .DATA_TC(1'b0), .SH({Oakhu6, G9khu6, Y7khu6, Q6khu6, 
        I5khu6}), .SH_TC(1'b0), .B(Ntkbx6) );
  cortexm0ds_logic_DW01_inc_1 add_3153 ( .A({vis_pc_o[30:2], n8014}), .SUM({
        N5fpw6, SYNOPSYS_UNCONNECTED__0}) );
  cortexm0ds_logic_DW01_add_3 add_3168 ( .A({1'b0, Idfpw6, 1'b0}), .B({1'b0, 
        D5epw6, Qbfpw6, n2535, I4epw6, B4epw6, U3epw6, N3epw6, G3epw6, Z2epw6, 
        L2epw6, X1epw6, Q1epw6, J1epw6, C1epw6, Qbfpw6_10, Q5phu6, W4epw6, 
        S2epw6, E2epw6, Qbfpw6_5, Qbfpw6_4, Qbfpw6_3, Qbfpw6_2, Qbfpw6_1, 
        Qbfpw6_0, 1'b1}), .CI(1'b0), .SUM({\Ozkbx6[33] , \Ozkbx6[32] , 
        \Ozkbx6[31] , \Ozkbx6[30] , \Ozkbx6[29] , \Ozkbx6[28] , \Ozkbx6[27] , 
        \Ozkbx6[26] , \Ozkbx6[25] , \Ozkbx6[24] , \Ozkbx6[23] , \Ozkbx6[22] , 
        \Ozkbx6[21] , \Ozkbx6[20] , \Ozkbx6[19] , \Ozkbx6[18] , \Ozkbx6[17] , 
        \Ozkbx6[16] , \Ozkbx6[15] , \Ozkbx6[14] , \Ozkbx6[13] , \Ozkbx6[12] , 
        \Ozkbx6[11] , \Ozkbx6[10] , \Ozkbx6[9] , \Ozkbx6[8] , \Ozkbx6[7] , 
        \Ozkbx6[6] , \Ozkbx6[5] , \Ozkbx6[4] , \Ozkbx6[3] , \Ozkbx6[2] , 
        \Ozkbx6[1] , SYNOPSYS_UNCONNECTED__1}) );
  cortexm0ds_logic_DW01_add_2 add_3159 ( .A({\Ozkbx6[33] , \Ozkbx6[32] , 
        \Ozkbx6[31] , \Ozkbx6[30] , \Ozkbx6[29] , \Ozkbx6[28] , \Ozkbx6[27] , 
        \Ozkbx6[26] , \Ozkbx6[25] , \Ozkbx6[24] , \Ozkbx6[23] , \Ozkbx6[22] , 
        \Ozkbx6[21] , \Ozkbx6[20] , \Ozkbx6[19] , \Ozkbx6[18] , \Ozkbx6[17] , 
        \Ozkbx6[16] , \Ozkbx6[15] , \Ozkbx6[14] , \Ozkbx6[13] , \Ozkbx6[12] , 
        \Ozkbx6[11] , \Ozkbx6[10] , \Ozkbx6[9] , \Ozkbx6[8] , \Ozkbx6[7] , 
        \Ozkbx6[6] , \Ozkbx6[5] , \Ozkbx6[4] , \Ozkbx6[3] , \Ozkbx6[2] , 
        \Ozkbx6[1] , 1'b0}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, Dqfhu6, 1'b1}), .CI(1'b0), .SUM({Nxkbx6, SYNOPSYS_UNCONNECTED__2}) );
  cortexm0ds_logic_DW02_mult_0 mult_3158 ( .A(Mifpw6), .B(Tgfpw6), .TC(1'b0), 
        .PRODUCT({SYNOPSYS_UNCONNECTED__3, SYNOPSYS_UNCONNECTED__4, 
        SYNOPSYS_UNCONNECTED__5, SYNOPSYS_UNCONNECTED__6, 
        SYNOPSYS_UNCONNECTED__7, SYNOPSYS_UNCONNECTED__8, 
        SYNOPSYS_UNCONNECTED__9, SYNOPSYS_UNCONNECTED__10, 
        SYNOPSYS_UNCONNECTED__11, SYNOPSYS_UNCONNECTED__12, 
        SYNOPSYS_UNCONNECTED__13, SYNOPSYS_UNCONNECTED__14, 
        SYNOPSYS_UNCONNECTED__15, SYNOPSYS_UNCONNECTED__16, 
        SYNOPSYS_UNCONNECTED__17, SYNOPSYS_UNCONNECTED__18, 
        SYNOPSYS_UNCONNECTED__19, SYNOPSYS_UNCONNECTED__20, 
        SYNOPSYS_UNCONNECTED__21, SYNOPSYS_UNCONNECTED__22, 
        SYNOPSYS_UNCONNECTED__23, SYNOPSYS_UNCONNECTED__24, 
        SYNOPSYS_UNCONNECTED__25, SYNOPSYS_UNCONNECTED__26, 
        SYNOPSYS_UNCONNECTED__27, SYNOPSYS_UNCONNECTED__28, 
        SYNOPSYS_UNCONNECTED__29, SYNOPSYS_UNCONNECTED__30, 
        SYNOPSYS_UNCONNECTED__31, SYNOPSYS_UNCONNECTED__32, 
        SYNOPSYS_UNCONNECTED__33, SYNOPSYS_UNCONNECTED__34, Affpw6}) );
  FA_X1 \add_3107/U1_2  ( .A(Tnhpw6[1]), .B(n4142), .CI(n408), .CO(
        \add_3107/carry[3] ), .S(Vrkbx6[2]) );
  FA_X1 \add_3107/U1_3  ( .A(Tnhpw6[2]), .B(\Aphpw6[2] ), .CI(
        \add_3107/carry[3] ), .CO(\add_3107/carry[4] ), .S(Vrkbx6[3]) );
  DFFR_X1 Qsfax6_reg ( .D(n7209), .CK(DCLK), .RN(DBGRESETn), .Q(Dtnhu6), .QN(
        n6913) );
  DFFR_X1 Dugax6_reg ( .D(Wexhu6), .CK(DCLK), .RN(DBGRESETn), .Q(\Aphpw6[2] ), 
        .QN(n7490) );
  DFFR_X1 Ksgax6_reg ( .D(Kfxhu6), .CK(DCLK), .RN(DBGRESETn), .Q(n4142), .QN(
        n7489) );
  DFFS_X1 Nj2qw6_reg ( .D(n7281), .CK(DCLK), .SN(DBGRESETn), .Q(n8176), .QN(
        n6655) );
  DFFS_X1 Jxgax6_reg ( .D(n4157), .CK(DCLK), .SN(DBGRESETn), .Q(n4158), .QN(
        n6909) );
  DFF_X1 Tceax6_reg ( .D(n7124), .CK(DCLK), .QN(n1399) );
  DFF_X1 Opbax6_reg ( .D(n7105), .CK(DCLK), .QN(n1516) );
  DFF_X1 Lx9ax6_reg ( .D(n7135), .CK(DCLK), .Q(K7hpw6[2]), .QN(n6845) );
  DFF_X1 Bvaax6_reg ( .D(n7075), .CK(DCLK), .Q(E1hpw6[2]), .QN(n6792) );
  DFF_X1 Hlcax6_reg ( .D(n7174), .CK(DCLK), .QN(n1122) );
  DFF_X1 Ahdax6_reg ( .D(n7196), .CK(DCLK), .QN(n1257) );
  DFF_X1 Wqdbx6_reg ( .D(n6959), .CK(DCLK), .Q(Trgpw6[20]), .QN(n6716) );
  DFF_X1 Kxeax6_reg ( .D(n6928), .CK(DCLK), .Q(Trgpw6[8]), .QN(n6697) );
  DFF_X1 Hqabx6_reg ( .D(n6943), .CK(DCLK), .Q(Trgpw6[14]), .QN(n6706) );
  DFF_X1 Zycbx6_reg ( .D(n6922), .CK(DCLK), .Q(Trgpw6[27]), .QN(n6690) );
  DFF_X1 Zodbx6_reg ( .D(n6958), .CK(DCLK), .Q(Gtgpw6[20]), .QN(n6715) );
  DFF_X1 Koabx6_reg ( .D(n6942), .CK(DCLK), .Q(Gtgpw6[14]), .QN(n6705) );
  DFF_X1 Facax6_reg ( .D(n6927), .CK(DCLK), .Q(Gtgpw6[8]), .QN(n6696) );
  DFF_X1 Cxcbx6_reg ( .D(n6921), .CK(DCLK), .Q(Gtgpw6[27]), .QN(n6689) );
  DFF_X1 Ureax6_reg ( .D(n7118), .CK(DCLK), .Q(Trgpw6[13]), .QN(n6830) );
  DFF_X1 Rteax6_reg ( .D(n7117), .CK(DCLK), .Q(Trgpw6[12]), .QN(n6829) );
  DFF_X1 N19bx6_reg ( .D(n7004), .CK(DCLK), .Q(Trgpw6[11]), .QN(n6754) );
  DFF_X1 Kpfbx6_reg ( .D(n6989), .CK(DCLK), .Q(Trgpw6[22]), .QN(n6739) );
  DFF_X1 Hpbbx6_reg ( .D(n7109), .CK(DCLK), .Q(Trgpw6[17]), .QN(n6823) );
  DFF_X1 Elgax6_reg ( .D(n7111), .CK(DCLK), .Q(Trgpw6[28]), .QN(n6825) );
  DFF_X1 Q1hbx6_reg ( .D(n6973), .CK(DCLK), .Q(Trgpw6[23]), .QN(n6732) );
  DFF_X1 Oveax6_reg ( .D(n6996), .CK(DCLK), .Q(Trgpw6[10]), .QN(n6747) );
  DFF_X1 Mgeax6_reg ( .D(n7122), .CK(DCLK), .Q(Trgpw6[25]), .QN(n6834) );
  DFF_X1 Jieax6_reg ( .D(n7121), .CK(DCLK), .Q(Trgpw6[24]), .QN(n6833) );
  DFF_X1 Gkeax6_reg ( .D(n6965), .CK(DCLK), .Q(Trgpw6[19]), .QN(n6723) );
  DFF_X1 Dmeax6_reg ( .D(n7120), .CK(DCLK), .Q(Trgpw6[18]), .QN(n6832) );
  DFF_X1 Daebx6_reg ( .D(n7107), .CK(DCLK), .Q(Trgpw6[21]), .QN(n6821) );
  DFF_X1 Xpeax6_reg ( .D(n7019), .CK(DCLK), .Q(Trgpw6[15]), .QN(n6764) );
  DFF_X1 B9jbx6_reg ( .D(n7106), .CK(DCLK), .Q(Trgpw6[9]), .QN(n6820) );
  DFF_X1 Wfcbx6_reg ( .D(n7108), .CK(DCLK), .Q(Trgpw6[26]), .QN(n6822) );
  DFF_X1 Aoeax6_reg ( .D(n7119), .CK(DCLK), .Q(Trgpw6[16]), .QN(n6831) );
  DFF_X1 Hi9bx6_reg ( .D(n7110), .CK(DCLK), .Q(Trgpw6[6]), .QN(n6824) );
  DFF_X1 Gzeax6_reg ( .D(n7116), .CK(DCLK), .Q(Trgpw6[7]), .QN(n6828) );
  DFF_X1 C1fax6_reg ( .D(n7064), .CK(DCLK), .Q(Trgpw6[5]), .QN(n6782) );
  DFF_X1 Y2fax6_reg ( .D(n7115), .CK(DCLK), .Q(Trgpw6[4]), .QN(n6827) );
  DFF_X1 U4fax6_reg ( .D(n7114), .CK(DCLK), .Q(Trgpw6[3]), .QN(n1397) );
  DFF_X1 Fldbx6_reg ( .D(n6961), .CK(DCLK), .Q(K7hpw6[20]), .QN(n6719) );
  DFF_X1 Ab9ax6_reg ( .D(n6967), .CK(DCLK), .Q(K7hpw6[19]), .QN(n6725) );
  DFF_X1 Qkabx6_reg ( .D(n6945), .CK(DCLK), .Q(K7hpw6[14]), .QN(n6709) );
  DFF_X1 Fo9ax6_reg ( .D(n6930), .CK(DCLK), .Q(K7hpw6[8]), .QN(n6699) );
  DFF_X1 Itcbx6_reg ( .D(n6924), .CK(DCLK), .Q(K7hpw6[27]), .QN(n6693) );
  DFF_X1 Rz8bx6_reg ( .D(n7003), .CK(DCLK), .Q(Gtgpw6[11]), .QN(n6753) );
  DFF_X1 P4cax6_reg ( .D(n7099), .CK(DCLK), .Q(Gtgpw6[13]), .QN(n6814) );
  DFF_X1 M6cax6_reg ( .D(n7098), .CK(DCLK), .Q(Gtgpw6[12]), .QN(n6813) );
  DFF_X1 Nnfbx6_reg ( .D(n6988), .CK(DCLK), .Q(Gtgpw6[22]), .QN(n6738) );
  DFF_X1 Knbbx6_reg ( .D(n7090), .CK(DCLK), .Q(Gtgpw6[17]), .QN(n6807) );
  DFF_X1 Hjgax6_reg ( .D(n7092), .CK(DCLK), .Q(Gtgpw6[28]), .QN(n6809) );
  DFF_X1 Yybax6_reg ( .D(n7101), .CK(DCLK), .Q(Gtgpw6[18]), .QN(n6816) );
  DFF_X1 Tzgbx6_reg ( .D(n6972), .CK(DCLK), .Q(Gtgpw6[23]), .QN(n6731) );
  DFF_X1 J8cax6_reg ( .D(n6995), .CK(DCLK), .Q(Gtgpw6[10]), .QN(n6746) );
  DFF_X1 Htbax6_reg ( .D(n7103), .CK(DCLK), .Q(Gtgpw6[25]), .QN(n6818) );
  DFF_X1 G8ebx6_reg ( .D(n7088), .CK(DCLK), .Q(Gtgpw6[21]), .QN(n6805) );
  DFF_X1 Evbax6_reg ( .D(n7102), .CK(DCLK), .Q(Gtgpw6[24]), .QN(n6817) );
  DFF_X1 Bxbax6_reg ( .D(n6964), .CK(DCLK), .Q(Gtgpw6[19]), .QN(n6722) );
  DFF_X1 S2cax6_reg ( .D(n7018), .CK(DCLK), .Q(Gtgpw6[15]), .QN(n6763) );
  DFF_X1 F7jbx6_reg ( .D(n7087), .CK(DCLK), .Q(Gtgpw6[9]), .QN(n6804) );
  DFF_X1 Zdcbx6_reg ( .D(n7089), .CK(DCLK), .Q(Gtgpw6[26]), .QN(n6806) );
  DFF_X1 V0cax6_reg ( .D(n7100), .CK(DCLK), .Q(Gtgpw6[16]), .QN(n6815) );
  DFF_X1 Lg9bx6_reg ( .D(n7091), .CK(DCLK), .Q(Gtgpw6[6]), .QN(n6808) );
  DFF_X1 Bccax6_reg ( .D(n7097), .CK(DCLK), .Q(Gtgpw6[7]), .QN(n6812) );
  DFF_X1 Xdcax6_reg ( .D(n7063), .CK(DCLK), .Q(Gtgpw6[5]), .QN(n6781) );
  DFF_X1 Tfcax6_reg ( .D(n7096), .CK(DCLK), .Q(Gtgpw6[4]), .QN(n6811) );
  DFF_X1 Phcax6_reg ( .D(n7095), .CK(DCLK), .Q(Gtgpw6[3]), .QN(n1515) );
  DFF_X1 Cndbx6_reg ( .D(n6960), .CK(DCLK), .Q(E1hpw6[20]), .QN(n6717) );
  DFF_X1 Q8aax6_reg ( .D(n6966), .CK(DCLK), .Q(E1hpw6[19]), .QN(n6724) );
  DFF_X1 Vlaax6_reg ( .D(n6929), .CK(DCLK), .Q(E1hpw6[8]), .QN(n6698) );
  DFF_X1 Nmabx6_reg ( .D(n6944), .CK(DCLK), .Q(E1hpw6[14]), .QN(n6707) );
  DFF_X1 Fvcbx6_reg ( .D(n6923), .CK(DCLK), .Q(E1hpw6[27]), .QN(n6691) );
  DFF_X1 Wahbx6_reg ( .D(n6969), .CK(DCLK), .Q(K7hpw6[29]), .QN(n6728) );
  DFF_X1 Xv8bx6_reg ( .D(n7006), .CK(DCLK), .Q(K7hpw6[11]), .QN(n6757) );
  DFF_X1 Oi9ax6_reg ( .D(n7140), .CK(DCLK), .Q(K7hpw6[13]), .QN(n6850) );
  DFF_X1 Lk9ax6_reg ( .D(n7139), .CK(DCLK), .Q(K7hpw6[12]), .QN(n6849) );
  DFF_X1 Tjfbx6_reg ( .D(n6991), .CK(DCLK), .Q(K7hpw6[22]), .QN(n6742) );
  DFF_X1 Qjbbx6_reg ( .D(n7130), .CK(DCLK), .Q(K7hpw6[17]), .QN(n6841) );
  DFF_X1 Nfgax6_reg ( .D(n7132), .CK(DCLK), .Q(K7hpw6[28]), .QN(n6843) );
  DFF_X1 Zvgbx6_reg ( .D(n6975), .CK(DCLK), .Q(K7hpw6[23]), .QN(n6734) );
  DFF_X1 Xc9ax6_reg ( .D(n7142), .CK(DCLK), .Q(K7hpw6[18]), .QN(n6852) );
  DFF_X1 M4ebx6_reg ( .D(n7128), .CK(DCLK), .Q(K7hpw6[21]), .QN(n6839) );
  DFF_X1 Im9ax6_reg ( .D(n6998), .CK(DCLK), .Q(K7hpw6[10]), .QN(n6749) );
  DFF_X1 G79ax6_reg ( .D(n7144), .CK(DCLK), .Q(K7hpw6[25]), .QN(n6854) );
  DFF_X1 D99ax6_reg ( .D(n7143), .CK(DCLK), .Q(K7hpw6[24]), .QN(n6853) );
  DFF_X1 Rg9ax6_reg ( .D(n7021), .CK(DCLK), .Q(K7hpw6[15]), .QN(n6767) );
  DFF_X1 N3jbx6_reg ( .D(n7127), .CK(DCLK), .Q(K7hpw6[9]), .QN(n6838) );
  DFF_X1 J59ax6_reg ( .D(n7145), .CK(DCLK), .Q(K7hpw6[30]), .QN(n6855) );
  DFF_X1 Facbx6_reg ( .D(n7129), .CK(DCLK), .Q(K7hpw6[26]), .QN(n6840) );
  DFF_X1 Q2gax6_reg ( .D(n7133), .CK(DCLK), .Q(K7hpw6[31]), .QN(n6844) );
  DFF_X1 Ue9ax6_reg ( .D(n7141), .CK(DCLK), .Q(K7hpw6[16]), .QN(n6851) );
  DFF_X1 Tc9bx6_reg ( .D(n7131), .CK(DCLK), .Q(K7hpw6[6]), .QN(n6842) );
  DFF_X1 Bq9ax6_reg ( .D(n7138), .CK(DCLK), .Q(K7hpw6[7]), .QN(n6848) );
  DFF_X1 Xr9ax6_reg ( .D(n7066), .CK(DCLK), .Q(K7hpw6[5]), .QN(n6784) );
  DFF_X1 Tt9ax6_reg ( .D(n7137), .CK(DCLK), .Q(K7hpw6[4]), .QN(n6847) );
  DFF_X1 Pv9ax6_reg ( .D(n7136), .CK(DCLK), .Q(K7hpw6[3]), .QN(n6846) );
  DFF_X1 Tchbx6_reg ( .D(n6968), .CK(DCLK), .Q(E1hpw6[29]), .QN(n6726) );
  DFF_X1 Ux8bx6_reg ( .D(n7005), .CK(DCLK), .Q(E1hpw6[11]), .QN(n6755) );
  DFF_X1 Egaax6_reg ( .D(n7080), .CK(DCLK), .Q(E1hpw6[13]), .QN(n6797) );
  DFF_X1 Biaax6_reg ( .D(n7079), .CK(DCLK), .Q(E1hpw6[12]), .QN(n6796) );
  DFF_X1 Qlfbx6_reg ( .D(n6990), .CK(DCLK), .Q(E1hpw6[22]), .QN(n6740) );
  DFF_X1 Nlbbx6_reg ( .D(n7070), .CK(DCLK), .Q(E1hpw6[17]), .QN(n6788) );
  DFF_X1 Khgax6_reg ( .D(n7072), .CK(DCLK), .Q(E1hpw6[28]), .QN(n6790) );
  DFF_X1 Yjaax6_reg ( .D(n6997), .CK(DCLK), .Q(E1hpw6[10]), .QN(n6748) );
  DFF_X1 Wxgbx6_reg ( .D(n6974), .CK(DCLK), .Q(E1hpw6[23]), .QN(n6733) );
  DFF_X1 W4aax6_reg ( .D(n7084), .CK(DCLK), .Q(E1hpw6[25]), .QN(n6801) );
  DFF_X1 T6aax6_reg ( .D(n7083), .CK(DCLK), .Q(E1hpw6[24]), .QN(n6800) );
  DFF_X1 Naaax6_reg ( .D(n7082), .CK(DCLK), .Q(E1hpw6[18]), .QN(n6799) );
  DFF_X1 J6ebx6_reg ( .D(n7068), .CK(DCLK), .Q(E1hpw6[21]), .QN(n6786) );
  DFF_X1 Heaax6_reg ( .D(n7020), .CK(DCLK), .Q(E1hpw6[15]), .QN(n6765) );
  DFF_X1 J5jbx6_reg ( .D(n7067), .CK(DCLK), .Q(E1hpw6[9]), .QN(n6785) );
  DFF_X1 Z2aax6_reg ( .D(n7085), .CK(DCLK), .Q(E1hpw6[30]), .QN(n6802) );
  DFF_X1 Cccbx6_reg ( .D(n7069), .CK(DCLK), .Q(E1hpw6[26]), .QN(n6787) );
  DFF_X1 N4gax6_reg ( .D(n7073), .CK(DCLK), .Q(E1hpw6[31]), .QN(n6791) );
  DFF_X1 Kcaax6_reg ( .D(n7081), .CK(DCLK), .Q(E1hpw6[16]), .QN(n6798) );
  DFF_X1 Rnaax6_reg ( .D(n7078), .CK(DCLK), .Q(E1hpw6[7]), .QN(n6795) );
  DFF_X1 Pe9bx6_reg ( .D(n7071), .CK(DCLK), .Q(E1hpw6[6]), .QN(n6789) );
  DFF_X1 Npaax6_reg ( .D(n7065), .CK(DCLK), .Q(E1hpw6[5]), .QN(n6783) );
  DFF_X1 Jraax6_reg ( .D(n7077), .CK(DCLK), .Q(E1hpw6[4]), .QN(n6794) );
  DFF_X1 Ftaax6_reg ( .D(n7076), .CK(DCLK), .Q(E1hpw6[3]), .QN(n6793) );
  DFF_X1 Qudbx6_reg ( .D(n6956), .CK(DCLK), .Q(Togpw6[20]), .QN(n6713) );
  DFF_X1 Y5dax6_reg ( .D(n6925), .CK(DCLK), .Q(Togpw6[8]), .QN(n6694) );
  DFF_X1 Buabx6_reg ( .D(n6940), .CK(DCLK), .Q(Togpw6[14]), .QN(n6703) );
  DFF_X1 T2dbx6_reg ( .D(n6919), .CK(DCLK), .Q(Togpw6[27]), .QN(n6687) );
  DFF_X1 Tsdbx6_reg ( .D(n6957), .CK(DCLK), .Q(Gqgpw6[20]), .QN(n6714) );
  DFF_X1 R1eax6_reg ( .D(n6926), .CK(DCLK), .Q(Gqgpw6[8]), .QN(n6695) );
  DFF_X1 Esabx6_reg ( .D(n6941), .CK(DCLK), .Q(Gqgpw6[14]), .QN(n6704) );
  DFF_X1 W0dbx6_reg ( .D(n6920), .CK(DCLK), .Q(Gqgpw6[27]), .QN(n6688) );
  DFF_X1 I0dax6_reg ( .D(n7169), .CK(DCLK), .Q(Togpw6[13]), .QN(n6867) );
  DFF_X1 F59bx6_reg ( .D(n7001), .CK(DCLK), .Q(Togpw6[11]), .QN(n6751) );
  DFF_X1 F2dax6_reg ( .D(n7168), .CK(DCLK), .Q(Togpw6[12]), .QN(n6866) );
  DFF_X1 Yogax6_reg ( .D(n7162), .CK(DCLK), .Q(Togpw6[28]), .QN(n6862) );
  DFF_X1 Etfbx6_reg ( .D(n6986), .CK(DCLK), .Q(Togpw6[22]), .QN(n6736) );
  DFF_X1 Btbbx6_reg ( .D(n7160), .CK(DCLK), .Q(Togpw6[17]), .QN(n6860) );
  DFF_X1 Xqcax6_reg ( .D(n7172), .CK(DCLK), .Q(Togpw6[24]), .QN(n6870) );
  DFF_X1 Xdebx6_reg ( .D(n7158), .CK(DCLK), .Q(Togpw6[21]), .QN(n6858) );
  DFF_X1 Uscax6_reg ( .D(n6962), .CK(DCLK), .Q(Togpw6[19]), .QN(n6720) );
  DFF_X1 Rucax6_reg ( .D(n7171), .CK(DCLK), .Q(Togpw6[18]), .QN(n6869) );
  DFF_X1 K5hbx6_reg ( .D(n6970), .CK(DCLK), .Q(Togpw6[23]), .QN(n6729) );
  DFF_X1 C4dax6_reg ( .D(n6993), .CK(DCLK), .Q(Togpw6[10]), .QN(n6744) );
  DFF_X1 Apcax6_reg ( .D(n7212), .CK(DCLK), .Q(Togpw6[25]), .QN(n6916) );
  DFF_X1 Lycax6_reg ( .D(n7016), .CK(DCLK), .Q(Togpw6[15]), .QN(n6761) );
  DFF_X1 Tcjbx6_reg ( .D(n7157), .CK(DCLK), .Q(Togpw6[9]), .QN(n6857) );
  DFF_X1 Qjcbx6_reg ( .D(n7159), .CK(DCLK), .Q(Togpw6[26]), .QN(n6859) );
  DFF_X1 Owcax6_reg ( .D(n7170), .CK(DCLK), .Q(Togpw6[16]), .QN(n6868) );
  DFF_X1 Zl9bx6_reg ( .D(n7161), .CK(DCLK), .Q(Togpw6[6]), .QN(n6861) );
  DFF_X1 U7dax6_reg ( .D(n7167), .CK(DCLK), .Q(Togpw6[7]), .QN(n6865) );
  DFF_X1 Q9dax6_reg ( .D(n7061), .CK(DCLK), .Q(Togpw6[5]), .QN(n6779) );
  DFF_X1 Mbdax6_reg ( .D(n7166), .CK(DCLK), .Q(Togpw6[4]), .QN(n6864) );
  DFF_X1 Iddax6_reg ( .D(n7165), .CK(DCLK), .Q(Togpw6[3]), .QN(n1119) );
  DFF_X1 Yxdax6_reg ( .D(n7178), .CK(DCLK), .Q(Gqgpw6[12]), .QN(n6876) );
  DFF_X1 J39bx6_reg ( .D(n7002), .CK(DCLK), .Q(Gqgpw6[11]), .QN(n6752) );
  DFF_X1 Bwdax6_reg ( .D(n7190), .CK(DCLK), .Q(Gqgpw6[13]), .QN(n6891) );
  DFF_X1 Hrfbx6_reg ( .D(n6987), .CK(DCLK), .Q(Gqgpw6[22]), .QN(n6737) );
  DFF_X1 Erbbx6_reg ( .D(n7182), .CK(DCLK), .Q(Gqgpw6[17]), .QN(n6880) );
  DFF_X1 Bngax6_reg ( .D(n7184), .CK(DCLK), .Q(Gqgpw6[28]), .QN(n6883) );
  DFF_X1 Vzdax6_reg ( .D(n6994), .CK(DCLK), .Q(Gqgpw6[10]), .QN(n6745) );
  DFF_X1 Tkdax6_reg ( .D(n7194), .CK(DCLK), .Q(Gqgpw6[25]), .QN(n6896) );
  DFF_X1 Qmdax6_reg ( .D(n7193), .CK(DCLK), .Q(Gqgpw6[24]), .QN(n6895) );
  DFF_X1 Nodax6_reg ( .D(n6963), .CK(DCLK), .Q(Gqgpw6[19]), .QN(n6721) );
  DFF_X1 N3hbx6_reg ( .D(n6971), .CK(DCLK), .Q(Gqgpw6[23]), .QN(n6730) );
  DFF_X1 Kqdax6_reg ( .D(n7192), .CK(DCLK), .Q(Gqgpw6[18]), .QN(n6893) );
  DFF_X1 Acebx6_reg ( .D(n7180), .CK(DCLK), .Q(Gqgpw6[21]), .QN(n6878) );
  DFF_X1 Eudax6_reg ( .D(n7017), .CK(DCLK), .Q(Gqgpw6[15]), .QN(n6762) );
  DFF_X1 Xajbx6_reg ( .D(n7179), .CK(DCLK), .Q(Gqgpw6[9]), .QN(n6877) );
  DFF_X1 Thcbx6_reg ( .D(n7181), .CK(DCLK), .Q(Gqgpw6[26]), .QN(n6879) );
  DFF_X1 Hsdax6_reg ( .D(n7191), .CK(DCLK), .Q(Gqgpw6[16]), .QN(n6892) );
  DFF_X1 N3eax6_reg ( .D(n7189), .CK(DCLK), .Q(Gqgpw6[7]), .QN(n6890) );
  DFF_X1 Dk9bx6_reg ( .D(n7183), .CK(DCLK), .Q(Gqgpw6[6]), .QN(n6881) );
  DFF_X1 J5eax6_reg ( .D(n7062), .CK(DCLK), .Q(Gqgpw6[5]), .QN(n6780) );
  DFF_X1 F7eax6_reg ( .D(n7188), .CK(DCLK), .Q(Gqgpw6[4]), .QN(n6888) );
  DFF_X1 B9eax6_reg ( .D(n7187), .CK(DCLK), .Q(Gqgpw6[3]), .QN(n1256) );
  DFF_X1 Yf1qw6_reg ( .D(n7913), .CK(DCLK), .Q(Jshpw6[9]), .QN(n7407) );
  DFF_X1 Ke1qw6_reg ( .D(n7914), .CK(DCLK), .Q(Jshpw6[8]), .QN(n7406) );
  DFF_X1 Vn9bx6_reg ( .D(n7916), .CK(DCLK), .Q(Jshpw6[6]), .QN(n7632) );
  DFF_X1 Nd3qw6_reg ( .D(n7915), .CK(DCLK), .Q(Jshpw6[7]), .QN(n7422) );
  DFF_X1 Bf3qw6_reg ( .D(n7917), .CK(DCLK), .Q(Jshpw6[5]), .QN(n7423) );
  DFF_X1 Vj3qw6_reg ( .D(n7854), .CK(DCLK), .Q(Tnhpw6[1]), .QN(n7426) );
  DFF_X1 Pg3qw6_reg ( .D(n7918), .CK(DCLK), .Q(Jshpw6[4]), .QN(n7424) );
  DFF_X1 P23qw6_reg ( .D(n7919), .CK(DCLK), .Q(Tnhpw6[3]), .QN(n7418) );
  DFF_X1 Xn7ax6_reg ( .D(n7920), .CK(DCLK), .Q(Tnhpw6[2]), .QN(n7441) );
  DFF_X1 Qehbx6_reg ( .D(n7921), .CK(DCLK), .Q(Tnhpw6[0]), .QN(n7683) );
  DFF_X1 X5bax6_reg ( .D(n7151), .CK(DCLK), .QN(n7458) );
  DFF_X1 T7bax6_reg ( .D(n7150), .CK(DCLK), .QN(n7459) );
  DFF_X1 Pkkbx6_reg ( .D(n7147), .CK(DCLK), .QN(n7708) );
  DFF_X1 Hdbax6_reg ( .D(n7156), .CK(DCLK), .QN(n7462) );
  DFF_X1 Dfbax6_reg ( .D(n7155), .CK(DCLK), .QN(n7463) );
  DFF_X1 Tikbx6_reg ( .D(n7152), .CK(DCLK), .QN(n7707) );
  DFF_X1 P9bax6_reg ( .D(n7149), .CK(DCLK), .QN(n7460) );
  DFF_X1 Lbbax6_reg ( .D(n7148), .CK(DCLK), .QN(n7461) );
  DFF_X1 Zgbax6_reg ( .D(n7154), .CK(DCLK), .QN(n7464) );
  DFF_X1 Vibax6_reg ( .D(n7153), .CK(DCLK), .QN(n7465) );
  DFF_X1 Hz9ax6_reg ( .D(n7134), .CK(DCLK), .Q(n4408), .QN(n7454) );
  DFF_X1 N39ax6_reg ( .D(n7146), .CK(DCLK), .QN(n6856) );
  DFF_X1 Xwaax6_reg ( .D(n7074), .CK(DCLK), .QN(n7455) );
  DFF_X1 D1aax6_reg ( .D(n7086), .CK(DCLK), .QN(n6803) );
  DFF_X1 Peeax6_reg ( .D(n7123), .CK(DCLK), .QN(n7474) );
  DFF_X1 H8gax6_reg ( .D(n7112), .CK(DCLK), .QN(n7484) );
  DFF_X1 Krbax6_reg ( .D(n7104), .CK(DCLK), .QN(n7468) );
  DFF_X1 K6gax6_reg ( .D(n7093), .CK(DCLK), .QN(n7483) );
  DFF_X1 Bt2qw6_reg ( .D(I0xhu6), .CK(DCLK), .QN(n7415) );
  DFF_X1 Fm7ax6_reg ( .D(P0xhu6), .CK(DCLK), .QN(n7440) );
  DFF_X1 Dncax6_reg ( .D(n7173), .CK(DCLK), .QN(n7470) );
  DFF_X1 Bcgax6_reg ( .D(n7163), .CK(DCLK), .QN(n7486) );
  DFF_X1 Widax6_reg ( .D(n7195), .CK(DCLK), .Q(n4335), .QN(n7472) );
  DFF_X1 Eagax6_reg ( .D(n7185), .CK(DCLK), .Q(n4336), .QN(n7485) );
  DFF_X1 A3ipw6_reg ( .D(X3yhu6), .CK(DCLK), .QN(n7250) );
  DFF_X1 Cq3qw6_reg ( .D(M9xhu6), .CK(DCLK), .Q(n8206), .QN(n7430) );
  DFF_X1 Kl8ax6_reg ( .D(Udxhu6), .CK(DCLK), .Q(n4145), .QN(n7447) );
  DFF_X1 Su8ax6_reg ( .D(Bexhu6), .CK(DCLK), .Q(n4402), .QN(n7450) );
  DFF_X1 B79bx6_reg ( .D(Iexhu6), .CK(DCLK), .Q(n8164), .QN(n7631) );
  DFF_X1 Yubbx6_reg ( .D(Scxhu6), .CK(DCLK), .QN(n7648) );
  DFF_X1 Vqgax6_reg ( .D(T9xhu6), .CK(DCLK), .QN(n7488) );
  DFF_X1 Nwdbx6_reg ( .D(Xbxhu6), .CK(DCLK), .QN(n7661) );
  DFF_X1 Bvfbx6_reg ( .D(Jbxhu6), .CK(DCLK), .QN(n7667) );
  DFF_X1 Ufebx6_reg ( .D(Qbxhu6), .CK(DCLK), .QN(n7664) );
  DFF_X1 Q2ibx6_reg ( .D(Oaxhu6), .CK(DCLK), .QN(n7693) );
  DFF_X1 No3qw6_reg ( .D(Vaxhu6), .CK(DCLK), .Q(n3389), .QN(n7429) );
  DFF_X1 H4ypw6_reg ( .D(Pexhu6), .CK(DCLK), .Q(n8172), .QN(n7397) );
  DFF_X1 Ym3qw6_reg ( .D(Ecxhu6), .CK(DCLK), .QN(n7428) );
  DFF_X1 Jl3qw6_reg ( .D(Lcxhu6), .CK(DCLK), .QN(n7427) );
  DFF_X1 H7hbx6_reg ( .D(Cbxhu6), .CK(DCLK), .QN(n7681) );
  DFF_X1 Yvabx6_reg ( .D(Ndxhu6), .CK(DCLK), .Q(n8253), .QN(n7641) );
  DFF_X1 Ad7ax6_reg ( .D(Gdxhu6), .CK(DCLK), .QN(n7437) );
  DFF_X1 Wc2qw6_reg ( .D(F9xhu6), .CK(DCLK), .Q(n4151), .QN(n7410) );
  DFF_X1 Nlcbx6_reg ( .D(Haxhu6), .CK(DCLK), .QN(n7655) );
  DFF_X1 Q4dbx6_reg ( .D(Aaxhu6), .CK(DCLK), .QN(n7657) );
  DFF_X1 Ydgax6_reg ( .D(O2yhu6), .CK(DCLK), .Q(n3880), .QN(n7487) );
  DFF_X1 Dpwpw6_reg ( .D(Zcxhu6), .CK(DCLK), .QN(n7387) );
  DFF_X1 Ceabx6_reg ( .D(n7895), .CK(DCLK), .QN(n7640) );
  DFF_X1 Idqpw6_reg ( .D(n7897), .CK(DCLK), .Q(n3004), .QN(n7345) );
  DFF_X1 L9bbx6_reg ( .D(n7900), .CK(DCLK), .QN(n7646) );
  DFF_X1 H3lpw6_reg ( .D(n7890), .CK(DCLK), .QN(n7292) );
  DFF_X1 Kswpw6_reg ( .D(n7891), .CK(DCLK), .Q(n4055), .QN(n7389) );
  DFF_X1 Vefax6_reg ( .D(n7909), .CK(DCLK), .Q(n4297), .QN(n6649) );
  DFF_X1 Rr3qw6_reg ( .D(n7896), .CK(DCLK), .Q(n8205) );
  DFF_X1 Gyxpw6_reg ( .D(n7905), .CK(DCLK), .QN(n7396) );
  DFF_X1 M81qw6_reg ( .D(n7907), .CK(DCLK), .QN(n7405) );
  DFF_X1 Cncbx6_reg ( .D(n7892), .CK(DCLK), .QN(n6658) );
  DFF_X1 Bu6bx6_reg ( .D(n7904), .CK(DCLK), .QN(n6652) );
  DFF_X1 X42qw6_reg ( .D(n7878), .CK(DCLK), .Q(n3125) );
  DFF_X1 Uunpw6_reg ( .D(n7898), .CK(DCLK), .Q(n3877) );
  DFF_X1 Gbvpw6_reg ( .D(n7899), .CK(DCLK), .QN(n6656) );
  DFF_X1 N0cbx6_reg ( .D(n7901), .CK(DCLK), .QN(n7650) );
  DFF_X1 Mh1qw6_reg ( .D(n7906), .CK(DCLK), .QN(n6651) );
  DFF_X1 F8dbx6_reg ( .D(n7855), .CK(DCLK), .QN(n7659) );
  DFF_X1 Ro8ax6_reg ( .D(n7873), .CK(DCLK), .QN(n7449) );
  DFF_X1 Z67ax6_reg ( .D(n7874), .CK(DCLK), .QN(n6666) );
  DFF_X1 Sd8ax6_reg ( .D(n7872), .CK(DCLK), .QN(n6667) );
  DFF_X1 Qwfbx6_reg ( .D(n7879), .CK(DCLK), .QN(n6662) );
  DFF_X1 Pdbbx6_reg ( .D(n7876), .CK(DCLK), .QN(n6664) );
  DFF_X1 Jhebx6_reg ( .D(n7893), .CK(DCLK), .QN(n7665) );
  DFF_X1 Cydbx6_reg ( .D(n7894), .CK(DCLK), .QN(n7662) );
  DFF_X1 Cjwpw6_reg ( .D(n7877), .CK(DCLK), .QN(n7386) );
  DFF_X1 Fl2qw6_reg ( .D(n7902), .CK(DCLK), .QN(n7413) );
  DFF_X1 Ggabx6_reg ( .D(n7875), .CK(DCLK), .Q(n3042), .QN(n6665) );
  DFFR_X1 Xxqpw6_reg ( .D(Q7ohu6), .CK(DCLK), .RN(DBGRESETn), .QN(n6914) );
  DFFR_X1 R19ax6_reg ( .D(L5xhu6), .CK(DCLK), .RN(DBGRESETn), .QN(n7453) );
  DFFR_X1 Vz8ax6_reg ( .D(n7350), .CK(DCLK), .RN(DBGRESETn), .QN(n6643) );
  DFFR_X1 Sbfax6_reg ( .D(n7125), .CK(DCLK), .RN(DBGRESETn), .QN(n6836) );
  DFFR_X1 Zx8ax6_reg ( .D(Z5xhu6), .CK(DCLK), .RN(DBGRESETn), .QN(n7452) );
  DFFR_X1 H4bax6_reg ( .D(n7208), .CK(DCLK), .RN(DBGRESETn), .Q(n4141), .QN(
        n7457) );
  DFFR_X1 Eafax6_reg ( .D(n7126), .CK(DCLK), .RN(DBGRESETn), .QN(n6837) );
  DFFR_X1 Xnbax6_reg ( .D(n7853), .CK(DCLK), .RN(DBGRESETn), .QN(n7467) );
  DFFR_X1 Q6fax6_reg ( .D(n7113), .CK(DCLK), .RN(DBGRESETn), .QN(n7475) );
  DFFR_X1 Ljcax6_reg ( .D(n7094), .CK(DCLK), .RN(DBGRESETn), .QN(n7469) );
  DFFR_X1 L2bax6_reg ( .D(n7175), .CK(DCLK), .RN(DBGRESETn), .QN(n6873) );
  DFFR_X1 P0bax6_reg ( .D(n7176), .CK(DCLK), .RN(DBGRESETn), .QN(n7456) );
  DFFR_X1 Tyaax6_reg ( .D(n7177), .CK(DCLK), .RN(DBGRESETn), .QN(n6874) );
  DFFR_X1 Hdfax6_reg ( .D(n6992), .CK(DCLK), .RN(DBGRESETn), .QN(n6743) );
  DFFR_X1 Tb3qw6_reg ( .D(Dfxhu6), .CK(DCLK), .RN(DBGRESETn), .Q(n4144), .QN(
        n7421) );
  DFFR_X1 Efdax6_reg ( .D(n7164), .CK(DCLK), .RN(DBGRESETn), .QN(n7471) );
  DFFR_X1 Xaeax6_reg ( .D(n7186), .CK(DCLK), .RN(DBGRESETn), .QN(n7473) );
  DFFR_X1 Gr2qw6_reg ( .D(W0xhu6), .CK(DCLK), .RN(DBGRESETn), .Q(n1840), .QN(
        n7414) );
  DFFR_X1 Thiax6_reg ( .D(n8012), .CK(DCLK), .RN(DBGRESETn), .Q(n8285), .QN(
        n6645) );
  DFFR_X1 Uh2qw6_reg ( .D(n7940), .CK(DCLK), .RN(DBGRESETn), .QN(n6653) );
  DFFR_X1 Hmbax6_reg ( .D(n8009), .CK(DCLK), .RN(DBGRESETn), .Q(n8162), .QN(
        n6647) );
  DFFR_X1 Wvgax6_reg ( .D(n7207), .CK(DCLK), .RN(DBGRESETn), .Q(n4152), .QN(
        n7491) );
  DFFR_X1 M8fax6_reg ( .D(n8011), .CK(DCLK), .RN(DBGRESETn), .Q(n4341), .QN(
        n7476) );
  DFFR_X1 Lmkbx6_reg ( .D(Pfphu6), .CK(DCLK), .RN(DBGRESETn), .QN(n6659) );
  DFFR_X1 Uofax6_reg ( .D(n7923), .CK(DCLK), .RN(DBGRESETn), .Q(n4112), .QN(
        n7480) );
  DFFR_X1 Sqfax6_reg ( .D(n2100), .CK(DCLK), .RN(DBGRESETn), .Q(n4116), .QN(
        n7481) );
  DFFR_X1 Dg2qw6_reg ( .D(n7883), .CK(DCLK), .RN(DBGRESETn), .Q(n4140), .QN(
        n7412) );
  DFFR_X1 Pe7ax6_reg ( .D(n7885), .CK(DCLK), .RN(DBGRESETn), .Q(n4329), .QN(
        n7438) );
  DFFR_X1 Le2qw6_reg ( .D(n7884), .CK(DCLK), .RN(DBGRESETn), .Q(n3913), .QN(
        n7411) );
  DFFR_X1 Hw8ax6_reg ( .D(n7882), .CK(DCLK), .RN(DBGRESETn), .Q(n4405), .QN(
        n7451) );
  DFFR_X1 Di3qw6_reg ( .D(n7887), .CK(DCLK), .RN(DBGRESETn), .Q(n4054), .QN(
        n7425) );
  DFFR_X1 Zm8ax6_reg ( .D(n7888), .CK(DCLK), .RN(DBGRESETn), .Q(n3882), .QN(
        n7448) );
  DFFR_X1 Sqwpw6_reg ( .D(n7889), .CK(DCLK), .RN(DBGRESETn), .Q(n3470), .QN(
        n7388) );
  DFFR_X1 D43qw6_reg ( .D(n7886), .CK(DCLK), .RN(DBGRESETn), .Q(n4406), .QN(
        n7419) );
  DFFR_X1 Pexpw6_reg ( .D(n7738), .CK(DCLK), .RN(DBGRESETn), .QN(n7392) );
  DFFR_X1 Jvvpw6_reg ( .D(n7737), .CK(DCLK), .RN(DBGRESETn), .QN(n7380) );
  DFFR_X1 Vpkpw6_reg ( .D(n7730), .CK(DCLK), .RN(DBGRESETn), .QN(n7291) );
  DFFR_X1 F4ibx6_reg ( .D(n7728), .CK(DCLK), .RN(DBGRESETn), .QN(n7694) );
  DFFR_X1 Rkbax6_reg ( .D(n7729), .CK(DCLK), .RN(DBGRESETn), .QN(n7466) );
  DFFS_X1 J0iax6_reg ( .D(n8013), .CK(HCLK), .SN(HRESETn), .Q(n5284), .QN(
        n7493) );
  DFFS_X1 L6lax6_reg ( .D(n7027), .CK(HCLK), .SN(HRESETn), .Q(n4667), .QN(
        n7532) );
  DFFS_X1 Tajax6_reg ( .D(n7025), .CK(HCLK), .SN(HRESETn), .Q(n4699), .QN(
        n6770) );
  DFFS_X1 P5vpw6_reg ( .D(n8004), .CK(HCLK), .SN(HRESETn), .Q(n479), .QN(n237)
         );
  DFFS_X1 Hgrpw6_reg ( .D(n7939), .CK(HCLK), .SN(HRESETn), .Q(n3549), .QN(
        n7354) );
  DFFS_X1 Dxvpw6_reg ( .D(n7936), .CK(HCLK), .SN(HRESETn), .Q(n476), .QN(n7381) );
  DFFS_X1 N4kax6_reg ( .D(n7929), .CK(HCLK), .SN(HRESETn), .Q(n4670), .QN(
        n7519) );
  DFFS_X1 Wkipw6_reg ( .D(n7925), .CK(HCLK), .SN(HRESETn), .Q(n4932), .QN(
        n7259) );
  DFFS_X1 Wfspw6_reg ( .D(n7935), .CK(HCLK), .SN(HRESETn), .Q(n3690), .QN(
        n7359) );
  DFFS_X1 S7mpw6_reg ( .D(n7852), .CK(HCLK), .SN(HRESETn), .Q(n4908), .QN(
        n7325) );
  DFFS_X1 Irmpw6_reg ( .D(n7924), .CK(HCLK), .SN(HRESETn), .Q(n4910), .QN(
        n7329) );
  DFFS_X1 U9ypw6_reg ( .D(n7938), .CK(HCLK), .SN(HRESETn), .Q(n4187), .QN(
        n7399) );
  DFFS_X1 Skjax6_reg ( .D(n7933), .CK(HCLK), .SN(HRESETn), .Q(n4635), .QN(
        n7510) );
  DFFS_X1 Rwjax6_reg ( .D(n7930), .CK(HCLK), .SN(HRESETn), .Q(n5042), .QN(
        n7516) );
  DFFS_X1 P0kax6_reg ( .D(n7934), .CK(HCLK), .SN(HRESETn), .Q(n4572), .QN(
        n7518) );
  DFFS_X1 W4jax6_reg ( .D(n7928), .CK(HCLK), .SN(HRESETn), .Q(n4993), .QN(
        n7505) );
  DFFS_X1 Ssjax6_reg ( .D(n7931), .CK(HCLK), .SN(HRESETn), .Q(n470), .QN(n7514) );
  DFFS_X1 Sojax6_reg ( .D(n7932), .CK(HCLK), .SN(HRESETn), .Q(n475), .QN(n270)
         );
  DFFS_X1 P14qw6_reg ( .D(n7937), .CK(HCLK), .SN(HRESETn), .Q(n2262), .QN(
        n7433) );
  DFFS_X1 Jgxpw6_reg ( .D(n7926), .CK(HCLK), .SN(HRESETn), .Q(n4978), .QN(
        n7393) );
  DFFS_X1 Jckax6_reg ( .D(n7927), .CK(HCLK), .SN(HRESETn), .Q(n4987), .QN(
        n7523) );
  DFFS_X1 F26bx6_reg ( .D(Ruphu6), .CK(HCLK), .SN(HRESETn), .QN(n7628) );
  DFFS_X1 Sz3qw6_reg ( .D(n7213), .CK(HCLK), .SN(HRESETn), .QN(n6769) );
  DFFR_X1 Mnmpw6_reg ( .D(n7957), .CK(HCLK), .RN(HRESETn), .Q(n6681), .QN(
        n3775) );
  DFFR_X1 Xfiax6_reg ( .D(Xdvhu6), .CK(HCLK), .RN(HRESETn), .Q(vis_primask_o), 
        .QN(n3114) );
  DFFR_X1 Npypw6_reg ( .D(Brrhu6), .CK(HCLK), .RN(HRESETn), .Q(vis_control_o), 
        .QN(n4364) );
  DFFR_X1 Qakbx6_reg ( .D(n8015), .CK(HCLK), .RN(HRESETn), .QN(n4546) );
  DFFR_X1 Halax6_reg ( .D(n8016), .CK(HCLK), .RN(HRESETn), .QN(n5256) );
  DFFR_X1 Vbkpw6_reg ( .D(n7849), .CK(HCLK), .RN(HRESETn), .Q(vis_ipsr_o[5]), 
        .QN(n5126) );
  DFFR_X1 Qhmpw6_reg ( .D(n7844), .CK(HCLK), .RN(HRESETn), .Q(vis_ipsr_o[3]), 
        .QN(n5088) );
  DFFR_X1 Aniax6_reg ( .D(n7847), .CK(HCLK), .RN(HRESETn), .Q(vis_ipsr_o[2]), 
        .QN(n5111) );
  DFFR_X1 Ijiax6_reg ( .D(n7845), .CK(HCLK), .RN(HRESETn), .Q(vis_ipsr_o[4]), 
        .QN(n5105) );
  DFFR_X1 Qijpw6_reg ( .D(Bgvhu6), .CK(HCLK), .RN(HRESETn), .Q(vis_apsr_o[1]), 
        .QN(n2729) );
  DFFR_X1 X5ibx6_reg ( .D(n7727), .CK(HCLK), .RN(HRESETn), .Q(vis_apsr_o[0]), 
        .QN(n8260) );
  DFF_X1 Vqjbx6_reg ( .D(n8023), .CK(HCLK), .Q(n6641), .QN(n4702) );
  DFF_X1 Usjbx6_reg ( .D(n8022), .CK(HCLK), .QN(n4701) );
  DFF_X1 Tujbx6_reg ( .D(n8021), .CK(HCLK), .QN(n4700) );
  DFF_X1 Tcjax6_reg ( .D(n8035), .CK(HCLK), .QN(n3673) );
  DFF_X1 Sejax6_reg ( .D(n8034), .CK(HCLK), .QN(n5270) );
  DFF_X1 O2kax6_reg ( .D(n8027), .CK(HCLK), .Q(n6640), .QN(n4708) );
  DFF_X1 Ua9bx6_reg ( .D(n7810), .CK(HCLK), .Q(n6679) );
  DFF_X1 I1lpw6_reg ( .D(n7828), .CK(HCLK), .Q(n6676), .QN(n3115) );
  DFF_X1 Y7upw6_reg ( .D(Zqqhu6), .CK(HCLK), .Q(vis_r0_o[17]), .QN(n6280) );
  DFF_X1 C5wpw6_reg ( .D(Kmqhu6), .CK(HCLK), .Q(vis_r0_o[16]), .QN(n6330) );
  DFF_X1 Wdmax6_reg ( .D(Exqhu6), .CK(HCLK), .Q(vis_r10_o[18]), .QN(n8191) );
  DFF_X1 V1vax6_reg ( .D(Sxqhu6), .CK(HCLK), .Q(vis_r4_o[18]), .QN(n8182) );
  DFF_X1 Uwqax6_reg ( .D(Cwqhu6), .CK(HCLK), .Q(vis_r2_o[18]), .QN(n8192) );
  DFF_X1 Tc0qw6_reg ( .D(Izqhu6), .CK(HCLK), .Q(vis_msp_o[16]), .QN(n8189) );
  DFF_X1 Pcxpw6_reg ( .D(Pzqhu6), .CK(HCLK), .Q(vis_psp_o[16]), .QN(n8184) );
  DFF_X1 Paxpw6_reg ( .D(Zxqhu6), .CK(HCLK), .Q(vis_r5_o[18]), .QN(n8178) );
  DFF_X1 P8xpw6_reg ( .D(Lxqhu6), .CK(HCLK), .Q(vis_r11_o[18]), .QN(n8187) );
  DFF_X1 P6xpw6_reg ( .D(Xwqhu6), .CK(HCLK), .Q(vis_r9_o[18]), .QN(n8179) );
  DFF_X1 P4xpw6_reg ( .D(Vvqhu6), .CK(HCLK), .Q(vis_r1_o[18]), .QN(n8180) );
  DFF_X1 P2xpw6_reg ( .D(Ovqhu6), .CK(HCLK), .Q(vis_r0_o[18]), .QN(n8185) );
  DFF_X1 O0sax6_reg ( .D(Qwqhu6), .CK(HCLK), .Q(vis_r8_o[18]), .QN(n8183) );
  DFF_X1 Nvnax6_reg ( .D(Bzqhu6), .CK(HCLK), .Q(vis_r14_o[18]), .QN(n8194) );
  DFF_X1 Llwax6_reg ( .D(Nyqhu6), .CK(HCLK), .Q(vis_r7_o[18]), .QN(n8186) );
  DFF_X1 Ektax6_reg ( .D(Uyqhu6), .CK(HCLK), .Q(vis_r12_o[18]), .QN(n8181) );
  DFF_X1 Edpax6_reg ( .D(Gyqhu6), .CK(HCLK), .Q(vis_r6_o[18]), .QN(n8190) );
  DFF_X1 Da6bx6_reg ( .D(Jwqhu6), .CK(HCLK), .Q(vis_r3_o[18]), .QN(n8188) );
  DFF_X1 Yhupw6_reg ( .D(Avqhu6), .CK(HCLK), .Q(vis_psp_o[15]), .QN(n3279) );
  DFF_X1 Yfupw6_reg ( .D(Ktqhu6), .CK(HCLK), .Q(vis_r5_o[17]), .QN(n6564) );
  DFF_X1 Ydupw6_reg ( .D(Wsqhu6), .CK(HCLK), .Q(vis_r11_o[17]), .QN(n8109) );
  DFF_X1 Ybupw6_reg ( .D(Isqhu6), .CK(HCLK), .Q(vis_r9_o[17]), .QN(n6150) );
  DFF_X1 Y9upw6_reg ( .D(Grqhu6), .CK(HCLK), .Q(vis_r1_o[17]), .QN(n6771) );
  DFF_X1 Whmax6_reg ( .D(Aoqhu6), .CK(HCLK), .Q(vis_r10_o[16]), .QN(n4004) );
  DFF_X1 Wfmax6_reg ( .D(Psqhu6), .CK(HCLK), .Q(vis_r10_o[17]), .QN(n8059) );
  DFF_X1 V5vax6_reg ( .D(Ooqhu6), .CK(HCLK), .Q(vis_r4_o[16]), .QN(n5386) );
  DFF_X1 V3vax6_reg ( .D(Dtqhu6), .CK(HCLK), .Q(vis_r4_o[17]), .QN(n5460) );
  DFF_X1 Uyqax6_reg ( .D(Nrqhu6), .CK(HCLK), .Q(vis_r2_o[17]), .QN(n5532) );
  DFF_X1 U0rax6_reg ( .D(Ymqhu6), .CK(HCLK), .Q(vis_r2_o[16]), .QN(n5465) );
  DFF_X1 Tg0qw6_reg ( .D(Eqqhu6), .CK(HCLK), .Q(vis_msp_o[14]), .QN(n5989) );
  DFF_X1 Te0qw6_reg ( .D(Tuqhu6), .CK(HCLK), .Q(vis_msp_o[15]), .QN(n5924) );
  DFF_X1 O4sax6_reg ( .D(Mnqhu6), .CK(HCLK), .Q(vis_r8_o[16]), .QN(n5875) );
  DFF_X1 O2sax6_reg ( .D(Bsqhu6), .CK(HCLK), .Q(vis_r8_o[17]), .QN(n5897) );
  DFF_X1 Nznax6_reg ( .D(Xpqhu6), .CK(HCLK), .Q(vis_r14_o[16]), .QN(n8075) );
  DFF_X1 Nxnax6_reg ( .D(Muqhu6), .CK(HCLK), .Q(vis_r14_o[17]), .QN(n8089) );
  DFF_X1 Lpwax6_reg ( .D(Jpqhu6), .CK(HCLK), .Q(vis_r7_o[16]), .QN(n7797) );
  DFF_X1 Lnwax6_reg ( .D(Ytqhu6), .CK(HCLK), .Q(vis_r7_o[17]), .QN(n7745) );
  DFF_X1 Eotax6_reg ( .D(Qpqhu6), .CK(HCLK), .Q(vis_r12_o[16]), .QN(n6218) );
  DFF_X1 Emtax6_reg ( .D(Fuqhu6), .CK(HCLK), .Q(vis_r12_o[17]), .QN(n6257) );
  DFF_X1 Ehpax6_reg ( .D(Cpqhu6), .CK(HCLK), .Q(vis_r6_o[16]), .QN(n5810) );
  DFF_X1 Efpax6_reg ( .D(Rtqhu6), .CK(HCLK), .Q(vis_r6_o[17]), .QN(n5709) );
  DFF_X1 De6bx6_reg ( .D(Fnqhu6), .CK(HCLK), .Q(vis_r3_o[16]), .QN(n7580) );
  DFF_X1 Dc6bx6_reg ( .D(Urqhu6), .CK(HCLK), .Q(vis_r3_o[17]), .QN(n7261) );
  DFF_X1 Cfwpw6_reg ( .D(Lqqhu6), .CK(HCLK), .Q(vis_psp_o[14]), .QN(n4003) );
  DFF_X1 Cdwpw6_reg ( .D(Voqhu6), .CK(HCLK), .Q(vis_r5_o[16]), .QN(n6478) );
  DFF_X1 Cbwpw6_reg ( .D(Hoqhu6), .CK(HCLK), .Q(vis_r11_o[16]), .QN(n8128) );
  DFF_X1 C9wpw6_reg ( .D(Tnqhu6), .CK(HCLK), .Q(vis_r9_o[16]), .QN(n6119) );
  DFF_X1 C7wpw6_reg ( .D(Rmqhu6), .CK(HCLK), .Q(vis_r1_o[16]), .QN(n6636) );
  DFF_X1 Zz7bx6_reg ( .D(Xiqhu6), .CK(HCLK), .Q(vis_r8_o[15]), .QN(n5825) );
  DFF_X1 Zx7bx6_reg ( .D(Qiqhu6), .CK(HCLK), .Q(vis_r3_o[15]), .QN(n7372) );
  DFF_X1 Zv7bx6_reg ( .D(Jiqhu6), .CK(HCLK), .Q(vis_r2_o[15]), .QN(n5552) );
  DFF_X1 Zt7bx6_reg ( .D(Ciqhu6), .CK(HCLK), .Q(vis_r1_o[15]), .QN(n6835) );
  DFF_X1 Zr7bx6_reg ( .D(Vhqhu6), .CK(HCLK), .Q(vis_r0_o[15]), .QN(n6292) );
  DFF_X1 Zl8bx6_reg ( .D(Wlqhu6), .CK(HCLK), .Q(vis_psp_o[13]), .QN(n3583) );
  DFF_X1 Zj8bx6_reg ( .D(Plqhu6), .CK(HCLK), .Q(vis_msp_o[13]), .QN(n5941) );
  DFF_X1 Zh8bx6_reg ( .D(Ilqhu6), .CK(HCLK), .Q(vis_r14_o[15]), .QN(n8096) );
  DFF_X1 Zf8bx6_reg ( .D(Blqhu6), .CK(HCLK), .Q(vis_r12_o[15]), .QN(n2490) );
  DFF_X1 Zd8bx6_reg ( .D(Ukqhu6), .CK(HCLK), .Q(vis_r7_o[15]), .QN(n7766) );
  DFF_X1 Zb8bx6_reg ( .D(Nkqhu6), .CK(HCLK), .Q(vis_r6_o[15]), .QN(n5729) );
  DFF_X1 Z98bx6_reg ( .D(Gkqhu6), .CK(HCLK), .Q(vis_r5_o[15]), .QN(n6585) );
  DFF_X1 Z78bx6_reg ( .D(Zjqhu6), .CK(HCLK), .Q(vis_r4_o[15]), .QN(n5317) );
  DFF_X1 Z58bx6_reg ( .D(Sjqhu6), .CK(HCLK), .Q(vis_r11_o[15]), .QN(n8115) );
  DFF_X1 Z38bx6_reg ( .D(Ljqhu6), .CK(HCLK), .Q(vis_r10_o[15]), .QN(n8065) );
  DFF_X1 Z18bx6_reg ( .D(Ejqhu6), .CK(HCLK), .Q(vis_r9_o[15]), .QN(n6168) );
  DFF_X1 Zrlax6_reg ( .D(Ehshu6), .CK(HCLK), .Q(vis_r10_o[6]), .QN(n8070) );
  DFF_X1 Z3spw6_reg ( .D(Xgshu6), .CK(HCLK), .Q(vis_r9_o[6]), .QN(n6039) );
  DFF_X1 Yfuax6_reg ( .D(Shshu6), .CK(HCLK), .Q(vis_r4_o[6]), .QN(n5352) );
  DFF_X1 Y5spw6_reg ( .D(Lhshu6), .CK(HCLK), .Q(vis_r11_o[6]), .QN(n8122) );
  DFF_X1 Xaqax6_reg ( .D(Jgshu6), .CK(HCLK), .Q(vis_r2_o[6]), .QN(n5555) );
  DFF_X1 X7spw6_reg ( .D(Zhshu6), .CK(HCLK), .Q(vis_r5_o[6]), .QN(n6394) );
  DFF_X1 W9spw6_reg ( .D(Dkshu6), .CK(HCLK), .Q(vis_r8_o[6]), .QN(n5894) );
  DFF_X1 Vszpw6_reg ( .D(Ijshu6), .CK(HCLK), .Q(vis_msp_o[4]), .QN(n5960) );
  DFF_X1 Pe5bx6_reg ( .D(Qgshu6), .CK(HCLK), .Q(vis_r3_o[6]), .QN(n7376) );
  DFF_X1 Pbnax6_reg ( .D(Bjshu6), .CK(HCLK), .Q(vis_r14_o[6]), .QN(n4280) );
  DFF_X1 Ozvax6_reg ( .D(Nishu6), .CK(HCLK), .Q(vis_r7_o[6]), .QN(n7781) );
  DFF_X1 Hysax6_reg ( .D(Uishu6), .CK(HCLK), .Q(vis_r12_o[6]), .QN(n6188) );
  DFF_X1 Hroax6_reg ( .D(Gishu6), .CK(HCLK), .Q(vis_r6_o[6]), .QN(n5793) );
  DFF_X1 B5zpw6_reg ( .D(Pjshu6), .CK(HCLK), .Q(vis_psp_o[4]), .QN(n4278) );
  DFF_X1 B0spw6_reg ( .D(Vfshu6), .CK(HCLK), .Q(vis_r0_o[6]), .QN(n6294) );
  DFF_X1 A2spw6_reg ( .D(Cgshu6), .CK(HCLK), .Q(vis_r1_o[6]), .QN(n6863) );
  DFF_X1 V1yax6_reg ( .D(Ibthu6), .CK(HCLK), .Q(vis_r3_o[0]), .QN(n7578) );
  DFF_X1 S5nax6_reg ( .D(O0thu6), .CK(HCLK), .Q(vis_r14_o[0]), .QN(n8088) );
  DFF_X1 Rtvax6_reg ( .D(W4thu6), .CK(HCLK), .Q(vis_r7_o[0]), .QN(n7760) );
  DFF_X1 Qukax6_reg ( .D(Cushu6), .CK(HCLK), .Q(vis_r9_o[0]), .QN(n6175) );
  DFF_X1 Qorax6_reg ( .D(Prrhu6), .CK(HCLK), .Q(vis_r8_o[0]), .QN(n5851) );
  DFF_X1 Pwkax6_reg ( .D(Ixshu6), .CK(HCLK), .Q(vis_r11_o[0]), .QN(n8127) );
  DFF_X1 Oykax6_reg ( .D(C8thu6), .CK(HCLK), .Q(vis_r5_o[0]), .QN(n3343) );
  DFF_X1 N0lax6_reg ( .D(Eevhu6), .CK(HCLK), .Q(vis_r0_o[0]), .QN(n6378) );
  DFF_X1 M2lax6_reg ( .D(Sevhu6), .CK(HCLK), .Q(vis_r1_o[0]), .QN(n6628) );
  DFF_X1 Kssax6_reg ( .D(Yyshu6), .CK(HCLK), .Q(vis_r12_o[0]), .QN(n6176) );
  DFF_X1 Kloax6_reg ( .D(M6thu6), .CK(HCLK), .Q(vis_r6_o[0]), .QN(n5730) );
  DFF_X1 Cmlax6_reg ( .D(Svshu6), .CK(HCLK), .Q(vis_r10_o[0]), .QN(n8055) );
  DFF_X1 Bauax6_reg ( .D(S9thu6), .CK(HCLK), .Q(vis_r4_o[0]), .QN(n5366) );
  DFF_X1 A5qax6_reg ( .D(Ycthu6), .CK(HCLK), .Q(vis_r2_o[0]), .QN(n5468) );
  DFF_X1 Gxmpw6_reg ( .D(Gpshu6), .CK(HCLK), .Q(vis_r0_o[3]), .QN(n6365) );
  DFF_X1 X3max6_reg ( .D(Xorhu6), .CK(HCLK), .Q(vis_r10_o[1]), .QN(n7922) );
  DFF_X1 Wruax6_reg ( .D(Lprhu6), .CK(HCLK), .Q(vis_r4_o[1]), .QN(n5403) );
  DFF_X1 Vmqax6_reg ( .D(Vnrhu6), .CK(HCLK), .Q(vis_r2_o[1]), .QN(n5484) );
  DFF_X1 Tdypw6_reg ( .D(Hnrhu6), .CK(HCLK), .Q(vis_r0_o[1]), .QN(n6351) );
  DFF_X1 Sfypw6_reg ( .D(Onrhu6), .CK(HCLK), .Q(vis_r1_o[1]), .QN(n6642) );
  DFF_X1 Rhypw6_reg ( .D(Qorhu6), .CK(HCLK), .Q(vis_r9_o[1]), .QN(n6121) );
  DFF_X1 Qjypw6_reg ( .D(Eprhu6), .CK(HCLK), .Q(vis_r11_o[1]), .QN(n8129) );
  DFF_X1 Pqrax6_reg ( .D(Jorhu6), .CK(HCLK), .Q(vis_r8_o[1]), .QN(n5876) );
  DFF_X1 Plypw6_reg ( .D(Sprhu6), .CK(HCLK), .Q(vis_r5_o[1]), .QN(n6479) );
  DFF_X1 Onypw6_reg ( .D(Uqrhu6), .CK(HCLK), .Q(vis_r14_o[1]), .QN(n8078) );
  DFF_X1 Nq5bx6_reg ( .D(Corhu6), .CK(HCLK), .Q(vis_r3_o[1]), .QN(n4352) );
  DFF_X1 Mbwax6_reg ( .D(Gqrhu6), .CK(HCLK), .Q(vis_r7_o[1]), .QN(n7800) );
  DFF_X1 Fatax6_reg ( .D(Nqrhu6), .CK(HCLK), .Q(vis_r12_o[1]), .QN(n6219) );
  DFF_X1 F3pax6_reg ( .D(Zprhu6), .CK(HCLK), .Q(vis_r6_o[1]), .QN(n5642) );
  DFF_X1 Z6qax6_reg ( .D(Upshu6), .CK(HCLK), .Q(vis_r2_o[3]), .QN(n5506) );
  DFF_X1 Xozpw6_reg ( .D(Tsshu6), .CK(HCLK), .Q(vis_msp_o[1]), .QN(n5928) );
  DFF_X1 U3yax6_reg ( .D(Bqshu6), .CK(HCLK), .Q(vis_r3_o[3]), .QN(n7668) );
  DFF_X1 R7nax6_reg ( .D(Msshu6), .CK(HCLK), .Q(vis_r14_o[3]), .QN(n8090) );
  DFF_X1 Qvvax6_reg ( .D(Yrshu6), .CK(HCLK), .Q(vis_r7_o[3]), .QN(n7748) );
  DFF_X1 Qpopw6_reg ( .D(Iqshu6), .CK(HCLK), .Q(vis_r9_o[3]), .QN(n6151) );
  DFF_X1 Qbmpw6_reg ( .D(Wqshu6), .CK(HCLK), .Q(vis_r11_o[3]), .QN(n8110) );
  DFF_X1 Pdmpw6_reg ( .D(Otshu6), .CK(HCLK), .Q(vis_r8_o[3]), .QN(n5865) );
  DFF_X1 Nbppw6_reg ( .D(Krshu6), .CK(HCLK), .Q(vis_r5_o[3]), .QN(n6570) );
  DFF_X1 Ktppw6_reg ( .D(Npshu6), .CK(HCLK), .Q(vis_r1_o[3]), .QN(n6657) );
  DFF_X1 Jusax6_reg ( .D(Fsshu6), .CK(HCLK), .Q(vis_r12_o[3]), .QN(n6260) );
  DFF_X1 Jnoax6_reg ( .D(Rrshu6), .CK(HCLK), .Q(vis_r6_o[3]), .QN(n5710) );
  DFF_X1 D1zpw6_reg ( .D(Atshu6), .CK(HCLK), .Q(vis_psp_o[1]), .QN(n3774) );
  DFF_X1 Bolax6_reg ( .D(Pqshu6), .CK(HCLK), .Q(vis_r10_o[3]), .QN(n8060) );
  DFF_X1 Acuax6_reg ( .D(Drshu6), .CK(HCLK), .Q(vis_r4_o[3]), .QN(n5461) );
  DFF_X1 Tu0qw6_reg ( .D(Nlphu6), .CK(HCLK), .Q(vis_r0_o[8]), .QN(n6329) );
  DFF_X1 Hkxpw6_reg ( .D(Yuphu6), .CK(HCLK), .Q(vis_r0_o[10]), .QN(n6281) );
  DFF_X1 Ebnpw6_reg ( .D(C4qhu6), .CK(HCLK), .Q(vis_r0_o[12]), .QN(n6387) );
  DFF_X1 C27bx6_reg ( .D(Nzphu6), .CK(HCLK), .Q(vis_r0_o[11]), .QN(n6328) );
  DFF_X1 Emrpw6_reg ( .D(Gbshu6), .CK(HCLK), .Q(vis_r0_o[7]), .QN(n6377) );
  DFF_X1 Vltpw6_reg ( .D(B9vhu6), .CK(HCLK), .Q(vis_r0_o[2]), .QN(n4273) );
  DFF_X1 Uwipw6_reg ( .D(Igvhu6), .CK(HCLK), .Q(vis_r0_o[4]), .QN(n6349) );
  DFF_X1 E9npw6_reg ( .D(R8qhu6), .CK(HCLK), .Q(vis_r0_o[13]), .QN(n6317) );
  DFF_X1 Sx7ax6_reg ( .D(Gdqhu6), .CK(HCLK), .Q(vis_r0_o[14]), .QN(n6372) );
  DFF_X1 Wpmax6_reg ( .D(Owphu6), .CK(HCLK), .Q(vis_r10_o[10]), .QN(n8062) );
  DFF_X1 Vtmax6_reg ( .D(Dnphu6), .CK(HCLK), .Q(vis_r10_o[8]), .QN(n8072) );
  DFF_X1 Vdvax6_reg ( .D(Cxphu6), .CK(HCLK), .Q(vis_r4_o[10]), .QN(n5463) );
  DFF_X1 Uhvax6_reg ( .D(Rnphu6), .CK(HCLK), .Q(vis_r4_o[8]), .QN(n5370) );
  DFF_X1 U8rax6_reg ( .D(Mvphu6), .CK(HCLK), .Q(vis_r2_o[10]), .QN(n5534) );
  DFF_X1 Tm0qw6_reg ( .D(Syphu6), .CK(HCLK), .Q(vis_msp_o[8]), .QN(n5938) );
  DFF_X1 Tcrax6_reg ( .D(Bmphu6), .CK(HCLK), .Q(vis_r2_o[8]), .QN(n5598) );
  DFF_X1 Sw0qw6_reg ( .D(Ulphu6), .CK(HCLK), .Q(vis_r1_o[8]), .QN(n6626) );
  DFF_X1 So0qw6_reg ( .D(Hpphu6), .CK(HCLK), .Q(vis_msp_o[6]), .QN(n5963) );
  DFF_X1 Ry0qw6_reg ( .D(Wmphu6), .CK(HCLK), .Q(vis_r9_o[8]), .QN(n6104) );
  DFF_X1 Q01qw6_reg ( .D(Knphu6), .CK(HCLK), .Q(vis_r11_o[8]), .QN(n8125) );
  DFF_X1 P21qw6_reg ( .D(Ynphu6), .CK(HCLK), .Q(vis_r5_o[8]), .QN(n6399) );
  DFF_X1 Ocsax6_reg ( .D(Awphu6), .CK(HCLK), .Q(vis_r8_o[10]), .QN(n3614) );
  DFF_X1 O41qw6_reg ( .D(Opphu6), .CK(HCLK), .Q(vis_psp_o[6]), .QN(n4007) );
  DFF_X1 Ngsax6_reg ( .D(Pmphu6), .CK(HCLK), .Q(vis_r8_o[8]), .QN(n5859) );
  DFF_X1 N9oax6_reg ( .D(Apphu6), .CK(HCLK), .Q(vis_r14_o[8]), .QN(n4008) );
  DFF_X1 N7oax6_reg ( .D(Lyphu6), .CK(HCLK), .Q(vis_r14_o[10]), .QN(n8093) );
  DFF_X1 Lzwax6_reg ( .D(Mophu6), .CK(HCLK), .Q(vis_r7_o[8]), .QN(n7787) );
  DFF_X1 Lxwax6_reg ( .D(Xxphu6), .CK(HCLK), .Q(vis_r7_o[10]), .QN(n7757) );
  DFF_X1 Huxpw6_reg ( .D(Zyphu6), .CK(HCLK), .Q(vis_psp_o[8]), .QN(n3611) );
  DFF_X1 Hsxpw6_reg ( .D(Jxphu6), .CK(HCLK), .Q(vis_r5_o[10]), .QN(n6574) );
  DFF_X1 Hqxpw6_reg ( .D(Vwphu6), .CK(HCLK), .Q(vis_r11_o[10]), .QN(n8113) );
  DFF_X1 Hoxpw6_reg ( .D(Hwphu6), .CK(HCLK), .Q(vis_r9_o[10]), .QN(n6153) );
  DFF_X1 Hmxpw6_reg ( .D(Fvphu6), .CK(HCLK), .Q(vis_r1_o[10]), .QN(n6810) );
  DFF_X1 Eytax6_reg ( .D(Tophu6), .CK(HCLK), .Q(vis_r12_o[8]), .QN(n6210) );
  DFF_X1 Ewtax6_reg ( .D(Eyphu6), .CK(HCLK), .Q(vis_r12_o[10]), .QN(n6267) );
  DFF_X1 Eppax6_reg ( .D(Qxphu6), .CK(HCLK), .Q(vis_r6_o[10]), .QN(n5718) );
  DFF_X1 Dtpax6_reg ( .D(Fophu6), .CK(HCLK), .Q(vis_r6_o[8]), .QN(n5799) );
  DFF_X1 Do6bx6_reg ( .D(Tvphu6), .CK(HCLK), .Q(vis_r3_o[10]), .QN(n7307) );
  DFF_X1 Cs6bx6_reg ( .D(Imphu6), .CK(HCLK), .Q(vis_r3_o[8]), .QN(n7577) );
  DFF_X1 Wnmax6_reg ( .D(S5qhu6), .CK(HCLK), .Q(vis_r10_o[12]), .QN(n8057) );
  DFF_X1 Vbvax6_reg ( .D(G6qhu6), .CK(HCLK), .Q(vis_r4_o[12]), .QN(n5449) );
  DFF_X1 U6rax6_reg ( .D(Q4qhu6), .CK(HCLK), .Q(vis_r2_o[12]), .QN(n5526) );
  DFF_X1 Tk0qw6_reg ( .D(W7qhu6), .CK(HCLK), .Q(vis_msp_o[10]), .QN(n5915) );
  DFF_X1 Oasax6_reg ( .D(E5qhu6), .CK(HCLK), .Q(vis_r8_o[12]), .QN(n5892) );
  DFF_X1 O3ppw6_reg ( .D(L5qhu6), .CK(HCLK), .Q(vis_r9_o[12]), .QN(n6144) );
  DFF_X1 N5oax6_reg ( .D(P7qhu6), .CK(HCLK), .Q(vis_r14_o[12]), .QN(n8087) );
  DFF_X1 Lvwax6_reg ( .D(B7qhu6), .CK(HCLK), .Q(vis_r7_o[12]), .QN(n4179) );
  DFF_X1 Lpppw6_reg ( .D(N6qhu6), .CK(HCLK), .Q(vis_r5_o[12]), .QN(n6526) );
  DFF_X1 I7qpw6_reg ( .D(J4qhu6), .CK(HCLK), .Q(vis_r1_o[12]), .QN(n6678) );
  DFF_X1 Eutax6_reg ( .D(I7qhu6), .CK(HCLK), .Q(vis_r12_o[12]), .QN(n6242) );
  DFF_X1 Enpax6_reg ( .D(U6qhu6), .CK(HCLK), .Q(vis_r6_o[12]), .QN(n5683) );
  DFF_X1 Dk6bx6_reg ( .D(X4qhu6), .CK(HCLK), .Q(vis_r3_o[12]), .QN(n6899) );
  DFF_X1 Bdjpw6_reg ( .D(D8qhu6), .CK(HCLK), .Q(vis_psp_o[10]), .QN(n4178) );
  DFF_X1 Bbjpw6_reg ( .D(Z5qhu6), .CK(HCLK), .Q(vis_r11_o[12]), .QN(n8102) );
  DFF_X1 Zr8bx6_reg ( .D(H3qhu6), .CK(HCLK), .Q(vis_msp_o[9]), .QN(n5964) );
  DFF_X1 Zp8bx6_reg ( .D(A3qhu6), .CK(HCLK), .Q(vis_r14_o[11]), .QN(n2816) );
  DFF_X1 Zn8bx6_reg ( .D(T2qhu6), .CK(HCLK), .Q(vis_r12_o[11]), .QN(n6212) );
  DFF_X1 Yt8bx6_reg ( .D(O3qhu6), .CK(HCLK), .Q(vis_psp_o[9]), .QN(n3591) );
  DFF_X1 Co7bx6_reg ( .D(M2qhu6), .CK(HCLK), .Q(vis_r7_o[11]), .QN(n7790) );
  DFF_X1 Cm7bx6_reg ( .D(F2qhu6), .CK(HCLK), .Q(vis_r6_o[11]), .QN(n5802) );
  DFF_X1 Ck7bx6_reg ( .D(Y1qhu6), .CK(HCLK), .Q(vis_r5_o[11]), .QN(n6425) );
  DFF_X1 Ci7bx6_reg ( .D(R1qhu6), .CK(HCLK), .Q(vis_r4_o[11]), .QN(n5372) );
  DFF_X1 Cg7bx6_reg ( .D(K1qhu6), .CK(HCLK), .Q(vis_r11_o[11]), .QN(n8126) );
  DFF_X1 Ce7bx6_reg ( .D(D1qhu6), .CK(HCLK), .Q(vis_r10_o[11]), .QN(n8073) );
  DFF_X1 Cc7bx6_reg ( .D(W0qhu6), .CK(HCLK), .Q(vis_r9_o[11]), .QN(n6105) );
  DFF_X1 Ca7bx6_reg ( .D(P0qhu6), .CK(HCLK), .Q(vis_r8_o[11]), .QN(n5860) );
  DFF_X1 C87bx6_reg ( .D(I0qhu6), .CK(HCLK), .Q(vis_r3_o[11]), .QN(n7579) );
  DFF_X1 C67bx6_reg ( .D(B0qhu6), .CK(HCLK), .Q(vis_r2_o[11]), .QN(n5606) );
  DFF_X1 C47bx6_reg ( .D(Uzphu6), .CK(HCLK), .Q(vis_r1_o[11]), .QN(n6607) );
  DFF_X1 Zvrpw6_reg ( .D(Ofshu6), .CK(HCLK), .Q(vis_r8_o[7]), .QN(n5872) );
  DFF_X1 Ytlax6_reg ( .D(Pcshu6), .CK(HCLK), .Q(vis_r10_o[7]), .QN(n8061) );
  DFF_X1 Xhuax6_reg ( .D(Ddshu6), .CK(HCLK), .Q(vis_r4_o[7]), .QN(n5462) );
  DFF_X1 Wcqax6_reg ( .D(Ubshu6), .CK(HCLK), .Q(vis_r2_o[7]), .QN(n5520) );
  DFF_X1 Uuzpw6_reg ( .D(Teshu6), .CK(HCLK), .Q(vis_msp_o[5]), .QN(n5935) );
  DFF_X1 Og5bx6_reg ( .D(Bcshu6), .CK(HCLK), .Q(vis_r3_o[7]), .QN(n7695) );
  DFF_X1 Odnax6_reg ( .D(Meshu6), .CK(HCLK), .Q(vis_r14_o[7]), .QN(n8091) );
  DFF_X1 N1wax6_reg ( .D(Ydshu6), .CK(HCLK), .Q(vis_r7_o[7]), .QN(n7751) );
  DFF_X1 Gtoax6_reg ( .D(Rdshu6), .CK(HCLK), .Q(vis_r6_o[7]), .QN(n5711) );
  DFF_X1 G0tax6_reg ( .D(Feshu6), .CK(HCLK), .Q(vis_r12_o[7]), .QN(n6264) );
  DFF_X1 Dorpw6_reg ( .D(Nbshu6), .CK(HCLK), .Q(vis_r1_o[7]), .QN(n6668) );
  DFF_X1 Cqrpw6_reg ( .D(Icshu6), .CK(HCLK), .Q(vis_r9_o[7]), .QN(n6152) );
  DFF_X1 Bsrpw6_reg ( .D(Wcshu6), .CK(HCLK), .Q(vis_r11_o[7]), .QN(n8112) );
  DFF_X1 Aurpw6_reg ( .D(Kdshu6), .CK(HCLK), .Q(vis_r5_o[7]), .QN(n6571) );
  DFF_X1 A7zpw6_reg ( .D(Afshu6), .CK(HCLK), .Q(vis_psp_o[5]), .QN(n4181) );
  DFF_X1 Zgzpw6_reg ( .D(G3thu6), .CK(HCLK), .Q(vis_msp_o[0]), .QN(n5976) );
  DFF_X1 Yftpw6_reg ( .D(Lvshu6), .CK(HCLK), .Q(vis_r9_o[2]), .QN(n6138) );
  DFF_X1 Xhtpw6_reg ( .D(Ryshu6), .CK(HCLK), .Q(vis_r11_o[2]), .QN(n8117) );
  DFF_X1 Wjtpw6_reg ( .D(L9thu6), .CK(HCLK), .Q(vis_r5_o[2]), .QN(n6537) );
  DFF_X1 Uvmax6_reg ( .D(X1thu6), .CK(HCLK), .Q(vis_r14_o[2]), .QN(n8076) );
  DFF_X1 Untpw6_reg ( .D(I9vhu6), .CK(HCLK), .Q(vis_r1_o[2]), .QN(n6686) );
  DFF_X1 Tjvax6_reg ( .D(F6thu6), .CK(HCLK), .Q(vis_r7_o[2]), .QN(n7809) );
  DFF_X1 Serax6_reg ( .D(Vtshu6), .CK(HCLK), .Q(vis_r8_o[2]), .QN(n5832) );
  DFF_X1 Misax6_reg ( .D(H0thu6), .CK(HCLK), .Q(vis_r12_o[2]), .QN(n6249) );
  DFF_X1 Mboax6_reg ( .D(V7thu6), .CK(HCLK), .Q(vis_r6_o[2]), .QN(n5673) );
  DFF_X1 K1xax6_reg ( .D(Rcthu6), .CK(HCLK), .Q(vis_r3_o[2]), .QN(n7370) );
  DFF_X1 Ftypw6_reg ( .D(P4thu6), .CK(HCLK), .Q(vis_psp_o[0]), .QN(n4272) );
  DFF_X1 Eclax6_reg ( .D(Bxshu6), .CK(HCLK), .Q(vis_r10_o[2]), .QN(n8074) );
  DFF_X1 D0uax6_reg ( .D(Bbthu6), .CK(HCLK), .Q(vis_r4_o[2]), .QN(n5464) );
  DFF_X1 Cvpax6_reg ( .D(Hethu6), .CK(HCLK), .Q(vis_r2_o[2]), .QN(n5562) );
  DFF_X1 Ymzpw6_reg ( .D(E2thu6), .CK(HCLK), .Q(vis_msp_o[2]), .QN(n5990) );
  DFF_X1 Vuipw6_reg ( .D(Kyshu6), .CK(HCLK), .Q(vis_r11_o[4]), .QN(n8124) );
  DFF_X1 Txmax6_reg ( .D(Q1thu6), .CK(HCLK), .Q(vis_r14_o[4]), .QN(n8085) );
  DFF_X1 Slvax6_reg ( .D(Y5thu6), .CK(HCLK), .Q(vis_r7_o[4]), .QN(n7754) );
  DFF_X1 Rjopw6_reg ( .D(Evshu6), .CK(HCLK), .Q(vis_r9_o[4]), .QN(n6167) );
  DFF_X1 Rgrax6_reg ( .D(Zoshu6), .CK(HCLK), .Q(vis_r8_o[4]), .QN(n5814) );
  DFF_X1 O5ppw6_reg ( .D(E9thu6), .CK(HCLK), .Q(vis_r5_o[4]), .QN(n6586) );
  DFF_X1 Lrppw6_reg ( .D(Zevhu6), .CK(HCLK), .Q(vis_r1_o[4]), .QN(n6600) );
  DFF_X1 Lksax6_reg ( .D(A0thu6), .CK(HCLK), .Q(vis_r12_o[4]), .QN(n2777) );
  DFF_X1 Ldoax6_reg ( .D(O7thu6), .CK(HCLK), .Q(vis_r6_o[4]), .QN(n5726) );
  DFF_X1 J3xax6_reg ( .D(Kcthu6), .CK(HCLK), .Q(vis_r3_o[4]), .QN(n7575) );
  DFF_X1 Ezypw6_reg ( .D(N3thu6), .CK(HCLK), .Q(vis_psp_o[2]), .QN(n3592) );
  DFF_X1 Delax6_reg ( .D(Uwshu6), .CK(HCLK), .Q(vis_r10_o[4]), .QN(n8019) );
  DFF_X1 C2uax6_reg ( .D(Uathu6), .CK(HCLK), .Q(vis_r4_o[4]), .QN(n5348) );
  DFF_X1 Bxpax6_reg ( .D(Aethu6), .CK(HCLK), .Q(vis_r2_o[4]), .QN(n5624) );
  DFF_X1 Wlmax6_reg ( .D(Haqhu6), .CK(HCLK), .Q(vis_r10_o[13]), .QN(n8068) );
  DFF_X1 Vnkpw6_reg ( .D(Scqhu6), .CK(HCLK), .Q(vis_psp_o[11]), .QN(n3588) );
  DFF_X1 Vlkpw6_reg ( .D(Oaqhu6), .CK(HCLK), .Q(vis_r11_o[13]), .QN(n8121) );
  DFF_X1 V9vax6_reg ( .D(Vaqhu6), .CK(HCLK), .Q(vis_r4_o[13]), .QN(n5334) );
  DFF_X1 U4rax6_reg ( .D(F9qhu6), .CK(HCLK), .Q(vis_r2_o[13]), .QN(n5584) );
  DFF_X1 Ti0qw6_reg ( .D(Lcqhu6), .CK(HCLK), .Q(vis_msp_o[11]), .QN(n5956) );
  DFF_X1 O8sax6_reg ( .D(T9qhu6), .CK(HCLK), .Q(vis_r8_o[13]), .QN(n5839) );
  DFF_X1 O1ppw6_reg ( .D(Aaqhu6), .CK(HCLK), .Q(vis_r9_o[13]), .QN(n3039) );
  DFF_X1 N3oax6_reg ( .D(Ecqhu6), .CK(HCLK), .Q(vis_r14_o[13]), .QN(n8099) );
  DFF_X1 Ltwax6_reg ( .D(Qbqhu6), .CK(HCLK), .Q(vis_r7_o[13]), .QN(n7778) );
  DFF_X1 Lnppw6_reg ( .D(Cbqhu6), .CK(HCLK), .Q(vis_r5_o[13]), .QN(n6595) );
  DFF_X1 I5qpw6_reg ( .D(Y8qhu6), .CK(HCLK), .Q(vis_r1_o[13]), .QN(n6603) );
  DFF_X1 Estax6_reg ( .D(Xbqhu6), .CK(HCLK), .Q(vis_r12_o[13]), .QN(n6183) );
  DFF_X1 Elpax6_reg ( .D(Jbqhu6), .CK(HCLK), .Q(vis_r6_o[13]), .QN(n5752) );
  DFF_X1 Di6bx6_reg ( .D(M9qhu6), .CK(HCLK), .Q(vis_r3_o[13]), .QN(n7573) );
  DFF_X1 Wjmax6_reg ( .D(Weqhu6), .CK(HCLK), .Q(vis_r10_o[14]), .QN(n8018) );
  DFF_X1 V7vax6_reg ( .D(Kfqhu6), .CK(HCLK), .Q(vis_r4_o[14]), .QN(n5410) );
  DFF_X1 U2rax6_reg ( .D(Udqhu6), .CK(HCLK), .Q(vis_r2_o[14]), .QN(n5507) );
  DFF_X1 Sz7ax6_reg ( .D(Ndqhu6), .CK(HCLK), .Q(vis_r1_o[14]), .QN(n6663) );
  DFF_X1 S98ax6_reg ( .D(Hhqhu6), .CK(HCLK), .Q(vis_psp_o[12]), .QN(n4167) );
  DFF_X1 S78ax6_reg ( .D(Ahqhu6), .CK(HCLK), .Q(vis_msp_o[12]), .QN(n8251) );
  DFF_X1 S58ax6_reg ( .D(Rfqhu6), .CK(HCLK), .Q(vis_r5_o[14]), .QN(n6484) );
  DFF_X1 S38ax6_reg ( .D(Dfqhu6), .CK(HCLK), .Q(vis_r11_o[14]), .QN(n8132) );
  DFF_X1 S18ax6_reg ( .D(Peqhu6), .CK(HCLK), .Q(vis_r9_o[14]), .QN(n6124) );
  DFF_X1 O6sax6_reg ( .D(Ieqhu6), .CK(HCLK), .Q(vis_r8_o[14]), .QN(n5886) );
  DFF_X1 N1oax6_reg ( .D(Tgqhu6), .CK(HCLK), .Q(vis_r14_o[14]), .QN(n8080) );
  DFF_X1 Lrwax6_reg ( .D(Fgqhu6), .CK(HCLK), .Q(vis_r7_o[14]), .QN(n7806) );
  DFF_X1 Eqtax6_reg ( .D(Mgqhu6), .CK(HCLK), .Q(vis_r12_o[14]), .QN(n6225) );
  DFF_X1 Ejpax6_reg ( .D(Yfqhu6), .CK(HCLK), .Q(vis_r6_o[14]), .QN(n5662) );
  DFF_X1 Dg6bx6_reg ( .D(Beqhu6), .CK(HCLK), .Q(vis_r3_o[14]), .QN(n4170) );
  DFF_X1 Fzmpw6_reg ( .D(Kkshu6), .CK(HCLK), .Q(vis_r0_o[5]), .QN(n6331) );
  DFF_X1 Zduax6_reg ( .D(Hmshu6), .CK(HCLK), .Q(vis_r4_o[5]), .QN(n5411) );
  DFF_X1 Y8qax6_reg ( .D(Ykshu6), .CK(HCLK), .Q(vis_r2_o[5]), .QN(n5467) );
  DFF_X1 Wqzpw6_reg ( .D(Xnshu6), .CK(HCLK), .Q(vis_msp_o[3]), .QN(n5899) );
  DFF_X1 T3kpw6_reg ( .D(Amshu6), .CK(HCLK), .Q(vis_r11_o[5]), .QN(n4109) );
  DFF_X1 S7yax6_reg ( .D(Flshu6), .CK(HCLK), .Q(vis_r3_o[5]), .QN(n7600) );
  DFF_X1 S5kpw6_reg ( .D(Soshu6), .CK(HCLK), .Q(vis_r8_o[5]), .QN(n5846) );
  DFF_X1 Q9nax6_reg ( .D(Qnshu6), .CK(HCLK), .Q(vis_r14_o[5]), .QN(n8081) );
  DFF_X1 Pxvax6_reg ( .D(Cnshu6), .CK(HCLK), .Q(vis_r7_o[5]), .QN(n7815) );
  DFF_X1 Propw6_reg ( .D(Mlshu6), .CK(HCLK), .Q(vis_r9_o[5]), .QN(n6128) );
  DFF_X1 Mdppw6_reg ( .D(Omshu6), .CK(HCLK), .Q(vis_r5_o[5]), .QN(n6487) );
  DFF_X1 Jvppw6_reg ( .D(Rkshu6), .CK(HCLK), .Q(vis_r1_o[5]), .QN(n6638) );
  DFF_X1 Iwsax6_reg ( .D(Jnshu6), .CK(HCLK), .Q(vis_r12_o[5]), .QN(n6229) );
  DFF_X1 Ipoax6_reg ( .D(Vmshu6), .CK(HCLK), .Q(vis_r6_o[5]), .QN(n5663) );
  DFF_X1 C3zpw6_reg ( .D(Eoshu6), .CK(HCLK), .Q(vis_psp_o[3]), .QN(n4086) );
  DFF_X1 Aqlax6_reg ( .D(Tlshu6), .CK(HCLK), .Q(vis_r10_o[5]), .QN(n8036) );
  DFF_X1 Wrmax6_reg ( .D(Srphu6), .CK(HCLK), .Q(vis_r10_o[9]), .QN(n8056) );
  DFF_X1 Vfvax6_reg ( .D(Gsphu6), .CK(HCLK), .Q(vis_r4_o[9]), .QN(n5428) );
  DFF_X1 Uarax6_reg ( .D(Qqphu6), .CK(HCLK), .Q(vis_r2_o[9]), .QN(n5523) );
  DFF_X1 Rvibx6_reg ( .D(Itphu6), .CK(HCLK), .Q(vis_r12_o[9]), .QN(n6241) );
  DFF_X1 Qxibx6_reg ( .D(Ptphu6), .CK(HCLK), .Q(vis_r14_o[9]), .QN(n8086) );
  DFF_X1 Pzibx6_reg ( .D(Wtphu6), .CK(HCLK), .Q(vis_msp_o[7]), .QN(n5914) );
  DFF_X1 Oesax6_reg ( .D(Erphu6), .CK(HCLK), .Q(vis_r8_o[9]), .QN(n5891) );
  DFF_X1 O1jbx6_reg ( .D(Duphu6), .CK(HCLK), .Q(vis_psp_o[7]), .QN(n3598) );
  DFF_X1 Jp1qw6_reg ( .D(Cqphu6), .CK(HCLK), .Q(vis_r0_o[9]), .QN(n6386) );
  DFF_X1 Ir1qw6_reg ( .D(Jqphu6), .CK(HCLK), .Q(vis_r1_o[9]), .QN(n6674) );
  DFF_X1 Ht1qw6_reg ( .D(Lrphu6), .CK(HCLK), .Q(vis_r9_o[9]), .QN(n6142) );
  DFF_X1 Gv1qw6_reg ( .D(Zrphu6), .CK(HCLK), .Q(vis_r11_o[9]), .QN(n8101) );
  DFF_X1 Fx1qw6_reg ( .D(Nsphu6), .CK(HCLK), .Q(vis_r5_o[9]), .QN(n6524) );
  DFF_X1 Ez1qw6_reg ( .D(Btphu6), .CK(HCLK), .Q(vis_r7_o[9]), .QN(n3341) );
  DFF_X1 Erpax6_reg ( .D(Usphu6), .CK(HCLK), .Q(vis_r6_o[9]), .QN(n5682) );
  DFF_X1 Dq6bx6_reg ( .D(Xqphu6), .CK(HCLK), .Q(vis_r3_o[9]), .QN(n6886) );
  DFF_X1 Jjvpw6_reg ( .D(D0rhu6), .CK(HCLK), .Q(vis_r0_o[19]), .QN(n6380) );
  DFF_X1 Wbmax6_reg ( .D(T1rhu6), .CK(HCLK), .Q(vis_r10_o[19]), .QN(n8040) );
  DFF_X1 Vzuax6_reg ( .D(H2rhu6), .CK(HCLK), .Q(vis_r4_o[19]), .QN(n5427) );
  DFF_X1 Uuqax6_reg ( .D(R0rhu6), .CK(HCLK), .Q(vis_r2_o[19]), .QN(n5522) );
  DFF_X1 Ta0qw6_reg ( .D(X3rhu6), .CK(HCLK), .Q(vis_msp_o[17]), .QN(n5905) );
  DFF_X1 Oyrax6_reg ( .D(F1rhu6), .CK(HCLK), .Q(vis_r8_o[19]), .QN(n5887) );
  DFF_X1 Ntnax6_reg ( .D(Q3rhu6), .CK(HCLK), .Q(vis_r14_o[19]), .QN(n8084) );
  DFF_X1 Ljwax6_reg ( .D(C3rhu6), .CK(HCLK), .Q(vis_r7_o[19]), .QN(n7821) );
  DFF_X1 Jtvpw6_reg ( .D(E4rhu6), .CK(HCLK), .Q(vis_psp_o[17]), .QN(n3864) );
  DFF_X1 Jrvpw6_reg ( .D(O2rhu6), .CK(HCLK), .Q(vis_r5_o[19]), .QN(n6518) );
  DFF_X1 Jpvpw6_reg ( .D(A2rhu6), .CK(HCLK), .Q(vis_r11_o[19]), .QN(n3865) );
  DFF_X1 Jnvpw6_reg ( .D(M1rhu6), .CK(HCLK), .Q(vis_r9_o[19]), .QN(n6136) );
  DFF_X1 Jlvpw6_reg ( .D(K0rhu6), .CK(HCLK), .Q(vis_r1_o[19]), .QN(n6669) );
  DFF_X1 Eitax6_reg ( .D(J3rhu6), .CK(HCLK), .Q(vis_r12_o[19]), .QN(n6239) );
  DFF_X1 Ebpax6_reg ( .D(V2rhu6), .CK(HCLK), .Q(vis_r6_o[19]), .QN(n5676) );
  DFF_X1 D86bx6_reg ( .D(Y0rhu6), .CK(HCLK), .Q(vis_r3_o[19]), .QN(n6871) );
  DFF_X1 Nwbbx6_reg ( .D(n7753), .CK(HCLK), .Q(n6680), .QN(n3335) );
  DFF_X1 E7npw6_reg ( .D(S4rhu6), .CK(HCLK), .Q(vis_r0_o[20]), .QN(n8212) );
  DFF_X1 X4jpw6_reg ( .D(T8rhu6), .CK(HCLK), .Q(vis_psp_o[18]), .QN(n8211) );
  DFF_X1 X2jpw6_reg ( .D(P6rhu6), .CK(HCLK), .Q(vis_r11_o[20]), .QN(n8214) );
  DFF_X1 W9max6_reg ( .D(I6rhu6), .CK(HCLK), .Q(vis_r10_o[20]), .QN(n8218) );
  DFF_X1 Vxuax6_reg ( .D(W6rhu6), .CK(HCLK), .Q(vis_r4_o[20]), .QN(n8209) );
  DFF_X1 Usqax6_reg ( .D(G5rhu6), .CK(HCLK), .Q(vis_r2_o[20]), .QN(n8219) );
  DFF_X1 T80qw6_reg ( .D(M8rhu6), .CK(HCLK), .Q(vis_msp_o[18]), .QN(n8216) );
  DFF_X1 Ozopw6_reg ( .D(B6rhu6), .CK(HCLK), .Q(vis_r9_o[20]), .QN(n8222) );
  DFF_X1 Owrax6_reg ( .D(U5rhu6), .CK(HCLK), .Q(vis_r8_o[20]), .QN(n8210) );
  DFF_X1 Nrnax6_reg ( .D(F8rhu6), .CK(HCLK), .Q(vis_r14_o[20]), .QN(n8220) );
  DFF_X1 Llppw6_reg ( .D(D7rhu6), .CK(HCLK), .Q(vis_r5_o[20]), .QN(n8221) );
  DFF_X1 Lhwax6_reg ( .D(R7rhu6), .CK(HCLK), .Q(vis_r7_o[20]), .QN(n8213) );
  DFF_X1 I3qpw6_reg ( .D(Z4rhu6), .CK(HCLK), .Q(vis_r1_o[20]), .QN(n8207) );
  DFF_X1 Egtax6_reg ( .D(Y7rhu6), .CK(HCLK), .Q(vis_r12_o[20]), .QN(n8208) );
  DFF_X1 E9pax6_reg ( .D(K7rhu6), .CK(HCLK), .Q(vis_r6_o[20]), .QN(n8217) );
  DFF_X1 D66bx6_reg ( .D(N5rhu6), .CK(HCLK), .Q(vis_r3_o[20]), .QN(n8215) );
  DFF_X1 W7max6_reg ( .D(Xarhu6), .CK(HCLK), .Q(vis_r10_o[21]), .QN(n8008) );
  DFF_X1 Vvuax6_reg ( .D(Lbrhu6), .CK(HCLK), .Q(vis_r4_o[21]), .QN(n5409) );
  DFF_X1 Uqqax6_reg ( .D(V9rhu6), .CK(HCLK), .Q(vis_r2_o[21]), .QN(n5485) );
  DFF_X1 T60qw6_reg ( .D(Bdrhu6), .CK(HCLK), .Q(vis_msp_o[19]), .QN(n3653) );
  DFF_X1 Rfkpw6_reg ( .D(Idrhu6), .CK(HCLK), .Q(vis_psp_o[19]), .QN(n3650) );
  DFF_X1 Rdkpw6_reg ( .D(Ebrhu6), .CK(HCLK), .Q(vis_r11_o[21]), .QN(n8130) );
  DFF_X1 Oxopw6_reg ( .D(Qarhu6), .CK(HCLK), .Q(vis_r9_o[21]), .QN(n6122) );
  DFF_X1 Ourax6_reg ( .D(Jarhu6), .CK(HCLK), .Q(vis_r8_o[21]), .QN(n5877) );
  DFF_X1 Npnax6_reg ( .D(Ucrhu6), .CK(HCLK), .Q(vis_r14_o[21]), .QN(n8079) );
  DFF_X1 Ljppw6_reg ( .D(Sbrhu6), .CK(HCLK), .Q(vis_r5_o[21]), .QN(n6480) );
  DFF_X1 Lfwax6_reg ( .D(Gcrhu6), .CK(HCLK), .Q(vis_r7_o[21]), .QN(n7802) );
  DFF_X1 I1qpw6_reg ( .D(O9rhu6), .CK(HCLK), .Q(vis_r1_o[21]), .QN(n6646) );
  DFF_X1 Eetax6_reg ( .D(Ncrhu6), .CK(HCLK), .Q(vis_r12_o[21]), .QN(n6220) );
  DFF_X1 E7pax6_reg ( .D(Zbrhu6), .CK(HCLK), .Q(vis_r6_o[21]), .QN(n5654) );
  DFF_X1 E5npw6_reg ( .D(H9rhu6), .CK(HCLK), .Q(vis_r0_o[21]), .QN(n6352) );
  DFF_X1 D46bx6_reg ( .D(Carhu6), .CK(HCLK), .Q(vis_r3_o[21]), .QN(n7644) );
  DFF_X1 Tnebx6_reg ( .D(Wdrhu6), .CK(HCLK), .Q(vis_r0_o[22]), .QN(n6290) );
  DFF_X1 Tzebx6_reg ( .D(Mfrhu6), .CK(HCLK), .Q(vis_r10_o[22]), .QN(n8064) );
  DFF_X1 Txebx6_reg ( .D(Ffrhu6), .CK(HCLK), .Q(vis_r9_o[22]), .QN(n6156) );
  DFF_X1 Tvebx6_reg ( .D(Yerhu6), .CK(HCLK), .Q(vis_r8_o[22]), .QN(n5822) );
  DFF_X1 Ttebx6_reg ( .D(Rerhu6), .CK(HCLK), .Q(vis_r3_o[22]), .QN(n7342) );
  DFF_X1 Trebx6_reg ( .D(Kerhu6), .CK(HCLK), .Q(vis_r2_o[22]), .QN(n5551) );
  DFF_X1 Tpebx6_reg ( .D(Derhu6), .CK(HCLK), .Q(vis_r1_o[22]), .QN(n6826) );
  DFF_X1 Thfbx6_reg ( .D(Xhrhu6), .CK(HCLK), .Q(vis_psp_o[20]), .QN(n3581) );
  DFF_X1 Tffbx6_reg ( .D(Qhrhu6), .CK(HCLK), .Q(vis_msp_o[20]), .QN(n5940) );
  DFF_X1 Tdfbx6_reg ( .D(Jhrhu6), .CK(HCLK), .Q(vis_r14_o[22]), .QN(n8094) );
  DFF_X1 Tbfbx6_reg ( .D(Chrhu6), .CK(HCLK), .Q(vis_r12_o[22]), .QN(n6271) );
  DFF_X1 T9fbx6_reg ( .D(Vgrhu6), .CK(HCLK), .Q(vis_r7_o[22]), .QN(n7763) );
  DFF_X1 T7fbx6_reg ( .D(Ogrhu6), .CK(HCLK), .Q(vis_r6_o[22]), .QN(n5725) );
  DFF_X1 T5fbx6_reg ( .D(Hgrhu6), .CK(HCLK), .Q(vis_r5_o[22]), .QN(n6583) );
  DFF_X1 T3fbx6_reg ( .D(Agrhu6), .CK(HCLK), .Q(vis_r4_o[22]), .QN(n2727) );
  DFF_X1 T1fbx6_reg ( .D(Tfrhu6), .CK(HCLK), .Q(vis_r11_o[22]), .QN(n8114) );
  DFF_X1 Vvxax6_reg ( .D(Dcthu6), .CK(HCLK), .Q(vis_r3_o[23]), .QN(n7643) );
  DFF_X1 Szmax6_reg ( .D(J1thu6), .CK(HCLK), .Q(vis_r14_o[23]), .QN(n8095) );
  DFF_X1 Rnvax6_reg ( .D(R5thu6), .CK(HCLK), .Q(vis_r7_o[23]), .QN(n7772) );
  DFF_X1 Qirax6_reg ( .D(Zashu6), .CK(HCLK), .Q(vis_r8_o[23]), .QN(n5820) );
  DFF_X1 P54qw6_reg ( .D(Dyshu6), .CK(HCLK), .Q(vis_r11_o[23]), .QN(n8131) );
  DFF_X1 P34qw6_reg ( .D(Xushu6), .CK(HCLK), .Q(vis_r9_o[23]), .QN(n5993) );
  DFF_X1 Kmsax6_reg ( .D(Tzshu6), .CK(HCLK), .Q(vis_r12_o[23]), .QN(n6207) );
  DFF_X1 Kfoax6_reg ( .D(H7thu6), .CK(HCLK), .Q(vis_r6_o[23]), .QN(n5789) );
  DFF_X1 Gx6ax6_reg ( .D(Davhu6), .CK(HCLK), .Q(vis_r1_o[23]), .QN(n3783) );
  DFF_X1 Gv6ax6_reg ( .D(W9vhu6), .CK(HCLK), .Q(vis_r0_o[23]), .QN(n6291) );
  DFF_X1 Gt6ax6_reg ( .D(X8thu6), .CK(HCLK), .Q(vis_r5_o[23]), .QN(n6452) );
  DFF_X1 Gr6ax6_reg ( .D(U3thu6), .CK(HCLK), .Q(vis_psp_o[21]), .QN(n3781) );
  DFF_X1 Gp6ax6_reg ( .D(L2thu6), .CK(HCLK), .Q(vis_msp_o[21]), .QN(n5959) );
  DFF_X1 Cglax6_reg ( .D(Nwshu6), .CK(HCLK), .Q(vis_r10_o[23]), .QN(n8063) );
  DFF_X1 B4uax6_reg ( .D(Nathu6), .CK(HCLK), .Q(vis_r4_o[23]), .QN(n5394) );
  DFF_X1 Azpax6_reg ( .D(Tdthu6), .CK(HCLK), .Q(vis_r2_o[23]), .QN(n5521) );
  DFF_X1 Ynspw6_reg ( .D(K6shu6), .CK(HCLK), .Q(vis_r0_o[24]), .QN(n6341) );
  DFF_X1 Z8zpw6_reg ( .D(Eashu6), .CK(HCLK), .Q(vis_psp_o[22]), .QN(n3596) );
  DFF_X1 Yxspw6_reg ( .D(Sashu6), .CK(HCLK), .Q(vis_r8_o[24]), .QN(n5848) );
  DFF_X1 Yvspw6_reg ( .D(O8shu6), .CK(HCLK), .Q(vis_r5_o[24]), .QN(n6504) );
  DFF_X1 Ytspw6_reg ( .D(A8shu6), .CK(HCLK), .Q(vis_r11_o[24]), .QN(n3482) );
  DFF_X1 Yrspw6_reg ( .D(M7shu6), .CK(HCLK), .Q(vis_r9_o[24]), .QN(n6129) );
  DFF_X1 Ypspw6_reg ( .D(R6shu6), .CK(HCLK), .Q(vis_r1_o[24]), .QN(n6639) );
  DFF_X1 Xvlax6_reg ( .D(T7shu6), .CK(HCLK), .Q(vis_r10_o[24]), .QN(n8038) );
  DFF_X1 Wjuax6_reg ( .D(H8shu6), .CK(HCLK), .Q(vis_r4_o[24]), .QN(n5419) );
  DFF_X1 Veqax6_reg ( .D(Y6shu6), .CK(HCLK), .Q(vis_r2_o[24]), .QN(n5470) );
  DFF_X1 Twzpw6_reg ( .D(X9shu6), .CK(HCLK), .Q(vis_msp_o[22]), .QN(n5901) );
  DFF_X1 Ni5bx6_reg ( .D(F7shu6), .CK(HCLK), .Q(vis_r3_o[24]), .QN(n7603) );
  DFF_X1 Nfnax6_reg ( .D(Q9shu6), .CK(HCLK), .Q(vis_r14_o[24]), .QN(n8083) );
  DFF_X1 M3wax6_reg ( .D(C9shu6), .CK(HCLK), .Q(vis_r7_o[24]), .QN(n7818) );
  DFF_X1 Fvoax6_reg ( .D(V8shu6), .CK(HCLK), .Q(vis_r6_o[24]), .QN(n5669) );
  DFF_X1 F2tax6_reg ( .D(J9shu6), .CK(HCLK), .Q(vis_r12_o[24]), .QN(n6234) );
  DFF_X1 Zbtpw6_reg ( .D(Tmrhu6), .CK(HCLK), .Q(vis_psp_o[23]), .QN(n3586) );
  DFF_X1 Z9tpw6_reg ( .D(Dlrhu6), .CK(HCLK), .Q(vis_r5_o[25]), .QN(n6588) );
  DFF_X1 Z7tpw6_reg ( .D(Pkrhu6), .CK(HCLK), .Q(vis_r11_o[25]), .QN(n8119) );
  DFF_X1 Z5tpw6_reg ( .D(Bkrhu6), .CK(HCLK), .Q(vis_r9_o[25]), .QN(n3324) );
  DFF_X1 Z3tpw6_reg ( .D(Zirhu6), .CK(HCLK), .Q(vis_r1_o[25]), .QN(n6599) );
  DFF_X1 Z1tpw6_reg ( .D(Sirhu6), .CK(HCLK), .Q(vis_r0_o[25]), .QN(n6313) );
  DFF_X1 W5max6_reg ( .D(Ikrhu6), .CK(HCLK), .Q(vis_r10_o[25]), .QN(n8066) );
  DFF_X1 Vtuax6_reg ( .D(Wkrhu6), .CK(HCLK), .Q(vis_r4_o[25]), .QN(n5326) );
  DFF_X1 Uoqax6_reg ( .D(Gjrhu6), .CK(HCLK), .Q(vis_r2_o[25]), .QN(n5579) );
  DFF_X1 T40qw6_reg ( .D(Mmrhu6), .CK(HCLK), .Q(vis_msp_o[23]), .QN(n5948) );
  DFF_X1 Osrax6_reg ( .D(Ujrhu6), .CK(HCLK), .Q(vis_r8_o[25]), .QN(n5834) );
  DFF_X1 Nnnax6_reg ( .D(Fmrhu6), .CK(HCLK), .Q(vis_r14_o[25]), .QN(n8097) );
  DFF_X1 Ldwax6_reg ( .D(Rlrhu6), .CK(HCLK), .Q(vis_r7_o[25]), .QN(n7769) );
  DFF_X1 Jy5bx6_reg ( .D(Njrhu6), .CK(HCLK), .Q(vis_r3_o[25]), .QN(n7571) );
  DFF_X1 Ectax6_reg ( .D(Ylrhu6), .CK(HCLK), .Q(vis_r12_o[25]), .QN(n6177) );
  DFF_X1 E5pax6_reg ( .D(Klrhu6), .CK(HCLK), .Q(vis_r6_o[25]), .QN(n5736) );
  DFF_X1 Xttpw6_reg ( .D(V1shu6), .CK(HCLK), .Q(vis_r0_o[26]), .QN(n6306) );
  DFF_X1 Zazpw6_reg ( .D(P5shu6), .CK(HCLK), .Q(vis_psp_o[24]), .QN(n4066) );
  DFF_X1 Xztpw6_reg ( .D(L3shu6), .CK(HCLK), .Q(vis_r11_o[26]), .QN(n8123) );
  DFF_X1 Xxtpw6_reg ( .D(X2shu6), .CK(HCLK), .Q(vis_r9_o[26]), .QN(n6080) );
  DFF_X1 Xxlax6_reg ( .D(E3shu6), .CK(HCLK), .Q(vis_r10_o[26]), .QN(n8071) );
  DFF_X1 Xvtpw6_reg ( .D(C2shu6), .CK(HCLK), .Q(vis_r1_o[26]), .QN(n4070) );
  DFF_X1 X3upw6_reg ( .D(D6shu6), .CK(HCLK), .Q(vis_r8_o[26]), .QN(n5895) );
  DFF_X1 X1upw6_reg ( .D(Z3shu6), .CK(HCLK), .Q(vis_r5_o[26]), .QN(n6395) );
  DFF_X1 Wluax6_reg ( .D(S3shu6), .CK(HCLK), .Q(vis_r4_o[26]), .QN(n5369) );
  DFF_X1 Vgqax6_reg ( .D(J2shu6), .CK(HCLK), .Q(vis_r2_o[26]), .QN(n5556) );
  DFF_X1 Tyzpw6_reg ( .D(I5shu6), .CK(HCLK), .Q(vis_msp_o[24]), .QN(n5961) );
  DFF_X1 Nk5bx6_reg ( .D(Q2shu6), .CK(HCLK), .Q(vis_r3_o[26]), .QN(n7377) );
  DFF_X1 Nhnax6_reg ( .D(B5shu6), .CK(HCLK), .Q(vis_r14_o[26]), .QN(n8282) );
  DFF_X1 M5wax6_reg ( .D(N4shu6), .CK(HCLK), .Q(vis_r7_o[26]), .QN(n7784) );
  DFF_X1 Fxoax6_reg ( .D(G4shu6), .CK(HCLK), .Q(vis_r6_o[26]), .QN(n5794) );
  DFF_X1 F4tax6_reg ( .D(U4shu6), .CK(HCLK), .Q(vis_r12_o[26]), .QN(n6202) );
  DFF_X1 E1npw6_reg ( .D(Gxrhu6), .CK(HCLK), .Q(vis_r0_o[27]), .QN(n6355) );
  DFF_X1 Zczpw6_reg ( .D(A1shu6), .CK(HCLK), .Q(vis_psp_o[25]), .QN(n3604) );
  DFF_X1 Xzlax6_reg ( .D(Pyrhu6), .CK(HCLK), .Q(vis_r10_o[27]), .QN(n8058) );
  DFF_X1 Wnuax6_reg ( .D(Dzrhu6), .CK(HCLK), .Q(vis_r4_o[27]), .QN(n5451) );
  DFF_X1 Viqax6_reg ( .D(Uxrhu6), .CK(HCLK), .Q(vis_r2_o[27]), .QN(n5493) );
  DFF_X1 T00qw6_reg ( .D(T0shu6), .CK(HCLK), .Q(vis_msp_o[25]), .QN(n5937) );
  DFF_X1 Otopw6_reg ( .D(Iyrhu6), .CK(HCLK), .Q(vis_r9_o[27]), .QN(n6148) );
  DFF_X1 Nm5bx6_reg ( .D(Byrhu6), .CK(HCLK), .Q(vis_r3_o[27]), .QN(n3607) );
  DFF_X1 Njnax6_reg ( .D(M0shu6), .CK(HCLK), .Q(vis_r14_o[27]), .QN(n8092) );
  DFF_X1 Mlmpw6_reg ( .D(O1shu6), .CK(HCLK), .Q(vis_r8_o[27]), .QN(n5873) );
  DFF_X1 Mjmpw6_reg ( .D(Wyrhu6), .CK(HCLK), .Q(vis_r11_o[27]), .QN(n8107) );
  DFF_X1 M7wax6_reg ( .D(Yzrhu6), .CK(HCLK), .Q(vis_r7_o[27]), .QN(n7704) );
  DFF_X1 Lfppw6_reg ( .D(Kzrhu6), .CK(HCLK), .Q(vis_r5_o[27]), .QN(n6560) );
  DFF_X1 Ixppw6_reg ( .D(Nxrhu6), .CK(HCLK), .Q(vis_r1_o[27]), .QN(n6650) );
  DFF_X1 Fzoax6_reg ( .D(Rzrhu6), .CK(HCLK), .Q(vis_r6_o[27]), .QN(n5689) );
  DFF_X1 F6tax6_reg ( .D(F0shu6), .CK(HCLK), .Q(vis_r12_o[27]), .QN(n6266) );
  DFF_X1 Ednpw6_reg ( .D(Rgphu6), .CK(HCLK), .Q(vis_r0_o[28]), .QN(n8267) );
  DFF_X1 Uqipw6_reg ( .D(Oiphu6), .CK(HCLK), .Q(vis_r11_o[28]), .QN(n8269) );
  DFF_X1 Rtibx6_reg ( .D(Skphu6), .CK(HCLK), .Q(vis_psp_o[26]), .QN(n8266) );
  DFF_X1 Rribx6_reg ( .D(Ekphu6), .CK(HCLK), .Q(vis_r14_o[28]), .QN(n8275) );
  DFF_X1 Rpibx6_reg ( .D(Xjphu6), .CK(HCLK), .Q(vis_r12_o[28]), .QN(n8263) );
  DFF_X1 Rnibx6_reg ( .D(Qjphu6), .CK(HCLK), .Q(vis_r7_o[28]), .QN(n8268) );
  DFF_X1 Rlibx6_reg ( .D(Jjphu6), .CK(HCLK), .Q(vis_r6_o[28]), .QN(n8272) );
  DFF_X1 Rjibx6_reg ( .D(Cjphu6), .CK(HCLK), .Q(vis_r5_o[28]), .QN(n8276) );
  DFF_X1 Rhibx6_reg ( .D(Viphu6), .CK(HCLK), .Q(vis_r4_o[28]), .QN(n8264) );
  DFF_X1 Rfibx6_reg ( .D(Hiphu6), .CK(HCLK), .Q(vis_r10_o[28]), .QN(n8273) );
  DFF_X1 Rdibx6_reg ( .D(Aiphu6), .CK(HCLK), .Q(vis_r9_o[28]), .QN(n8277) );
  DFF_X1 Rbibx6_reg ( .D(Thphu6), .CK(HCLK), .Q(vis_r8_o[28]), .QN(n8265) );
  DFF_X1 R9ibx6_reg ( .D(Mhphu6), .CK(HCLK), .Q(vis_r3_o[28]), .QN(n8270) );
  DFF_X1 R7ibx6_reg ( .D(Fhphu6), .CK(HCLK), .Q(vis_r2_o[28]), .QN(n8274) );
  DFF_X1 Pejbx6_reg ( .D(Lkphu6), .CK(HCLK), .Q(vis_msp_o[26]), .QN(n8271) );
  DFF_X1 I9qpw6_reg ( .D(Ygphu6), .CK(HCLK), .Q(vis_r1_o[28]), .QN(n8262) );
  DFF_X1 E3npw6_reg ( .D(Ysrhu6), .CK(HCLK), .Q(vis_r0_o[29]), .QN(n6289) );
  DFF_X1 Zezpw6_reg ( .D(Swrhu6), .CK(HCLK), .Q(vis_psp_o[27]), .QN(n3587) );
  DFF_X1 X1max6_reg ( .D(Hurhu6), .CK(HCLK), .Q(vis_r10_o[29]), .QN(n8067) );
  DFF_X1 Wpuax6_reg ( .D(Vurhu6), .CK(HCLK), .Q(vis_r4_o[29]), .QN(n5333) );
  DFF_X1 Vkqax6_reg ( .D(Mtrhu6), .CK(HCLK), .Q(vis_r2_o[29]), .QN(n5540) );
  DFF_X1 T20qw6_reg ( .D(Lwrhu6), .CK(HCLK), .Q(vis_msp_o[27]), .QN(n5955) );
  DFF_X1 Ovopw6_reg ( .D(Aurhu6), .CK(HCLK), .Q(vis_r9_o[29]), .QN(n3031) );
  DFF_X1 No5bx6_reg ( .D(Ttrhu6), .CK(HCLK), .Q(vis_r3_o[29]), .QN(n7341) );
  DFF_X1 Nlnax6_reg ( .D(Ewrhu6), .CK(HCLK), .Q(vis_r14_o[29]), .QN(n8098) );
  DFF_X1 M9wax6_reg ( .D(Qvrhu6), .CK(HCLK), .Q(vis_r7_o[29]), .QN(n7775) );
  DFF_X1 Lhppw6_reg ( .D(Cvrhu6), .CK(HCLK), .Q(vis_r5_o[29]), .QN(n6590) );
  DFF_X1 Kmjpw6_reg ( .D(Zwrhu6), .CK(HCLK), .Q(vis_r8_o[29]), .QN(n5811) );
  DFF_X1 Kkjpw6_reg ( .D(Ourhu6), .CK(HCLK), .Q(vis_r11_o[29]), .QN(n8120) );
  DFF_X1 Izppw6_reg ( .D(Ftrhu6), .CK(HCLK), .Q(vis_r1_o[29]), .QN(n6819) );
  DFF_X1 F8tax6_reg ( .D(Xvrhu6), .CK(HCLK), .Q(vis_r12_o[29]), .QN(n6178) );
  DFF_X1 F1pax6_reg ( .D(Jvrhu6), .CK(HCLK), .Q(vis_r6_o[29]), .QN(n5739) );
  DFF_X1 Gvmpw6_reg ( .D(Ocvhu6), .CK(HCLK), .Q(vis_r0_o[30]), .QN(n6324) );
  DFF_X1 Ykzpw6_reg ( .D(S2thu6), .CK(HCLK), .Q(vis_msp_o[28]), .QN(n5939) );
  DFF_X1 Weipw6_reg ( .D(Vcvhu6), .CK(HCLK), .Q(vis_r1_o[30]), .QN(n6605) );
  DFF_X1 Vxxax6_reg ( .D(Wbthu6), .CK(HCLK), .Q(vis_r3_o[30]), .QN(n6918) );
  DFF_X1 Uoipw6_reg ( .D(Wxshu6), .CK(HCLK), .Q(vis_r11_o[30]), .QN(n8108) );
  DFF_X1 S1nax6_reg ( .D(C1thu6), .CK(HCLK), .Q(vis_r14_o[30]), .QN(n8100) );
  DFF_X1 Rpvax6_reg ( .D(K5thu6), .CK(HCLK), .Q(vis_r7_o[30]), .QN(n7793) );
  DFF_X1 Qlopw6_reg ( .D(Qushu6), .CK(HCLK), .Q(vis_r9_o[30]), .QN(n6120) );
  DFF_X1 Qkrax6_reg ( .D(Rsrhu6), .CK(HCLK), .Q(vis_r8_o[30]), .QN(n5849) );
  DFF_X1 N7ppw6_reg ( .D(Q8thu6), .CK(HCLK), .Q(vis_r5_o[30]), .QN(n6486) );
  DFF_X1 Kosax6_reg ( .D(Mzshu6), .CK(HCLK), .Q(vis_r12_o[30]), .QN(n6221) );
  DFF_X1 Khoax6_reg ( .D(A7thu6), .CK(HCLK), .Q(vis_r6_o[30]), .QN(n2758) );
  DFF_X1 Exypw6_reg ( .D(B4thu6), .CK(HCLK), .Q(vis_psp_o[28]), .QN(n3601) );
  DFF_X1 Cilax6_reg ( .D(Gwshu6), .CK(HCLK), .Q(vis_r10_o[30]), .QN(n8069) );
  DFF_X1 B6uax6_reg ( .D(Gathu6), .CK(HCLK), .Q(vis_r4_o[30]), .QN(n5433) );
  DFF_X1 A1qax6_reg ( .D(Mdthu6), .CK(HCLK), .Q(vis_r2_o[30]), .QN(n5541) );
  DFF_X1 Yizpw6_reg ( .D(Z2thu6), .CK(HCLK), .Q(vis_msp_o[29]), .QN(n5898) );
  DFF_X1 Vzxax6_reg ( .D(Pbthu6), .CK(HCLK), .Q(vis_r3_o[31]), .QN(n7512) );
  DFF_X1 S3nax6_reg ( .D(V0thu6), .CK(HCLK), .Q(vis_r14_o[31]), .QN(n8077) );
  DFF_X1 Rrvax6_reg ( .D(D5thu6), .CK(HCLK), .Q(vis_r7_o[31]), .QN(n7811) );
  DFF_X1 Qnopw6_reg ( .D(Jushu6), .CK(HCLK), .Q(vis_r9_o[31]), .QN(n6146) );
  DFF_X1 Qmrax6_reg ( .D(Wrrhu6), .CK(HCLK), .Q(vis_r8_o[31]), .QN(n5829) );
  DFF_X1 N9ppw6_reg ( .D(J8thu6), .CK(HCLK), .Q(vis_r5_o[31]), .QN(n6577) );
  DFF_X1 Kqsax6_reg ( .D(Fzshu6), .CK(HCLK), .Q(vis_r12_o[31]), .QN(n6253) );
  DFF_X1 Kjoax6_reg ( .D(T6thu6), .CK(HCLK), .Q(vis_r6_o[31]), .QN(n5684) );
  DFF_X1 Evypw6_reg ( .D(I4thu6), .CK(HCLK), .Q(vis_psp_o[29]), .QN(n3593) );
  DFF_X1 Ejnpw6_reg ( .D(Jdvhu6), .CK(HCLK), .Q(vis_r1_o[31]), .QN(n6677) );
  DFF_X1 Ehnpw6_reg ( .D(Cdvhu6), .CK(HCLK), .Q(vis_r0_o[31]), .QN(n2815) );
  DFF_X1 Efnpw6_reg ( .D(Pxshu6), .CK(HCLK), .Q(vis_r11_o[31]), .QN(n8118) );
  DFF_X1 Cklax6_reg ( .D(Zvshu6), .CK(HCLK), .Q(vis_r10_o[31]), .QN(n7824) );
  DFF_X1 B8uax6_reg ( .D(Z9thu6), .CK(HCLK), .Q(vis_r4_o[31]), .QN(n5319) );
  DFF_X1 A3qax6_reg ( .D(Fdthu6), .CK(HCLK), .Q(vis_r2_o[31]), .QN(n5580) );
  DFFS_X1 Eliax6_reg ( .D(n7848), .CK(HCLK), .SN(HRESETn), .Q(vis_ipsr_o[0]), 
        .QN(n5112) );
  DFFS_X1 Pcrpw6_reg ( .D(n7846), .CK(HCLK), .SN(HRESETn), .Q(vis_ipsr_o[1]), 
        .QN(n3968) );
  DFFS_X1 Lerpw6_reg ( .D(n7827), .CK(HCLK), .SN(HRESETn), .Q(vis_pc_o[0]), 
        .QN(n4548) );
  DFFS_X1 Zshax6_reg ( .D(n7813), .CK(HCLK), .SN(HRESETn), .Q(vis_pc_o[4]), 
        .QN(n4782) );
  DFFS_X1 Cq7bx6_reg ( .D(n7785), .CK(HCLK), .SN(HRESETn), .Q(vis_pc_o[14]), 
        .QN(n4776) );
  DFFS_X1 Zdhax6_reg ( .D(n7776), .CK(HCLK), .SN(HRESETn), .Q(vis_pc_o[17]), 
        .QN(n8174) );
  DFFS_X1 Wfhax6_reg ( .D(n7779), .CK(HCLK), .SN(HRESETn), .Q(vis_pc_o[16]), 
        .QN(n4773) );
  DFFS_X1 Thhax6_reg ( .D(n7782), .CK(HCLK), .SN(HRESETn), .Q(vis_pc_o[15]), 
        .QN(n4774) );
  DFFS_X1 Nxabx6_reg ( .D(n7764), .CK(HCLK), .SN(HRESETn), .Q(vis_pc_o[21]), 
        .QN(n4766) );
  DFFS_X1 I8hax6_reg ( .D(n7767), .CK(HCLK), .SN(HRESETn), .Q(vis_pc_o[20]), 
        .QN(n4772) );
  DFFS_X1 Fahax6_reg ( .D(n7770), .CK(HCLK), .SN(HRESETn), .Q(vis_pc_o[19]), 
        .QN(n4184) );
  DFFS_X1 Cchax6_reg ( .D(n7773), .CK(HCLK), .SN(HRESETn), .Q(vis_pc_o[18]), 
        .QN(n8193) );
  DFFS_X1 C37ax6_reg ( .D(n7761), .CK(HCLK), .SN(HRESETn), .Q(vis_pc_o[22]), 
        .QN(n4765) );
  DFFS_X1 Drhax6_reg ( .D(n7812), .CK(HCLK), .SN(HRESETn), .Q(vis_pc_o[5]), 
        .QN(n4816) );
  DFFS_X1 Rwhax6_reg ( .D(n7819), .CK(HCLK), .SN(HRESETn), .Q(vis_pc_o[2]), 
        .QN(n4787) );
  DFFS_X1 P7bbx6_reg ( .D(n7798), .CK(HCLK), .SN(HRESETn), .Q(vis_pc_o[9]), 
        .QN(n4807) );
  DFFS_X1 Hphax6_reg ( .D(n7804), .CK(HCLK), .SN(HRESETn), .Q(vis_pc_o[7]), 
        .QN(n4810) );
  DFFS_X1 Knhax6_reg ( .D(n7794), .CK(HCLK), .SN(HRESETn), .Q(vis_pc_o[11]), 
        .QN(n4805) );
  DFFS_X1 Mw5bx6_reg ( .D(n7795), .CK(HCLK), .SN(HRESETn), .Q(vis_pc_o[10]), 
        .QN(n4806) );
  DFFS_X1 Equpw6_reg ( .D(n7807), .CK(HCLK), .SN(HRESETn), .Q(vis_pc_o[6]), 
        .QN(n4811) );
  DFFS_X1 Qjhax6_reg ( .D(n7788), .CK(HCLK), .SN(HRESETn), .Q(vis_pc_o[13]), 
        .QN(n4801) );
  DFFS_X1 Nlhax6_reg ( .D(n7791), .CK(HCLK), .SN(HRESETn), .Q(vis_pc_o[12]), 
        .QN(n4802) );
  DFFS_X1 J06bx6_reg ( .D(n7803), .CK(HCLK), .SN(HRESETn), .Q(vis_pc_o[8]), 
        .QN(n4777) );
  DFFS_X1 Nyhax6_reg ( .D(n7822), .CK(HCLK), .SN(HRESETn), .Q(vis_pc_o[1]), 
        .QN(n4795) );
  DFFS_X1 Vuhax6_reg ( .D(n7816), .CK(HCLK), .SN(HRESETn), .Q(vis_pc_o[3]), 
        .QN(n4783) );
  DFFS_X1 L6hax6_reg ( .D(n7758), .CK(HCLK), .SN(HRESETn), .Q(vis_pc_o[23]), 
        .QN(n4764) );
  DFFS_X1 O4hax6_reg ( .D(n7755), .CK(HCLK), .SN(HRESETn), .Q(vis_pc_o[24]), 
        .QN(n4799) );
  DFFS_X1 Pzkpw6_reg ( .D(Nfvhu6), .CK(HCLK), .SN(HRESETn), .Q(vis_tbit_o), 
        .QN(n3486) );
  DFFS_X1 R2hax6_reg ( .D(n7752), .CK(HCLK), .SN(HRESETn), .Q(vis_pc_o[25]), 
        .QN(n4797) );
  DFFS_X1 U0hax6_reg ( .D(n7749), .CK(HCLK), .SN(HRESETn), .Q(vis_pc_o[26]), 
        .QN(n3871) );
  DFFS_X1 D12qw6_reg ( .D(n7746), .CK(HCLK), .SN(HRESETn), .Q(vis_pc_o[27]), 
        .QN(n4110) );
  DFFS_X1 Lqjpw6_reg ( .D(n7743), .CK(HCLK), .SN(HRESETn), .Q(vis_pc_o[28]), 
        .QN(n4761) );
  DFFS_X1 A32qw6_reg ( .D(n7741), .CK(HCLK), .SN(HRESETn), .Q(vis_pc_o[29]), 
        .QN(n3124) );
  DFFS_X1 Awupw6_reg ( .D(n7739), .CK(HCLK), .SN(HRESETn), .Q(vis_pc_o[30]), 
        .QN(n3875) );
  DFFS_X1 Arnpw6_reg ( .D(Kgphu6), .CK(HCLK), .SN(HRESETn), .Q(vis_apsr_o[3]), 
        .QN(n2812) );
  DFFS_X1 Bfjpw6_reg ( .D(Ksrhu6), .CK(HCLK), .SN(HRESETn), .Q(vis_apsr_o[2]), 
        .QN(n2778) );
  DFFR_X1 Zszax6_reg ( .D(n7015), .CK(HCLK), .RN(HRESETn), .Q(n8154), .QN(
        n6760) );
  DFFR_X1 Kqhbx6_reg ( .D(n7029), .CK(HCLK), .RN(HRESETn), .Q(n4535), .QN(
        n7688) );
  DFFR_X1 Lp7ax6_reg ( .D(n7723), .CK(HCLK), .RN(HRESETn), .QN(n7442) );
  DFFR_X1 I2zax6_reg ( .D(n7721), .CK(HCLK), .RN(HRESETn), .Q(n8133), .QN(
        n7560) );
  DFFR_X1 G0zax6_reg ( .D(n7718), .CK(HCLK), .RN(HRESETn), .Q(n4491), .QN(
        n7559) );
  DFFR_X1 Avzax6_reg ( .D(n7720), .CK(HCLK), .RN(HRESETn), .Q(n8155), .QN(
        n7570) );
  DFFR_X1 Owhbx6_reg ( .D(n7960), .CK(HCLK), .RN(HRESETn), .Q(n8144), .QN(
        n7690) );
  DFFR_X1 C3wpw6_reg ( .D(n7947), .CK(HCLK), .RN(HRESETn), .Q(n8136), .QN(
        n7384) );
  DFFR_X1 Ikhbx6_reg ( .D(n7964), .CK(HCLK), .RN(HRESETn), .Q(n8146), .QN(
        n7685) );
  DFFR_X1 Czzax6_reg ( .D(n7968), .CK(HCLK), .RN(HRESETn), .Q(n8281), .QN(
        n7572) );
  DFFR_X1 L1bbx6_reg ( .D(n7955), .CK(HCLK), .RN(HRESETn), .Q(n8142) );
  DFFR_X1 Z9abx6_reg ( .D(n7057), .CK(HCLK), .RN(HRESETn), .QN(n7638) );
  DFFR_X1 X7abx6_reg ( .D(n7050), .CK(HCLK), .RN(HRESETn), .QN(n7637) );
  DFFR_X1 V5abx6_reg ( .D(n7037), .CK(HCLK), .RN(HRESETn), .QN(n6773) );
  DFFR_X1 T3abx6_reg ( .D(n7011), .CK(HCLK), .RN(HRESETn), .QN(n7636) );
  DFFR_X1 R1abx6_reg ( .D(n7053), .CK(HCLK), .RN(HRESETn), .QN(n6778) );
  DFFR_X1 Pz9bx6_reg ( .D(n7043), .CK(HCLK), .RN(HRESETn), .QN(n6775) );
  DFFR_X1 Nv9bx6_reg ( .D(n7033), .CK(HCLK), .RN(HRESETn), .QN(n7634) );
  DFFR_X1 Bcabx6_reg ( .D(n7007), .CK(HCLK), .RN(HRESETn), .QN(n7639) );
  DFFR_X1 Yqzax6_reg ( .D(n6946), .CK(HCLK), .RN(HRESETn), .Q(n8236), .QN(
        n7569) );
  DFFR_X1 Wu3bx6_reg ( .D(n6949), .CK(HCLK), .RN(HRESETn), .Q(n8233), .QN(
        n6711) );
  DFFR_X1 Sn4bx6_reg ( .D(n6948), .CK(HCLK), .RN(HRESETn), .Q(n8234), .QN(
        n6710) );
  DFFR_X1 S3mpw6_reg ( .D(n6954), .CK(HCLK), .RN(HRESETn), .Q(n8228), .QN(
        n7323) );
  DFFR_X1 Mfyax6_reg ( .D(n6950), .CK(HCLK), .RN(HRESETn), .Q(n8232), .QN(
        n7551) );
  DFFR_X1 I74bx6_reg ( .D(n6953), .CK(HCLK), .RN(HRESETn), .Q(n8229), .QN(
        n7610) );
  DFFR_X1 H4zax6_reg ( .D(n6951), .CK(HCLK), .RN(HRESETn), .Q(n8231), .QN(
        n6712) );
  DFFR_X1 E05bx6_reg ( .D(n6952), .CK(HCLK), .RN(HRESETn), .Q(n8230), .QN(
        n7621) );
  DFFR_X1 Cxzax6_reg ( .D(n7851), .CK(HCLK), .RN(HRESETn), .Q(n8134) );
  DFFR_X1 Nt9bx6_reg ( .D(n7971), .CK(HCLK), .RN(HRESETn), .Q(n8149), .QN(
        n7633) );
  DFFR_X1 C10bx6_reg ( .D(n7975), .CK(HCLK), .RN(HRESETn), .Q(n8237) );
  DFFR_X1 Ih0bx6_reg ( .D(n7950), .CK(HCLK), .RN(HRESETn), .Q(n8139), .QN(
        n6634) );
  DFFR_X1 Kl0bx6_reg ( .D(n7954), .CK(HCLK), .RN(HRESETn), .Q(n8141), .QN(
        n6631) );
  DFFR_X1 Kojpw6_reg ( .D(n7966), .CK(HCLK), .RN(HRESETn), .Q(n8147), .QN(
        n7280) );
  DFFR_X1 Oxkpw6_reg ( .D(n7948), .CK(HCLK), .RN(HRESETn), .Q(n8137) );
  DFFR_X1 Pv0bx6_reg ( .D(n7977), .CK(HCLK), .RN(HRESETn), .Q(n8152), .QN(
        n7581) );
  DFFR_X1 Jj0bx6_reg ( .D(n7976), .CK(HCLK), .RN(HRESETn), .Q(n8151), .QN(
        n7576) );
  DFFR_X1 Ln0bx6_reg ( .D(n7959), .CK(HCLK), .RN(HRESETn), .Q(n8143) );
  DFFR_X1 Mp0bx6_reg ( .D(n7963), .CK(HCLK), .RN(HRESETn), .Q(n8225) );
  DFFR_X1 Nr0bx6_reg ( .D(n7967), .CK(HCLK), .RN(HRESETn), .Q(n8148) );
  DFFR_X1 Usipw6_reg ( .D(n7962), .CK(HCLK), .RN(HRESETn), .Q(n8278) );
  DFFR_X1 Fb0bx6_reg ( .D(n7965), .CK(HCLK), .RN(HRESETn), .QN(n7574) );
  DFFR_X1 E90bx6_reg ( .D(n7961), .CK(HCLK), .RN(HRESETn), .Q(n8145), .QN(
        n6629) );
  DFFR_X1 D70bx6_reg ( .D(n7956), .CK(HCLK), .RN(HRESETn), .Q(n8165), .QN(
        n6630) );
  DFFR_X1 C50bx6_reg ( .D(n7951), .CK(HCLK), .RN(HRESETn), .Q(n8169), .QN(
        n6633) );
  DFFR_X1 Tngbx6_reg ( .D(n6977), .CK(HCLK), .RN(HRESETn), .QN(n7678) );
  DFFR_X1 Rlgbx6_reg ( .D(n6978), .CK(HCLK), .RN(HRESETn), .QN(n7677) );
  DFFR_X1 Pjgbx6_reg ( .D(n6979), .CK(HCLK), .RN(HRESETn), .Q(n8199), .QN(
        n6735) );
  DFFR_X1 Nhgbx6_reg ( .D(n6980), .CK(HCLK), .RN(HRESETn), .QN(n7676) );
  DFFR_X1 Lfgbx6_reg ( .D(n6981), .CK(HCLK), .RN(HRESETn), .Q(n8198), .QN(
        n7675) );
  DFFR_X1 Jdgbx6_reg ( .D(n6982), .CK(HCLK), .RN(HRESETn), .QN(n7674) );
  DFFR_X1 Hbgbx6_reg ( .D(n6983), .CK(HCLK), .RN(HRESETn), .QN(n7673) );
  DFFR_X1 C5gbx6_reg ( .D(n6985), .CK(HCLK), .RN(HRESETn), .QN(n7670) );
  DFFR_X1 Yt4bx6_reg ( .D(n7046), .CK(HCLK), .RN(HRESETn), .Q(n4468), .QN(
        n7619) );
  DFFR_X1 Vkzax6_reg ( .D(n7034), .CK(HCLK), .RN(HRESETn), .Q(n4487), .QN(
        n7566) );
  DFFR_X1 Slyax6_reg ( .D(n7014), .CK(HCLK), .RN(HRESETn), .Q(n8157), .QN(
        n7554) );
  DFFR_X1 Od4bx6_reg ( .D(n7060), .CK(HCLK), .RN(HRESETn), .Q(n4433), .QN(
        n7612) );
  DFFR_X1 Nazax6_reg ( .D(n7040), .CK(HCLK), .RN(HRESETn), .Q(n4474), .QN(
        n7563) );
  DFFR_X1 K65bx6_reg ( .D(n7047), .CK(HCLK), .RN(HRESETn), .Q(n4467), .QN(
        n6777) );
  DFFR_X1 C14bx6_reg ( .D(n7056), .CK(HCLK), .RN(HRESETn), .QN(n7607) );
  DFFR_X1 Auyax6_reg ( .D(n7010), .CK(HCLK), .RN(HRESETn), .Q(n8159), .QN(
        n7557) );
  DFFR_X1 Vpgbx6_reg ( .D(n6976), .CK(HCLK), .RN(HRESETn), .Q(n8200), .QN(
        n7679) );
  DFFR_X1 Gz6ax6_reg ( .D(n7211), .CK(HCLK), .RN(HRESETn), .Q(n3785), .QN(
        n7434) );
  DFFR_X1 B3gbx6_reg ( .D(n7970), .CK(HCLK), .RN(HRESETn), .Q(n8201) );
  DFFR_X1 Ot0bx6_reg ( .D(n7974), .CK(HCLK), .RN(HRESETn), .Q(n8292) );
  DFFR_X1 Tkjbx6_reg ( .D(n7978), .CK(HCLK), .RN(HRESETn), .Q(n8153), .QN(
        n7697) );
  DFFR_X1 C30bx6_reg ( .D(n7949), .CK(HCLK), .RN(HRESETn), .Q(n8138), .QN(
        n6635) );
  DFFR_X1 X5upw6_reg ( .D(n7953), .CK(HCLK), .RN(HRESETn), .Q(n8140), .QN(
        n6632) );
  DFFR_X1 Qx0bx6_reg ( .D(n7958), .CK(HCLK), .RN(HRESETn), .Q(n8295), .QN(
        n7582) );
  DFFR_X1 Yw3bx6_reg ( .D(n6936), .CK(HCLK), .RN(HRESETn), .Q(n8255), .QN(
        n7605) );
  DFFR_X1 Xozax6_reg ( .D(n6939), .CK(HCLK), .RN(HRESETn), .Q(n8254), .QN(
        n7568) );
  DFFR_X1 Vbspw6_reg ( .D(n6931), .CK(HCLK), .RN(HRESETn), .Q(n8256), .QN(
        n6700) );
  DFFR_X1 Up4bx6_reg ( .D(n6937), .CK(HCLK), .RN(HRESETn), .QN(n7617) );
  DFFR_X1 Ohyax6_reg ( .D(n6935), .CK(HCLK), .RN(HRESETn), .QN(n7552) );
  DFFR_X1 K94bx6_reg ( .D(n6932), .CK(HCLK), .RN(HRESETn), .QN(n6701) );
  DFFR_X1 J6zax6_reg ( .D(n6934), .CK(HCLK), .RN(HRESETn), .QN(n7561) );
  DFFR_X1 G25bx6_reg ( .D(n6933), .CK(HCLK), .RN(HRESETn), .QN(n6702) );
  DFFR_X1 Unyax6_reg ( .D(n7013), .CK(HCLK), .RN(HRESETn), .QN(n6759) );
  DFFR_X1 Uizax6_reg ( .D(n7035), .CK(HCLK), .RN(HRESETn), .QN(n6772) );
  DFFR_X1 Qf4bx6_reg ( .D(n7059), .CK(HCLK), .RN(HRESETn), .QN(n7613) );
  DFFR_X1 Pczax6_reg ( .D(n7039), .CK(HCLK), .RN(HRESETn), .QN(n6774) );
  DFFR_X1 M85bx6_reg ( .D(n7048), .CK(HCLK), .RN(HRESETn), .QN(n7623) );
  DFFR_X1 E34bx6_reg ( .D(n7055), .CK(HCLK), .RN(HRESETn), .Q(n4442), .QN(
        n7608) );
  DFFR_X1 Cwyax6_reg ( .D(n7009), .CK(HCLK), .RN(HRESETn), .Q(n8160), .QN(
        n6758) );
  DFFR_X1 Aw4bx6_reg ( .D(n7045), .CK(HCLK), .RN(HRESETn), .QN(n6776) );
  DFFR_X1 Wpyax6_reg ( .D(n7012), .CK(HCLK), .RN(HRESETn), .Q(n8158), .QN(
        n7555) );
  DFFR_X1 Tgzax6_reg ( .D(n7036), .CK(HCLK), .RN(HRESETn), .Q(n4482), .QN(
        n7565) );
  DFFR_X1 Sh4bx6_reg ( .D(n7058), .CK(HCLK), .RN(HRESETn), .Q(n4434), .QN(
        n7614) );
  DFFR_X1 Rezax6_reg ( .D(n7038), .CK(HCLK), .RN(HRESETn), .Q(n4478), .QN(
        n7564) );
  DFFR_X1 Oa5bx6_reg ( .D(n7049), .CK(HCLK), .RN(HRESETn), .Q(n4466), .QN(
        n7624) );
  DFFR_X1 G54bx6_reg ( .D(n7054), .CK(HCLK), .RN(HRESETn), .Q(n4453), .QN(
        n7609) );
  DFFR_X1 Eyyax6_reg ( .D(n7008), .CK(HCLK), .RN(HRESETn), .Q(n8161), .QN(
        n7558) );
  DFFR_X1 Cy4bx6_reg ( .D(n7044), .CK(HCLK), .RN(HRESETn), .Q(n4470), .QN(
        n7620) );
  DFFR_X1 Wgipw6_reg ( .D(n7042), .CK(HCLK), .RN(HRESETn), .QN(n7257) );
  DFFR_X1 Tl4bx6_reg ( .D(n7051), .CK(HCLK), .RN(HRESETn), .Q(n4459), .QN(
        n7616) );
  DFFR_X1 Gd0bx6_reg ( .D(n7969), .CK(HCLK), .RN(HRESETn), .Q(n8257), .QN(
        n6627) );
  DFFR_X1 Yryax6_reg ( .D(n7709), .CK(HCLK), .RN(HRESETn), .Q(n8241), .QN(
        n7556) );
  DFFR_X1 Wr4bx6_reg ( .D(n7715), .CK(HCLK), .RN(HRESETn), .Q(n8247), .QN(
        n7618) );
  DFFR_X1 Wmzax6_reg ( .D(n7717), .CK(HCLK), .RN(HRESETn), .Q(n8248), .QN(
        n7567) );
  DFFR_X1 Qjyax6_reg ( .D(n7710), .CK(HCLK), .RN(HRESETn), .Q(n8242), .QN(
        n7553) );
  DFFR_X1 Mb4bx6_reg ( .D(n7711), .CK(HCLK), .RN(HRESETn), .Q(n8243), .QN(
        n7611) );
  DFFR_X1 L8zax6_reg ( .D(n7713), .CK(HCLK), .RN(HRESETn), .Q(n8245), .QN(
        n7562) );
  DFFR_X1 I45bx6_reg ( .D(n7712), .CK(HCLK), .RN(HRESETn), .Q(n8244), .QN(
        n7622) );
  DFFR_X1 Az3bx6_reg ( .D(n7714), .CK(HCLK), .RN(HRESETn), .Q(n8246), .QN(
        n7606) );
  DFFR_X1 Uj4bx6_reg ( .D(n7052), .CK(HCLK), .RN(HRESETn), .Q(n4454), .QN(
        n7615) );
  DFFR_X1 Elnpw6_reg ( .D(n7041), .CK(HCLK), .RN(HRESETn), .Q(n4473), .QN(
        n7331) );
  DFFR_X1 Rz0bx6_reg ( .D(n7881), .CK(HCLK), .RN(HRESETn), .Q(n8135), .QN(
        n6660) );
  DFFR_X1 S0kbx6_reg ( .D(n7973), .CK(HCLK), .RN(HRESETn), .Q(n8150), .QN(
        n7701) );
  DFFR_X1 Hf0bx6_reg ( .D(n7972), .CK(HCLK), .RN(HRESETn), .Q(n8240) );
  DFFR_X1 F17ax6_reg ( .D(n7943), .CK(HCLK), .RN(HRESETn), .Q(n8291), .QN(
        n7435) );
  DFFR_X1 T8kbx6_reg ( .D(n7850), .CK(HCLK), .RN(HRESETn), .Q(n4673), .QN(
        n7705) );
  DFFR_X1 I8lax6_reg ( .D(n7032), .CK(HCLK), .RN(HRESETn), .QN(n7533) );
  DFFR_X1 U8jax6_reg ( .D(n7026), .CK(HCLK), .RN(HRESETn), .QN(n7507) );
  DFFR_X1 R3vpw6_reg ( .D(n7941), .CK(HCLK), .RN(HRESETn), .Q(n486), .QN(n7375) );
  DFFR_X1 Aujpw6_reg ( .D(n7942), .CK(HCLK), .RN(HRESETn), .Q(n265), .QN(n7282) );
  DFFR_X1 Vygax6_reg ( .D(n7825), .CK(HCLK), .RN(HRESETn), .Q(n4512), .QN(
        n7492) );
  DFFR_X1 S4kbx6_reg ( .D(Levhu6), .CK(HCLK), .RN(HRESETn), .Q(n4694), .QN(
        n7703) );
  DFFR_X1 Ms5bx6_reg ( .D(Lirhu6), .CK(HCLK), .RN(HRESETn), .Q(n8175), .QN(
        n7626) );
  DFFR_X1 Xxupw6_reg ( .D(Qrohu6), .CK(HCLK), .RN(HRESETn), .Q(n508), .QN(n267) );
  DFFR_X1 Zdiax6_reg ( .D(n7024), .CK(HCLK), .RN(HRESETn), .Q(n4753), .QN(
        n6768) );
  DFFR_X1 Hirpw6_reg ( .D(n7944), .CK(HCLK), .RN(HRESETn), .Q(n254), .QN(n7355) );
  DFFR_X1 Daiax6_reg ( .D(n8017), .CK(HCLK), .RN(HRESETn), .Q(n4826), .QN(
        n7497) );
  DFFR_X1 Ufopw6_reg ( .D(n7946), .CK(HCLK), .RN(HRESETn), .Q(n523), .QN(n228)
         );
  DFFR_X1 F9vpw6_reg ( .D(n7023), .CK(HCLK), .RN(HRESETn), .Q(n5225), .QN(
        n7378) );
  DFFR_X1 T1vpw6_reg ( .D(Crohu6), .CK(HCLK), .RN(HRESETn), .Q(n272), .QN(
        n7374) );
  DFFR_X1 Vzupw6_reg ( .D(Jrohu6), .CK(HCLK), .RN(HRESETn), .Q(n266), .QN(
        n7373) );
  DFFR_X1 Yvjpw6_reg ( .D(Twohu6), .CK(HCLK), .RN(HRESETn), .Q(n4263), .QN(
        n7283) );
  DFFR_X1 X7ypw6_reg ( .D(L0vhu6), .CK(HCLK), .RN(HRESETn), .Q(n2234), .QN(
        n6637) );
  DFFR_X1 C1wpw6_reg ( .D(Hyuhu6), .CK(HCLK), .RN(HRESETn), .Q(n3634), .QN(
        n7383) );
  DFFR_X1 Ztupw6_reg ( .D(n7732), .CK(HCLK), .RN(HRESETn), .Q(n4182), .QN(
        n7371) );
  DFFR_X1 W5ypw6_reg ( .D(n7731), .CK(HCLK), .RN(HRESETn), .Q(n4160), .QN(
        n7398) );
  DFFR_X1 R9yax6_reg ( .D(n7733), .CK(HCLK), .RN(HRESETn), .Q(n4410), .QN(
        n7548) );
  DFFR_X1 Yzspw6_reg ( .D(n7735), .CK(HCLK), .RN(HRESETn), .QN(n7363) );
  DFFR_X1 I5xax6_reg ( .D(n7734), .CK(HCLK), .RN(HRESETn), .Q(n4395), .QN(
        n7534) );
  DFFR_X1 Ydopw6_reg ( .D(n7726), .CK(HCLK), .RN(HRESETn), .Q(n529), .QN(n225)
         );
  DFF_X1 Oyhbx6_reg ( .D(n7031), .CK(HCLK), .QN(n7691) );
  DFF_X1 M6rpw6_reg ( .D(n7030), .CK(HCLK), .QN(n7351) );
  DFF_X1 Imhbx6_reg ( .D(n7028), .CK(HCLK), .Q(n4545), .QN(n7686) );
  DFF_X1 X5opw6_reg ( .D(n7210), .CK(HCLK), .QN(n7338) );
  DFF_X1 Vlxax6_reg ( .D(n7722), .CK(HCLK), .QN(n7542) );
  DFF_X1 Wnxax6_reg ( .D(n7719), .CK(HCLK), .QN(n7543) );
  DFF_X1 Ox9bx6_reg ( .D(n7197), .CK(HCLK), .QN(n7635) );
  DFF_X1 Thxax6_reg ( .D(n6947), .CK(HCLK), .Q(n8235), .QN(n7540) );
  DFF_X1 Tyipw6_reg ( .D(n7022), .CK(HCLK), .Q(n8104), .QN(n7275) );
  DFF_X1 Tptpw6_reg ( .D(n6999), .CK(HCLK), .QN(n7365) );
  DFF_X1 R7kpw6_reg ( .D(n7206), .CK(HCLK), .Q(n4161), .QN(n7287) );
  DFF_X1 Ofmpw6_reg ( .D(n7000), .CK(HCLK), .QN(n7327) );
  DFF_X1 Ujspw6_reg ( .D(n7204), .CK(HCLK), .QN(n7361) );
  DFF_X1 Lywpw6_reg ( .D(n7201), .CK(HCLK), .Q(n4163), .QN(n7390) );
  DFF_X1 Yjupw6_reg ( .D(n7203), .CK(HCLK), .QN(n7367) );
  DFF_X1 Hhvpw6_reg ( .D(n7202), .CK(HCLK), .QN(n7379) );
  DFF_X1 X6jpw6_reg ( .D(n6955), .CK(HCLK), .QN(n7277) );
  DFF_X1 Rhkpw6_reg ( .D(n7205), .CK(HCLK), .QN(n7289) );
  DFF_X1 D7gbx6_reg ( .D(n6984), .CK(HCLK), .Q(n8197), .QN(n7671) );
  DFF_X1 J7xax6_reg ( .D(n7199), .CK(HCLK), .QN(n7535) );
  DFF_X1 Tmjbx6_reg ( .D(n7198), .CK(HCLK), .QN(n7698) );
  DFF_X1 Rq0qw6_reg ( .D(n7200), .CK(HCLK), .QN(n7402) );
  DFF_X1 Pdxax6_reg ( .D(n6938), .CK(HCLK), .QN(n7538) );
  DFF_X1 L9xax6_reg ( .D(n7716), .CK(HCLK), .QN(n7536) );
  DFF_X1 Fpnpw6_reg ( .D(n8007), .CK(HCLK), .Q(n5257), .QN(n7332) );
  DFF_X1 Wxjpw6_reg ( .D(Mwohu6), .CK(HCLK), .Q(n5302), .QN(n7284) );
  DFF_X1 Shopw6_reg ( .D(Ntohu6), .CK(HCLK), .Q(n5304), .QN(n7343) );
  DFF_X1 M6kax6_reg ( .D(Gfohu6), .CK(HCLK), .Q(n5307), .QN(n7520) );
  DFF_X1 Dzvpw6_reg ( .D(Aqohu6), .CK(HCLK), .Q(n2466), .QN(n7382) );
  DFF_X1 Swjbx6_reg ( .D(n3520), .CK(HCLK), .Q(n8298) );
  DFF_X1 Jrypw6_reg ( .D(P9vhu6), .CK(HCLK), .Q(n4394), .QN(n7401) );
  DFF_X1 Vhspw6_reg ( .D(Lsohu6), .CK(HCLK), .Q(n5313), .QN(n7360) );
  DFF_X1 Iixpw6_reg ( .D(Q4xhu6), .CK(HCLK), .Q(n5312), .QN(n7394) );
  DFF_X1 Htmpw6_reg ( .D(Wuohu6), .CK(HCLK), .QN(n7330) );
  DFF_X1 Vmipw6_reg ( .D(Vxohu6), .CK(HCLK), .Q(n5291), .QN(n7274) );
  DFF_X1 V6jax6_reg ( .D(Miohu6), .CK(HCLK), .Q(n4637), .QN(n7506) );
  DFF_X1 Umkax6_reg ( .D(Leohu6), .CK(HCLK), .QN(n7527) );
  DFF_X1 Fkrpw6_reg ( .D(Ssohu6), .CK(HCLK), .Q(n5074), .QN(n7356) );
  DFF_X1 Ubypw6_reg ( .D(n7945), .CK(HCLK), .Q(n5070), .QN(n7400) );
  DFF_X1 Tokax6_reg ( .D(n8024), .CK(HCLK), .Q(n4703), .QN(n7528) );
  DFF_X1 Sujax6_reg ( .D(n8029), .CK(HCLK), .Q(n4720), .QN(n7515) );
  DFF_X1 Sqjax6_reg ( .D(n8030), .CK(HCLK), .Q(n4721), .QN(n7513) );
  DFF_X1 Smjax6_reg ( .D(n8031), .CK(HCLK), .Q(n4724), .QN(n7511) );
  DFF_X1 Sijax6_reg ( .D(n8032), .CK(HCLK), .Q(n5258), .QN(n7509) );
  DFF_X1 Sgjax6_reg ( .D(n8033), .CK(HCLK), .Q(n5266), .QN(n7508) );
  DFF_X1 Qyjax6_reg ( .D(n8028), .CK(HCLK), .Q(n4713), .QN(n7517) );
  DFF_X1 L8kax6_reg ( .D(n8026), .CK(HCLK), .Q(n4707), .QN(n7521) );
  DFF_X1 Kakax6_reg ( .D(n8025), .CK(HCLK), .Q(n4704), .QN(n7522) );
  DFF_X1 Rkkax6_reg ( .D(Cfthu6), .CK(HCLK), .Q(n4506), .QN(n6601) );
  DFF_X1 Iekax6_reg ( .D(Xfthu6), .CK(HCLK), .Q(n3571), .QN(n7524) );
  DFF_X1 Lgkax6_reg ( .D(n8005), .CK(HCLK), .Q(n5065), .QN(n7525) );
  DFF_X1 U1kpw6_reg ( .D(Vethu6), .CK(HCLK), .Q(n5299), .QN(n7286) );
  DFF_X1 Sqkax6_reg ( .D(Pgvhu6), .CK(HCLK), .Q(n5293), .QN(n7529) );
  DFF_X1 Rskax6_reg ( .D(Oethu6), .CK(HCLK), .Q(n3083), .QN(n7530) );
  DFF_X1 R9mpw6_reg ( .D(L7vhu6), .CK(HCLK), .Q(n5294), .QN(n7326) );
  DFF_X1 Oikax6_reg ( .D(n8006), .CK(HCLK), .Q(n3576), .QN(n7526) );
  DFF_X1 Xrxax6_reg ( .D(n7823), .CK(HCLK), .Q(n8168), .QN(n7545) );
  DFF_X1 N61qw6_reg ( .D(n7805), .CK(HCLK), .Q(n4009), .QN(n7404) );
  DFF_X1 Gwxpw6_reg ( .D(n7799), .CK(HCLK), .Q(n8171), .QN(n7395) );
  DFF_X1 Dm6bx6_reg ( .D(n7792), .CK(HCLK), .Q(n8103), .QN(n7629) );
  DFF_X1 C07bx6_reg ( .D(n7796), .CK(HCLK), .Q(n8163), .QN(n7630) );
  DFF_X1 Asupw6_reg ( .D(n7808), .CK(HCLK), .Q(n4940) );
  DFF_X1 Xpxax6_reg ( .D(n7789), .CK(HCLK), .Q(n3041), .QN(n7544) );
  DFF_X1 Qc5bx6_reg ( .D(n7814), .CK(HCLK), .Q(n8082), .QN(n7625) );
  DFF_X1 Wtxax6_reg ( .D(n7817), .CK(HCLK), .Q(n8167), .QN(n7546) );
  DFF_X1 T5yax6_reg ( .D(n7820), .CK(HCLK), .Q(n8111), .QN(n7547) );
  DFF_X1 Nu5bx6_reg ( .D(n7826), .CK(HCLK), .Q(n4348), .QN(n7627) );
  DFF_X1 Kn1qw6_reg ( .D(n7801), .CK(HCLK), .Q(n8173), .QN(n7408) );
  DFF_X1 Sb8ax6_reg ( .D(n7786), .CK(HCLK), .Q(n8252), .QN(n7446) );
  DFF_X1 Z47ax6_reg ( .D(n7783), .CK(HCLK), .Q(n8116), .QN(n7436) );
  DFF_X1 Chwpw6_reg ( .D(n7780), .CK(HCLK), .Q(n4185), .QN(n7385) );
  DFF_X1 Pbbbx6_reg ( .D(n7777), .CK(HCLK), .Q(n3280), .QN(n7647) );
  DFF_X1 Syjbx6_reg ( .D(n7774), .CK(HCLK), .Q(n8177), .QN(n7700) );
  DFF_X1 T6kbx6_reg ( .D(n7771), .CK(HCLK), .Q(n8224) );
  DFF_X1 Fjdbx6_reg ( .D(n7768), .CK(HCLK), .Q(n8223), .QN(n7660) );
  DFF_X1 M2ebx6_reg ( .D(n7765), .CK(HCLK), .Q(n3672), .QN(n7663) );
  DFF_X1 Tlebx6_reg ( .D(n7762), .CK(HCLK), .Q(n8196), .QN(n7666) );
  DFF_X1 Ztgbx6_reg ( .D(n7759), .CK(HCLK), .Q(n8195), .QN(n7680) );
  DFF_X1 Tgkbx6_reg ( .D(n7756), .CK(HCLK), .Q(n3484), .QN(n7706) );
  DFF_X1 F8cbx6_reg ( .D(n7750), .CK(HCLK), .Q(n8283), .QN(n7654) );
  DFF_X1 Nybbx6_reg ( .D(n7747), .CK(HCLK), .Q(n8297), .QN(n7649) );
  DFF_X1 Ibqpw6_reg ( .D(n7744), .CK(HCLK), .Q(n8261), .QN(n7344) );
  DFF_X1 Sx3qw6_reg ( .D(n7742), .CK(HCLK), .Q(n8204), .QN(n7432) );
  DFF_X1 F6dbx6_reg ( .D(n7740), .CK(HCLK), .Q(n2779), .QN(n7658) );
  DFF_X1 Usnpw6_reg ( .D(n7736), .CK(HCLK), .Q(n2814), .QN(n7333) );
  DFF_X1 Vgjpw6_reg ( .D(Oxohu6), .CK(HCLK), .Q(n2731), .QN(n7279) );
  DFF_X1 Z8jpw6_reg ( .D(n7983), .CK(SCLK), .Q(Tzfpw6[20]), .QN(n7278) );
  DFF_X1 Y7opw6_reg ( .D(n7997), .CK(SCLK), .Q(Tzfpw6[5]), .QN(n7339) );
  DFF_X1 Wlspw6_reg ( .D(n7987), .CK(SCLK), .Q(Tzfpw6[16]), .QN(n7362) );
  DFF_X1 Vrtpw6_reg ( .D(n7992), .CK(SCLK), .Q(Tzfpw6[10]), .QN(n7366) );
  DFF_X1 V0jpw6_reg ( .D(n7979), .CK(SCLK), .Q(Tzfpw6[12]), .QN(n7276) );
  DFF_X1 Uojbx6_reg ( .D(n7993), .CK(SCLK), .Q(Tzfpw6[9]), .QN(n7699) );
  DFF_X1 Ujxax6_reg ( .D(n7995), .CK(SCLK), .Q(Tzfpw6[7]), .QN(n7541) );
  DFF_X1 Tjkpw6_reg ( .D(n7982), .CK(SCLK), .Q(Tzfpw6[21]), .QN(n7290) );
  DFF_X1 T9kpw6_reg ( .D(n7990), .CK(SCLK), .Q(Tzfpw6[13]), .QN(n7288) );
  DFF_X1 Ss0qw6_reg ( .D(n7994), .CK(SCLK), .Q(Tzfpw6[8]), .QN(n7403) );
  DFF_X1 Rv7ax6_reg ( .D(n7996), .CK(SCLK), .Q(Tzfpw6[6]), .QN(n7445) );
  DFF_X1 Rfxax6_reg ( .D(n7989), .CK(SCLK), .Q(Tzfpw6[14]), .QN(n7539) );
  DFF_X1 Pt7ax6_reg ( .D(n7991), .CK(SCLK), .Q(Tzfpw6[11]), .QN(n7444) );
  DFF_X1 P0ibx6_reg ( .D(n7999), .CK(SCLK), .Q(Tzfpw6[3]), .QN(n7692) );
  DFF_X1 Oarpw6_reg ( .D(n8001), .CK(SCLK), .Q(Tzfpw6[1]), .QN(n7353) );
  DFF_X1 Nr7ax6_reg ( .D(n7984), .CK(SCLK), .Q(Tzfpw6[19]), .QN(n7443) );
  DFF_X1 Nbxax6_reg ( .D(n7988), .CK(SCLK), .Q(Tzfpw6[15]), .QN(n7537) );
  DFF_X1 N8rpw6_reg ( .D(n8002), .CK(SCLK), .Q(Tzfpw6[0]), .QN(n7352) );
  DFF_X1 N0xpw6_reg ( .D(n7985), .CK(SCLK), .Q(Tzfpw6[18]), .QN(n7391) );
  DFF_X1 Kzabx6_reg ( .D(n8000), .CK(SCLK), .Q(Tzfpw6[2]), .QN(n7642) );
  DFF_X1 Johbx6_reg ( .D(n7998), .CK(SCLK), .Q(Tzfpw6[4]), .QN(n7687) );
  DFF_X1 F9gbx6_reg ( .D(n7981), .CK(SCLK), .Q(Tzfpw6[22]), .QN(n7672) );
  DFF_X1 Coupw6_reg ( .D(n7980), .CK(SCLK), .Q(Tzfpw6[23]), .QN(n7369) );
  DFF_X1 Amupw6_reg ( .D(n7986), .CK(SCLK), .Q(Tzfpw6[17]), .QN(n7368) );
  DFFR_X1 Ok2bx6_reg ( .D(Ppthu6), .CK(SCLK), .RN(HRESETn), .QN(n6589) );
  DFFR_X1 Oi1bx6_reg ( .D(Nothu6), .CK(SCLK), .RN(HRESETn), .QN(n6587) );
  DFFR_X1 Ie1bx6_reg ( .D(Znthu6), .CK(SCLK), .RN(HRESETn), .QN(n6606) );
  DFFR_X1 Ca1bx6_reg ( .D(Snthu6), .CK(SCLK), .RN(HRESETn), .QN(n6594) );
  DFFR_X1 Sbyax6_reg ( .D(n2479), .CK(SCLK), .RN(HRESETn), .QN(n7549) );
  DFFR_X1 M13bx6_reg ( .D(n2486), .CK(SCLK), .RN(HRESETn), .QN(n6573) );
  DFFR_X1 At2bx6_reg ( .D(n2485), .CK(SCLK), .RN(HRESETn), .QN(n6580) );
  DFFR_X1 Z71bx6_reg ( .D(R2phu6), .CK(SCLK), .RN(HRESETn), .Q(n8106), .QN(
        n7583) );
  DFFR_X1 Lg1bx6_reg ( .D(Y2phu6), .CK(SCLK), .RN(HRESETn), .Q(n8166), .QN(
        n7585) );
  DFFR_X1 Rk1bx6_reg ( .D(K2phu6), .CK(SCLK), .RN(HRESETn), .QN(n7586) );
  DFFR_X1 Fc1bx6_reg ( .D(F3phu6), .CK(SCLK), .RN(HRESETn), .Q(n8170), .QN(
        n7584) );
  DFFR_X1 P33bx6_reg ( .D(Ezohu6), .CK(SCLK), .RN(HRESETn), .Q(n8296), .QN(
        n7598) );
  DFFR_X1 Dv2bx6_reg ( .D(Nwdpw6), .CK(SCLK), .RN(HRESETn), .Q(n3121), .QN(
        n7597) );
  DFFR_X1 Um1bx6_reg ( .D(Uothu6), .CK(SCLK), .RN(HRESETn), .Q(n8258), .QN(
        n6598) );
  DFFR_X1 Qaipw6_reg ( .D(Sgthu6), .CK(SCLK), .RN(HRESETn), .Q(n5175), .QN(
        n6593) );
  DFFR_X1 Gx2bx6_reg ( .D(Wpthu6), .CK(SCLK), .RN(HRESETn), .Q(n5148), .QN(
        n6602) );
  DFFR_X1 Ee3bx6_reg ( .D(Q6vhu6), .CK(SCLK), .RN(HRESETn), .Q(n5180), .QN(
        n6591) );
  DFFR_X1 Xo1bx6_reg ( .D(D2phu6), .CK(SCLK), .RN(HRESETn), .Q(n8259), .QN(
        n7587) );
  DFFR_X1 Tcipw6_reg ( .D(Jyohu6), .CK(SCLK), .RN(HRESETn), .Q(n2811), .QN(
        n7255) );
  DFFR_X1 Jz2bx6_reg ( .D(Lzohu6), .CK(SCLK), .RN(HRESETn), .Q(n5154), .QN(
        n6581) );
  DFFR_X1 Hg3bx6_reg ( .D(Cyohu6), .CK(SCLK), .RN(HRESETn), .Q(n5192), .QN(
        n7602) );
  DFFR_X1 Pdyax6_reg ( .D(Npghu6), .CK(SCLK), .RN(HRESETn), .Q(n2500), .QN(
        n7550) );
  DFFR_X1 W51bx6_reg ( .D(Gothu6), .CK(SCLK), .RN(HRESETn), .Q(n8105), .QN(
        n6579) );
  DFFR_X1 Woiax6_reg ( .D(Bpthu6), .CK(SCLK), .RN(HRESETn), .Q(n8249) );
  DFFR_X1 Y93bx6_reg ( .D(J6vhu6), .CK(SCLK), .RN(HRESETn), .Q(n8288) );
  DFFR_X1 Vyfbx6_reg ( .D(Uuuhu6), .CK(SCLK), .RN(HRESETn), .Q(n8202) );
  DFFR_X1 Pgjbx6_reg ( .D(Lnthu6), .CK(SCLK), .RN(HRESETn), .Q(n8290) );
  DFFR_X1 L3bbx6_reg ( .D(Jmthu6), .CK(SCLK), .RN(HRESETn), .Q(n5216) );
  DFFR_X1 Ki3bx6_reg ( .D(Hsthu6), .CK(SCLK), .RN(HRESETn), .Q(n8289) );
  DFFR_X1 S32bx6_reg ( .D(Xsuhu6), .CK(SCLK), .RN(HRESETn), .Q(n5128) );
  DFFR_X1 Om3bx6_reg ( .D(Vsthu6), .CK(SCLK), .RN(HRESETn), .Q(n8238) );
  DFFR_X1 Kshbx6_reg ( .D(Trthu6), .CK(SCLK), .RN(HRESETn), .Q(n5209) );
  DFFR_X1 Gv1bx6_reg ( .D(Zgthu6), .CK(SCLK), .RN(HRESETn), .Q(n5129) );
  DFFR_X1 Ar1bx6_reg ( .D(Vruhu6), .CK(SCLK), .RN(HRESETn), .Q(n8286) );
  DFFR_X1 Y72bx6_reg ( .D(Cmthu6), .CK(SCLK), .RN(HRESETn), .Q(n3268) );
  DFFR_X1 Uo2bx6_reg ( .D(Pvuhu6), .CK(SCLK), .RN(HRESETn), .Q(n8293) );
  DFFR_X1 Sq3bx6_reg ( .D(Enthu6), .CK(SCLK), .RN(HRESETn), .Q(n5198) );
  DFFR_X1 S11bx6_reg ( .D(Mivhu6), .CK(SCLK), .RN(HRESETn), .Q(n4839) );
  DFFR_X1 Mz1bx6_reg ( .D(Jsuhu6), .CK(SCLK), .RN(HRESETn), .Q(n5134) );
  DFFR_X1 Jp9bx6_reg ( .D(Osthu6), .CK(SCLK), .RN(HRESETn), .Q(n4281) );
  DFFR_X1 Ig2bx6_reg ( .D(Ztuhu6), .CK(SCLK), .RN(HRESETn), .Q(n8287) );
  DFFR_X1 Eghbx6_reg ( .D(Asthu6), .CK(SCLK), .RN(HRESETn), .Q(n5193) );
  DFFR_X1 Cc2bx6_reg ( .D(Ltuhu6), .CK(SCLK), .RN(HRESETn), .Q(n8226) );
  DFFR_X1 S53bx6_reg ( .D(Kqthu6), .CK(SCLK), .RN(HRESETn), .Q(n8279), .QN(
        n6584) );
  DFFR_X1 Rm2bx6_reg ( .D(n2646), .CK(SCLK), .RN(HRESETn), .QN(n7595) );
  DFFR_X1 Us3bx6_reg ( .D(n7266), .CK(SCLK), .RN(HRESETn), .Q(n4010), .QN(
        n7604) );
  DFFR_X1 Y0gbx6_reg ( .D(Zzohu6), .CK(SCLK), .RN(HRESETn), .Q(n8203), .QN(
        n7669) );
  DFFR_X1 Qo3bx6_reg ( .D(n7272), .CK(SCLK), .RN(HRESETn), .Q(n8239), .QN(
        n6582) );
  DFFR_X1 Fe2bx6_reg ( .D(n7260), .CK(SCLK), .RN(HRESETn), .Q(n8227), .QN(
        n7593) );
  DFFR_X1 Dt1bx6_reg ( .D(n7265), .CK(SCLK), .RN(HRESETn), .Q(n3310), .QN(
        n7588) );
  DFFR_X1 P12bx6_reg ( .D(n7264), .CK(SCLK), .RN(HRESETn), .Q(n4061), .QN(
        n7590) );
  DFFR_X1 Lr9bx6_reg ( .D(n7273), .CK(SCLK), .RN(HRESETn), .Q(n4293), .QN(
        n6578) );
  DFFR_X1 Aa2bx6_reg ( .D(n7254), .CK(SCLK), .RN(HRESETn), .Q(n3276), .QN(
        n7592) );
  DFFR_X1 U31bx6_reg ( .D(n7268), .CK(SCLK), .RN(HRESETn), .Q(n4001), .QN(
        n6575) );
  DFFR_X1 Rijbx6_reg ( .D(Uwdpw6), .CK(SCLK), .RN(HRESETn), .Q(n3930), .QN(
        n7696) );
  DFFR_X1 Xq2bx6_reg ( .D(n7270), .CK(SCLK), .RN(HRESETn), .Q(n8294), .QN(
        n7596) );
  DFFR_X1 Muhbx6_reg ( .D(n7263), .CK(SCLK), .RN(HRESETn), .Q(n5210), .QN(
        n7689) );
  DFFR_X1 Bc3bx6_reg ( .D(Qyohu6), .CK(SCLK), .RN(HRESETn), .Q(n3037), .QN(
        n7601) );
  DFFR_X1 N5bbx6_reg ( .D(V4phu6), .CK(SCLK), .RN(HRESETn), .Q(n3030), .QN(
        n7645) );
  DFFR_X1 Jx1bx6_reg ( .D(n7267), .CK(SCLK), .RN(HRESETn), .Q(n4005), .QN(
        n7589) );
  DFFR_X1 Gihbx6_reg ( .D(H4phu6), .CK(SCLK), .RN(HRESETn), .Q(n5197), .QN(
        n7684) );
  DFFR_X1 V52bx6_reg ( .D(n7262), .CK(SCLK), .RN(HRESETn), .Q(n3870), .QN(
        n7591) );
  DFFR_X1 Li2bx6_reg ( .D(n7269), .CK(SCLK), .RN(HRESETn), .Q(n3669), .QN(
        n7594) );
  DFFR_X1 V73bx6_reg ( .D(n2651), .CK(SCLK), .RN(HRESETn), .Q(n8280), .QN(
        n7599) );
  DFFR_X1 Yxrpw6_reg ( .D(n7271), .CK(SCLK), .RN(HRESETn), .Q(n8250), .QN(
        n7357) );
  DFFR_X1 T2kbx6_reg ( .D(n8003), .CK(SCLK), .RN(HRESETn), .QN(n7702) );
  DFFR_X1 Zdtpw6_reg ( .D(n7952), .CK(SCLK), .RN(HRESETn), .Q(n3617), .QN(
        n7364) );
  DFFR_X1 Z9opw6_reg ( .D(J4xhu6), .CK(SCLK), .RN(HRESETn), .Q(n2502), .QN(
        n6684) );
  DFFR_X1 Cokbx6_reg ( .D(n6917), .CK(SCLK), .RN(HRESETn), .Q(n221), .QN(n6685) );
  DFFR_X1 Vzjpw6_reg ( .D(Fivhu6), .CK(SCLK), .RN(HRESETn), .Q(n2233), .QN(
        n7285) );
  DFFS_X1 Fnnpw6_reg ( .D(n7256), .CK(SCLK), .SN(HRESETn), .Q(n4674), .QN(
        n6682) );
  DFFS_X1 L4lax6_reg ( .D(Wfphu6), .CK(SCLK), .SN(HRESETn), .Q(n3533), .QN(
        n7531) );
  DFF_X1 W8hbx6_reg ( .D(Yhvhu6), .CK(SCLK), .QN(n7682) );
  DFF_X1 Zqiax6_reg ( .D(n7862), .CK(SCLK), .Q(n3538), .QN(n7498) );
  DFF_X1 Ysiax6_reg ( .D(n7863), .CK(SCLK), .Q(n3540), .QN(n7499) );
  DFF_X1 Xuiax6_reg ( .D(n7864), .CK(SCLK), .Q(n3543), .QN(n7500) );
  DFF_X1 Wyiax6_reg ( .D(n7866), .CK(SCLK), .Q(n3545), .QN(n7502) );
  DFF_X1 Wwiax6_reg ( .D(n7865), .CK(SCLK), .Q(n3544), .QN(n7501) );
  DFF_X1 W2jax6_reg ( .D(n7868), .CK(SCLK), .Q(n3534), .QN(n7504) );
  DFF_X1 W0jax6_reg ( .D(n7867), .CK(SCLK), .Q(n3546), .QN(n7503) );
  DFF_X1 E8iax6_reg ( .D(n7861), .CK(SCLK), .Q(n3535), .QN(n7496) );
  DFF_X1 Xiipw6_reg ( .D(n7858), .CK(SCLK), .Q(n4855), .QN(n7258) );
  DFF_X1 Xdspw6_reg ( .D(n7869), .CK(SCLK), .Q(n2232), .QN(n7358) );
  DFF_X1 T5mpw6_reg ( .D(n7856), .CK(SCLK), .Q(n4841), .QN(n7324) );
  DFF_X1 Jpmpw6_reg ( .D(n7857), .CK(SCLK), .Q(n3065), .QN(n7328) );
  DFF_X1 G2iax6_reg ( .D(n7859), .CK(SCLK), .QN(n7494) );
  DFF_X1 F4iax6_reg ( .D(n7860), .CK(SCLK), .QN(n7495) );
  DFFR_X1 T0ipw6_reg ( .D(O5ohu6), .CK(SWCLKTCK), .RN(Fmdhu6), .Q(n1817), .QN(
        n7249) );
  DFFR_X1 Qwfax6_reg ( .D(S3ohu6), .CK(SWCLKTCK), .RN(Fmdhu6), .QN(n6604) );
  DFFR_X1 Cjqpw6_reg ( .D(n7829), .CK(SWCLKTCK), .RN(Fmdhu6), .Q(n4041), .QN(
        n7348) );
  DFFR_X1 Pmlpw6_reg ( .D(n8054), .CK(SWCLKTCK), .RN(Fmdhu6), .Q(n4016), .QN(
        n7315) );
  DFFR_X1 Jflpw6_reg ( .D(n8052), .CK(SWCLKTCK), .RN(Fmdhu6), .Q(n4024), .QN(
        n7311) );
  DFFR_X1 Gylpw6_reg ( .D(n7252), .CK(SWCLKTCK), .RN(Fmdhu6), .QN(n6622) );
  DFFR_X1 Yklpw6_reg ( .D(n7840), .CK(SWCLKTCK), .RN(Fmdhu6), .Q(n3201), .QN(
        n7314) );
  DFFR_X1 Ryfax6_reg ( .D(n7831), .CK(SWCLKTCK), .RN(Fmdhu6), .Q(n4136), .QN(
        n7482) );
  DFFR_X1 Oulpw6_reg ( .D(Sqxhu6), .CK(SWCLKTCK), .RN(Fmdhu6), .Q(n4036), .QN(
        n7320) );
  DFFR_X1 A5ipw6_reg ( .D(n7835), .CK(SWCLKTCK), .RN(Fmdhu6), .Q(n3242), .QN(
        n6673) );
  DFFR_X1 I0opw6_reg ( .D(n7832), .CK(SWCLKTCK), .RN(Fmdhu6), .Q(n3233), .QN(
        n7336) );
  DFFR_X1 Ry2qw6_reg ( .D(n7836), .CK(SWCLKTCK), .RN(Fmdhu6), .QN(n7417) );
  DFFR_X1 B7lpw6_reg ( .D(Fwohu6), .CK(SWCLKTCK), .RN(Fmdhu6), .Q(n4138), .QN(
        n7305) );
  DFFR_X1 T82qw6_reg ( .D(n7251), .CK(SWCLKTCK), .RN(Fmdhu6), .Q(n4038), .QN(
        n6608) );
  DFFR_X1 Hpcbx6_reg ( .D(Mgxhu6), .CK(SWCLKTCK), .RN(Fmdhu6), .QN(n7656) );
  DFFR_X1 Ehqpw6_reg ( .D(Fgxhu6), .CK(SWCLKTCK), .RN(Fmdhu6), .Q(n4040), .QN(
        n7347) );
  DFFR_X1 Kwlpw6_reg ( .D(Tgxhu6), .CK(SWCLKTCK), .RN(Fmdhu6), .QN(n7321) );
  DFFR_X1 Qynpw6_reg ( .D(Hvxhu6), .CK(SWCLKTCK), .RN(Fmdhu6), .Q(n3127), .QN(
        n7335) );
  DFFR_X1 Bclpw6_reg ( .D(n7837), .CK(SWCLKTCK), .RN(Fmdhu6), .Q(n4028), .QN(
        n7309) );
  DFFS_X1 Kalpw6_reg ( .D(n8053), .CK(SWCLKTCK), .SN(Fmdhu6), .Q(n4029), .QN(
        n7308) );
  DFFS_X1 Ahlpw6_reg ( .D(n7839), .CK(SWCLKTCK), .SN(n956), .QN(n7312) );
  DFFS_X1 Sdlpw6_reg ( .D(n7838), .CK(SWCLKTCK), .SN(n956), .Q(n3212), .QN(
        n7310) );
  DFFS_X1 Rilpw6_reg ( .D(n3139), .CK(SWCLKTCK), .SN(n956), .Q(n4022), .QN(
        n7313) );
  DFF_X1 Krlpw6_reg ( .D(n7725), .CK(SWCLKTCK), .Q(n4034), .QN(n7318) );
  DFF_X1 Zslpw6_reg ( .D(n7724), .CK(SWCLKTCK), .Q(n4035), .QN(n7319) );
  DFF_X1 Golpw6_reg ( .D(Yvohu6), .CK(SWCLKTCK), .Q(n4032), .QN(n7316) );
  DFF_X1 Vplpw6_reg ( .D(Rvohu6), .CK(SWCLKTCK), .Q(n4033), .QN(n7317) );
  DFF_X1 Z73qw6_reg ( .D(n3129), .CK(SWCLKTCK), .Q(n3884), .QN(n7420) );
  DFF_X1 Stkpw6_reg ( .D(n3128), .CK(SWCLKTCK), .QN(n6625) );
  DFF_X1 Li7ax6_reg ( .D(n3009), .CK(SWCLKTCK), .QN(n7439) );
  DFF_X1 J4cbx6_reg ( .D(n7294), .CK(SWCLKTCK), .QN(n7652) );
  DFF_X1 Wq8ax6_reg ( .D(n8042), .CK(SWCLKTCK), .QN(n6619) );
  DFF_X1 Sddbx6_reg ( .D(n8045), .CK(SWCLKTCK), .QN(n6610) );
  DFF_X1 S2cbx6_reg ( .D(n8047), .CK(SWCLKTCK), .QN(n7651) );
  DFF_X1 Kn2qw6_reg ( .D(n8046), .CK(SWCLKTCK), .QN(n6624) );
  DFF_X1 Kadbx6_reg ( .D(n8020), .CK(SWCLKTCK), .QN(n6623) );
  DFF_X1 Jfdbx6_reg ( .D(n8044), .CK(SWCLKTCK), .QN(n6611) );
  DFF_X1 Hlwpw6_reg ( .D(n8043), .CK(SWCLKTCK), .QN(n6615) );
  DFF_X1 Yzlpw6_reg ( .D(n8051), .CK(SWCLKTCK), .Q(n4042), .QN(n7322) );
  DFF_X1 L0ypw6_reg ( .D(n8041), .CK(SWCLKTCK), .QN(n6621) );
  DFF_X1 Bx2qw6_reg ( .D(n8037), .CK(SWCLKTCK), .QN(n7416) );
  DFF_X1 Xf8ax6_reg ( .D(n7300), .CK(SWCLKTCK), .QN(n6617) );
  DFF_X1 Ufbbx6_reg ( .D(n7298), .CK(SWCLKTCK), .QN(n6614) );
  DFF_X1 Qj1qw6_reg ( .D(n7303), .CK(SWCLKTCK), .QN(n6671) );
  DFF_X1 Qa1qw6_reg ( .D(n7304), .CK(SWCLKTCK), .QN(n6672) );
  DFF_X1 Puwpw6_reg ( .D(n7297), .CK(SWCLKTCK), .QN(n6613) );
  DFF_X1 Oh8ax6_reg ( .D(n7301), .CK(SWCLKTCK), .QN(n6618) );
  DFF_X1 Ldvpw6_reg ( .D(n7296), .CK(SWCLKTCK), .QN(n6612) );
  DFF_X1 Gw6bx6_reg ( .D(n7302), .CK(SWCLKTCK), .QN(n6620) );
  DFF_X1 E97ax6_reg ( .D(n7299), .CK(SWCLKTCK), .QN(n6616) );
  DFF_X1 Bcdbx6_reg ( .D(n7295), .CK(SWCLKTCK), .QN(n6609) );
  DFF_X1 Y8lpw6_reg ( .D(n7834), .CK(SWCLKTCK), .Q(n4027), .QN(n7306) );
  DFF_X1 Zgfax6_reg ( .D(n3130), .CK(SWCLKTCK), .QN(n7477) );
  DFF_X1 W6ipw6_reg ( .D(n7842), .CK(SWCLKTCK), .QN(n7253) );
  DFF_X1 D2opw6_reg ( .D(n8039), .CK(SWCLKTCK), .QN(n7337) );
  DFF_X1 L5lpw6_reg ( .D(n7843), .CK(SWCLKTCK), .QN(n7293) );
  DFF_X1 Okfax6_reg ( .D(Isxhu6), .CK(SWCLKTCK), .QN(n7478) );
  DFF_X1 Lhbbx6_reg ( .D(n7216), .CK(SWCLKTCK), .QN(n6905) );
  DFF_X1 D2rpw6_reg ( .D(n7217), .CK(SWCLKTCK), .QN(n6882) );
  DFF_X1 Q89bx6_reg ( .D(n7215), .CK(SWCLKTCK), .QN(n6900) );
  DFF_X1 Nmfax6_reg ( .D(Xpxhu6), .CK(SWCLKTCK), .QN(n7479) );
  DFF_X1 J0gax6_reg ( .D(n7240), .CK(SWCLKTCK), .QN(n6597) );
  DFF_X1 Nv3qw6_reg ( .D(n7243), .CK(SWCLKTCK), .QN(n6727) );
  DFF_X1 Gnqpw6_reg ( .D(n7214), .CK(SWCLKTCK), .QN(n6569) );
  DFF_X1 H0ebx6_reg ( .D(n7248), .CK(SWCLKTCK), .QN(n6907) );
  DFF_X1 C2ypw6_reg ( .D(n7247), .CK(SWCLKTCK), .QN(n6750) );
  DFF_X1 Bp2qw6_reg ( .D(n7246), .CK(SWCLKTCK), .Q(n3618), .QN(n6915) );
  DFF_X1 Liabx6_reg ( .D(n7245), .CK(SWCLKTCK), .QN(n6708) );
  DFF_X1 Yzqpw6_reg ( .D(n7242), .CK(SWCLKTCK), .Q(n3879), .QN(n6884) );
  DFF_X1 L03qw6_reg ( .D(n7244), .CK(SWCLKTCK), .Q(n4049), .QN(n6885) );
  DFF_X1 Nrqpw6_reg ( .D(n7221), .CK(SWCLKTCK), .QN(n6572) );
  DFF_X1 M8ipw6_reg ( .D(n7228), .CK(SWCLKTCK), .QN(n6872) );
  DFF_X1 I4rpw6_reg ( .D(n7224), .CK(SWCLKTCK), .QN(n6910) );
  DFF_X1 Gpqpw6_reg ( .D(n7236), .CK(SWCLKTCK), .QN(n6592) );
  DFF_X1 Bk7ax6_reg ( .D(n7218), .CK(SWCLKTCK), .QN(n6898) );
  DFF_X1 Xx6bx6_reg ( .D(n7237), .CK(SWCLKTCK), .QN(n6756) );
  DFF_X1 Ns8ax6_reg ( .D(n7229), .CK(SWCLKTCK), .QN(n6875) );
  DFF_X1 Fj8ax6_reg ( .D(n7219), .CK(SWCLKTCK), .QN(n6908) );
  DFF_X1 Ojebx6_reg ( .D(n7238), .CK(SWCLKTCK), .QN(n6741) );
  DFF_X1 Ahdbx6_reg ( .D(n7223), .CK(SWCLKTCK), .QN(n6718) );
  DFF_X1 Urgbx6_reg ( .D(n7230), .CK(SWCLKTCK), .QN(n6912) );
  DFF_X1 Jvkpw6_reg ( .D(n7220), .CK(SWCLKTCK), .Q(n3388), .QN(n6894) );
  DFF_X1 Gwwpw6_reg ( .D(n7241), .CK(SWCLKTCK), .QN(n6903) );
  DFF_X1 Cfvpw6_reg ( .D(n7232), .CK(SWCLKTCK), .QN(n6904) );
  DFF_X1 Va7ax6_reg ( .D(n7235), .CK(SWCLKTCK), .QN(n6766) );
  DFF_X1 Gc1qw6_reg ( .D(n7231), .CK(SWCLKTCK), .QN(n6902) );
  DFF_X1 Gl1qw6_reg ( .D(n7222), .CK(SWCLKTCK), .Q(n3922), .QN(n6901) );
  DFF_X1 Ra2qw6_reg ( .D(n7233), .CK(SWCLKTCK), .QN(n6897) );
  DFF_X1 A6cbx6_reg ( .D(Qixhu6), .CK(SWCLKTCK), .QN(n7653) );
  DFF_X1 Drcbx6_reg ( .D(n7227), .CK(SWCLKTCK), .QN(n6692) );
  DFF_X1 Ymwpw6_reg ( .D(n7226), .CK(SWCLKTCK), .QN(n6906) );
  DFF_X1 O1mpw6_reg ( .D(n7239), .CK(SWCLKTCK), .QN(n6889) );
  DFF_X1 T3opw6_reg ( .D(n7225), .CK(SWCLKTCK), .Q(n4409), .QN(n6911) );
  DFF_X1 P93qw6_reg ( .D(n7234), .CK(SWCLKTCK), .Q(n4139), .QN(n6887) );
  DFF_X1 Wt3qw6_reg ( .D(n7833), .CK(SWCLKTCK), .QN(n7431) );
  DFF_X1 Zwnpw6_reg ( .D(n8050), .CK(SWCLKTCK), .QN(n7334) );
  DFF_X1 Nfqpw6_reg ( .D(n8048), .CK(SWCLKTCK), .QN(n7346) );
  DFF_X1 C72qw6_reg ( .D(n8049), .CK(SWCLKTCK), .QN(n7409) );
  DFFS_X2 Xbopw6_reg ( .D(n1855), .CK(SCLK), .SN(HRESETn), .Q(SLEEPHOLDACKn), 
        .QN(n7340) );
  INV_X1 U3 ( .A(1'b1), .ZN(WICENACK) );
  INV_X1 U5 ( .A(1'b1), .ZN(WICSENSE[0]) );
  INV_X1 U7 ( .A(1'b1), .ZN(WICSENSE[1]) );
  INV_X1 U9 ( .A(1'b1), .ZN(WICSENSE[2]) );
  INV_X1 U15 ( .A(1'b1), .ZN(WICSENSE[3]) );
  INV_X1 U17 ( .A(1'b1), .ZN(WICSENSE[4]) );
  INV_X1 U19 ( .A(1'b1), .ZN(WICSENSE[5]) );
  INV_X1 U21 ( .A(1'b1), .ZN(WICSENSE[6]) );
  INV_X1 U23 ( .A(1'b1), .ZN(WICSENSE[7]) );
  INV_X1 U25 ( .A(1'b1), .ZN(WICSENSE[8]) );
  INV_X1 U27 ( .A(1'b1), .ZN(WICSENSE[9]) );
  INV_X1 U29 ( .A(1'b1), .ZN(WICSENSE[10]) );
  INV_X1 U31 ( .A(1'b1), .ZN(WICSENSE[11]) );
  INV_X1 U33 ( .A(1'b1), .ZN(WICSENSE[12]) );
  INV_X1 U35 ( .A(1'b1), .ZN(WICSENSE[13]) );
  INV_X1 U37 ( .A(1'b1), .ZN(WICSENSE[14]) );
  INV_X1 U39 ( .A(1'b1), .ZN(WICSENSE[15]) );
  INV_X1 U42 ( .A(1'b1), .ZN(WICSENSE[16]) );
  INV_X1 U44 ( .A(1'b1), .ZN(WICSENSE[17]) );
  INV_X1 U46 ( .A(1'b1), .ZN(WICSENSE[18]) );
  INV_X1 U48 ( .A(1'b1), .ZN(WICSENSE[19]) );
  INV_X1 U50 ( .A(1'b1), .ZN(WICSENSE[20]) );
  INV_X1 U52 ( .A(1'b1), .ZN(WICSENSE[21]) );
  INV_X1 U54 ( .A(1'b1), .ZN(WICSENSE[22]) );
  INV_X1 U56 ( .A(1'b1), .ZN(WICSENSE[23]) );
  INV_X1 U58 ( .A(1'b1), .ZN(WICSENSE[24]) );
  INV_X1 U60 ( .A(1'b1), .ZN(WICSENSE[25]) );
  INV_X1 U63 ( .A(1'b1), .ZN(WICSENSE[26]) );
  INV_X1 U65 ( .A(1'b1), .ZN(WICSENSE[27]) );
  INV_X1 U67 ( .A(1'b1), .ZN(WICSENSE[28]) );
  INV_X1 U69 ( .A(1'b1), .ZN(WICSENSE[29]) );
  INV_X1 U71 ( .A(1'b1), .ZN(WICSENSE[30]) );
  INV_X1 U73 ( .A(1'b1), .ZN(WICSENSE[31]) );
  INV_X1 U75 ( .A(1'b1), .ZN(WICSENSE[32]) );
  INV_X1 U77 ( .A(1'b1), .ZN(WICSENSE[33]) );
  INV_X1 U80 ( .A(1'b1), .ZN(WAKEUP) );
  INV_X1 U82 ( .A(1'b1), .ZN(nTDOEN) );
  INV_X1 U84 ( .A(1'b1), .ZN(TDO) );
  INV_X1 U86 ( .A(1'b1), .ZN(HTRANS[0]) );
  INV_X1 U88 ( .A(1'b1), .ZN(HSIZE[2]) );
  INV_X1 U90 ( .A(1'b0), .ZN(HPROT[1]) );
  INV_X1 U92 ( .A(1'b1), .ZN(HMASTLOCK) );
  INV_X1 U94 ( .A(1'b1), .ZN(HBURST[0]) );
  INV_X1 U96 ( .A(1'b1), .ZN(HBURST[1]) );
  INV_X1 U98 ( .A(1'b1), .ZN(HBURST[2]) );
  AND2_X1 U100 ( .A1(n5236), .A2(n221), .ZN(SLEEPING) );
  AOI211_X1 U101 ( .C1(n6238), .C2(n6217), .A(n6632), .B(n6581), .ZN(n6216) );
  NOR2_X1 U104 ( .A1(n4451), .A2(n6601), .ZN(n4426) );
  NAND2_X1 U105 ( .A1(n7461), .A2(n2307), .ZN(Msmhu6) );
  NAND2_X1 U106 ( .A1(n7465), .A2(n2333), .ZN(Oakhu6) );
  AOI22_X1 U107 ( .A1(n6193), .A2(n6194), .B1(n6171), .B2(n6195), .ZN(n5309)
         );
  NOR3_X1 U108 ( .A1(n4160), .A2(n4410), .A3(n4182), .ZN(n1856) );
  NOR2_X1 U109 ( .A1(n5112), .A2(vis_ipsr_o[1]), .ZN(n5867) );
  NOR2_X1 U111 ( .A1(vis_ipsr_o[0]), .A2(vis_ipsr_o[1]), .ZN(n5243) );
  AOI221_X1 U112 ( .B1(n172), .B2(HADDR[7]), .C1(n173), .C2(HADDR[6]), .A(
        HADDR[9]), .ZN(n171) );
  NOR2_X1 U114 ( .A1(n266), .A2(n538), .ZN(n1620) );
  NOR3_X1 U115 ( .A1(n491), .A2(n529), .A3(n522), .ZN(n1455) );
  NOR2_X1 U116 ( .A1(n254), .A2(n7283), .ZN(n435) );
  AOI221_X1 U117 ( .B1(n3365), .B2(n4717), .C1(n4691), .C2(HRDATA[6]), .A(
        n5527), .ZN(n4522) );
  AOI222_X1 U118 ( .A1(n3359), .A2(n3725), .B1(n1219), .B2(n4705), .C1(n4691), 
        .C2(HRDATA[8]), .ZN(n4393) );
  AOI222_X1 U119 ( .A1(n2391), .A2(n3725), .B1(n4691), .B2(HRDATA[15]), .C1(
        n837), .C2(n4705), .ZN(n4344) );
  AOI221_X1 U120 ( .B1(n2826), .B2(n4705), .C1(n3371), .C2(n4690), .A(n5338), 
        .ZN(n4593) );
  OAI211_X1 U121 ( .C1(n2722), .C2(n3081), .A(n6038), .B(n5576), .ZN(n4269) );
  NOR3_X1 U122 ( .A1(n4410), .A2(n7371), .A3(n4160), .ZN(n1325) );
  NOR3_X1 U123 ( .A1(n3913), .A2(n7388), .A3(n3882), .ZN(n1182) );
  NOR2_X1 U124 ( .A1(n485), .A2(n7283), .ZN(n2562) );
  OAI21_X1 U125 ( .B1(n7533), .B2(n2439), .A(n7491), .ZN(n3876) );
  OAI21_X1 U126 ( .B1(n2693), .B2(n7533), .A(n7491), .ZN(n4906) );
  NOR2_X1 U127 ( .A1(n254), .A2(n237), .ZN(n474) );
  NOR2_X1 U128 ( .A1(n2193), .A2(n7383), .ZN(n2089) );
  NOR2_X1 U129 ( .A1(n2200), .A2(n7383), .ZN(n2105) );
  NOR2_X1 U130 ( .A1(n2199), .A2(n7383), .ZN(n2101) );
  NOR2_X1 U131 ( .A1(n2198), .A2(n7383), .ZN(n2099) );
  NOR2_X1 U132 ( .A1(n2194), .A2(n7383), .ZN(n2097) );
  NOR2_X1 U133 ( .A1(n2197), .A2(n7383), .ZN(n2095) );
  NOR2_X1 U134 ( .A1(n2196), .A2(n7383), .ZN(n2093) );
  NOR2_X1 U135 ( .A1(n2195), .A2(n7383), .ZN(n2091) );
  INV_X1 U136 ( .A(Nxkbx6[30]), .ZN(n1575) );
  INV_X1 U137 ( .A(Nxkbx6[29]), .ZN(n1581) );
  INV_X1 U138 ( .A(Nxkbx6[28]), .ZN(n1590) );
  INV_X1 U139 ( .A(Nxkbx6[27]), .ZN(n1597) );
  INV_X1 U140 ( .A(Nxkbx6[26]), .ZN(n1604) );
  INV_X1 U141 ( .A(Nxkbx6[25]), .ZN(n1608) );
  INV_X1 U142 ( .A(Nxkbx6[5]), .ZN(n1795) );
  INV_X1 U143 ( .A(Nxkbx6[3]), .ZN(n1804) );
  INV_X1 U144 ( .A(Nxkbx6[10]), .ZN(n1770) );
  INV_X1 U145 ( .A(Nxkbx6[14]), .ZN(n1717) );
  INV_X1 U146 ( .A(Nxkbx6[15]), .ZN(n1696) );
  INV_X1 U147 ( .A(Nxkbx6[8]), .ZN(n1783) );
  INV_X1 U148 ( .A(Nxkbx6[12]), .ZN(n1764) );
  INV_X1 U149 ( .A(Nxkbx6[13]), .ZN(n1719) );
  INV_X1 U150 ( .A(Nxkbx6[9]), .ZN(n1775) );
  INV_X1 U151 ( .A(Nxkbx6[11]), .ZN(n1767) );
  INV_X1 U152 ( .A(Nxkbx6[4]), .ZN(n1801) );
  INV_X1 U153 ( .A(Nxkbx6[7]), .ZN(n1786) );
  INV_X1 U154 ( .A(Nxkbx6[2]), .ZN(n1809) );
  XOR2_X1 U155 ( .A(n6914), .B(n6913), .Z(n1371) );
  AND2_X1 U156 ( .A1(n1365), .A2(n3923), .ZN(n222) );
  AND2_X1 U157 ( .A1(n5544), .A2(n1325), .ZN(n226) );
  AND3_X1 U158 ( .A1(n5723), .A2(n4394), .A3(n5724), .ZN(n229) );
  OR2_X1 U159 ( .A1(n5236), .A2(n7340), .ZN(n230) );
  AND4_X1 U160 ( .A1(n914), .A2(n354), .A3(n3258), .A4(n4844), .ZN(n233) );
  AND2_X1 U161 ( .A1(n906), .A2(n3568), .ZN(n234) );
  AND3_X1 U162 ( .A1(n7305), .A2(n3158), .A3(n2177), .ZN(n236) );
  AND2_X1 U163 ( .A1(n1293), .A2(n1108), .ZN(n239) );
  OR4_X1 U164 ( .A1(n5635), .A2(n5636), .A3(n5637), .A4(n5638), .ZN(n242) );
  OR3_X1 U165 ( .A1(n7355), .A2(n7279), .A3(n4598), .ZN(n243) );
  AND2_X1 U166 ( .A1(n7312), .A2(n4016), .ZN(n244) );
  OR2_X1 U167 ( .A1(n989), .A2(n7412), .ZN(n247) );
  OR2_X1 U168 ( .A1(n1004), .A2(n7412), .ZN(n249) );
  OR2_X1 U169 ( .A1(n985), .A2(n7412), .ZN(n250) );
  OR2_X1 U170 ( .A1(n1006), .A2(n7412), .ZN(n253) );
  OR2_X1 U171 ( .A1(n377), .A2(n380), .ZN(HADDR[18]) );
  OR2_X1 U172 ( .A1(n373), .A2(n376), .ZN(HADDR[19]) );
  OR2_X1 U173 ( .A1(n370), .A2(n371), .ZN(HADDR[24]) );
  INV_X1 U174 ( .A(n365), .ZN(HADDR[3]) );
  XOR2_X1 U175 ( .A(\add_3107/B[1] ), .B(Tnhpw6[0]), .Z(n277) );
  XOR2_X1 U176 ( .A(Jshpw6[4]), .B(n424), .Z(n279) );
  XOR2_X1 U177 ( .A(Jshpw6[6]), .B(n423), .Z(n281) );
  XOR2_X1 U178 ( .A(Jshpw6[5]), .B(n422), .Z(n283) );
  XOR2_X1 U179 ( .A(Jshpw6[8]), .B(n421), .Z(n285) );
  XOR2_X1 U180 ( .A(Tnhpw6[3]), .B(\add_3107/carry[4] ), .Z(n287) );
  XOR2_X1 U181 ( .A(Jshpw6[7]), .B(n425), .Z(n288) );
  XOR2_X1 U182 ( .A(Jshpw6[9]), .B(n430), .Z(n290) );
  INV_X1 U183 ( .A(n8373), .ZN(n293) );
  INV_X1 U184 ( .A(n293), .ZN(HADDR[21]) );
  OAI22_X1 U185 ( .A1(n952), .A2(n1631), .B1(n7664), .B2(n946), .ZN(n8373) );
  INV_X1 U186 ( .A(n8372), .ZN(n298) );
  INV_X1 U187 ( .A(n298), .ZN(HADDR[25]) );
  OAI22_X1 U188 ( .A1(n952), .A2(n1603), .B1(n7693), .B2(n950), .ZN(n8372) );
  INV_X1 U189 ( .A(n8371), .ZN(n303) );
  INV_X1 U190 ( .A(n303), .ZN(HADDR[26]) );
  OAI22_X1 U191 ( .A1(n952), .A2(n1596), .B1(n7655), .B2(n950), .ZN(n8371) );
  INV_X1 U192 ( .A(n8370), .ZN(n308) );
  INV_X1 U193 ( .A(n308), .ZN(HADDR[27]) );
  OAI22_X1 U194 ( .A1(n952), .A2(n1582), .B1(n7657), .B2(n950), .ZN(n8370) );
  INV_X1 U195 ( .A(n8369), .ZN(n313) );
  INV_X1 U196 ( .A(n313), .ZN(HADDR[28]) );
  OAI22_X1 U197 ( .A1(n1580), .A2(n952), .B1(n7488), .B2(n950), .ZN(n8369) );
  INV_X1 U198 ( .A(n8375), .ZN(n316) );
  INV_X1 U199 ( .A(n316), .ZN(HADDR[6]) );
  AOI22_X1 U200 ( .A1(n1785), .A2(n941), .B1(n955), .B2(n7632), .ZN(n8375) );
  INV_X1 U201 ( .A(n8384), .ZN(n320) );
  INV_X1 U202 ( .A(n320), .ZN(HWDATA[15]) );
  OAI222_X1 U203 ( .A1(n6766), .A2(n670), .B1(n4180), .B2(n3874), .C1(n2478), 
        .C2(n3876), .ZN(n8384) );
  INV_X1 U204 ( .A(n8376), .ZN(n323) );
  INV_X1 U205 ( .A(n323), .ZN(HADDR[5]) );
  AOI22_X1 U206 ( .A1(n1788), .A2(n941), .B1(n955), .B2(n7423), .ZN(n8376) );
  INV_X1 U207 ( .A(n8374), .ZN(n328) );
  INV_X1 U208 ( .A(n328), .ZN(HADDR[10]) );
  AOI22_X1 U209 ( .A1(n1766), .A2(n941), .B1(n955), .B2(n7397), .ZN(n8374) );
  INV_X1 U210 ( .A(n8385), .ZN(n332) );
  INV_X1 U211 ( .A(n332), .ZN(HWDATA[14]) );
  OAI222_X1 U212 ( .A1(n6708), .A2(n670), .B1(n4275), .B2(n3874), .C1(n4164), 
        .C2(n3876), .ZN(n8385) );
  INV_X1 U213 ( .A(n8387), .ZN(n335) );
  INV_X1 U214 ( .A(n335), .ZN(HWDATA[8]) );
  OAI222_X1 U215 ( .A1(n6902), .A2(n670), .B1(n3885), .B2(n3874), .C1(n4006), 
        .C2(n3876), .ZN(n8387) );
  INV_X1 U216 ( .A(n8386), .ZN(n339) );
  INV_X1 U217 ( .A(n339), .ZN(HWDATA[9]) );
  OAI222_X1 U218 ( .A1(n6901), .A2(n670), .B1(n3873), .B2(n3874), .C1(n3337), 
        .C2(n3876), .ZN(n8386) );
  INV_X1 U219 ( .A(n8383), .ZN(n344) );
  INV_X1 U220 ( .A(n344), .ZN(HWDATA[26]) );
  OAI221_X1 U221 ( .B1(n3881), .B2(n3874), .C1(n7653), .C2(n670), .A(n4957), 
        .ZN(n8383) );
  INV_X1 U222 ( .A(n8381), .ZN(n349) );
  INV_X1 U223 ( .A(n349), .ZN(HWDATA[30]) );
  OAI221_X1 U224 ( .B1(n4275), .B2(n3874), .C1(n6897), .C2(n3872), .A(n4887), 
        .ZN(n8381) );
  INV_X1 U225 ( .A(n8382), .ZN(n352) );
  INV_X1 U226 ( .A(n352), .ZN(HWDATA[27]) );
  OAI221_X1 U227 ( .B1(n3773), .B2(n3874), .C1(n6692), .C2(n3872), .A(n4937), 
        .ZN(n8382) );
  INV_X1 U228 ( .A(n8380), .ZN(n356) );
  INV_X1 U229 ( .A(n356), .ZN(HWDATA[31]) );
  OAI221_X1 U230 ( .B1(n4180), .B2(n3874), .C1(n6884), .C2(n3872), .A(n4889), 
        .ZN(n8380) );
  AOI22_X4 U231 ( .A1(n1780), .A2(n941), .B1(n955), .B2(n7422), .ZN(HADDR[7])
         );
  INV_X1 U232 ( .A(n8378), .ZN(n360) );
  INV_X2 U233 ( .A(n360), .ZN(HADDR[2]) );
  AOI22_X1 U234 ( .A1(n1802), .A2(n941), .B1(n3894), .B2(n955), .ZN(n8378) );
  INV_X1 U235 ( .A(n8377), .ZN(n365) );
  AOI22_X1 U236 ( .A1(n1798), .A2(n941), .B1(n3886), .B2(n955), .ZN(n8377) );
  OAI22_X4 U237 ( .A1(n222), .A2(n1610), .B1(n7681), .B2(n950), .ZN(HADDR[23])
         );
  OAI22_X4 U238 ( .A1(n952), .A2(n1633), .B1(n7661), .B2(n946), .ZN(HADDR[20])
         );
  OAI221_X4 U239 ( .B1(n4078), .B2(n3874), .C1(n6727), .C2(n3872), .A(n4877), 
        .ZN(HWDATA[29]) );
  NOR2_X1 U240 ( .A1(n7429), .A2(n950), .ZN(n370) );
  NOR2_X1 U241 ( .A1(n955), .A2(n1606), .ZN(n371) );
  NOR2_X1 U242 ( .A1(n7428), .A2(n946), .ZN(n373) );
  NOR2_X1 U243 ( .A1(n952), .A2(n1639), .ZN(n376) );
  OAI22_X4 U244 ( .A1(n3956), .A2(n3878), .B1(n6887), .B2(n3872), .ZN(
        HWDATA[4]) );
  OAI222_X4 U245 ( .A1(n6906), .A2(n670), .B1(n3885), .B2(n4906), .C1(n4002), 
        .C2(n2692), .ZN(HWDATA[16]) );
  OAI22_X4 U246 ( .A1(n952), .A2(n1616), .B1(n7667), .B2(n950), .ZN(HADDR[22])
         );
  NOR2_X1 U247 ( .A1(n7427), .A2(n946), .ZN(n377) );
  NOR2_X1 U248 ( .A1(n222), .A2(n1652), .ZN(n380) );
  OAI22_X4 U249 ( .A1(n3873), .A2(n3878), .B1(n7491), .B2(n3259), .ZN(
        HWDATA[1]) );
  OAI221_X4 U250 ( .B1(n3885), .B2(n3874), .C1(n6894), .C2(n3872), .A(n4954), 
        .ZN(HWDATA[24]) );
  NOR3_X4 U251 ( .A1(n3411), .A2(n635), .A3(n341), .ZN(n2340) );
  OAI222_X4 U252 ( .A1(n6903), .A2(n670), .B1(n3881), .B2(n4906), .C1(n4379), 
        .C2(n2692), .ZN(HWDATA[18]) );
  OAI22_X4 U253 ( .A1(n222), .A2(n1656), .B1(n7648), .B2(n946), .ZN(HADDR[17])
         );
  OAI221_X4 U254 ( .B1(n1530), .B2(n3887), .C1(n3850), .C2(n950), .A(n3888), 
        .ZN(HTRANS[1]) );
  OAI22_X4 U255 ( .A1(n3773), .A2(n3878), .B1(n6885), .B2(n3872), .ZN(
        HWDATA[3]) );
  NOR3_X4 U256 ( .A1(n3418), .A2(n635), .A3(n331), .ZN(n2331) );
  OAI222_X4 U257 ( .A1(n6718), .A2(n670), .B1(n3956), .B2(n4906), .C1(n4378), 
        .C2(n2692), .ZN(HWDATA[20]) );
  OAI222_X4 U258 ( .A1(n6908), .A2(n670), .B1(n4078), .B2(n3874), .C1(n3040), 
        .C2(n3876), .ZN(HWDATA[13]) );
  OAI22_X4 U259 ( .A1(n955), .A2(n1671), .B1(n7387), .B2(n946), .ZN(HADDR[16])
         );
  OAI22_X4 U260 ( .A1(n7410), .A2(n941), .B1(n955), .B2(n1545), .ZN(HADDR[30])
         );
  OAI22_X4 U261 ( .A1(n2617), .A2(n952), .B1(n911), .B2(n950), .ZN(HWRITE) );
  OAI22_X4 U262 ( .A1(n4078), .A2(n3878), .B1(n6911), .B2(n3872), .ZN(
        HWDATA[5]) );
  NOR3_X4 U263 ( .A1(n3401), .A2(n2150), .A3(n2206), .ZN(n2269) );
  NOR3_X4 U264 ( .A1(n3429), .A2(n635), .A3(n347), .ZN(n2205) );
  OAI222_X4 U265 ( .A1(n6904), .A2(n670), .B1(n3773), .B2(n4906), .C1(n3863), 
        .C2(n2692), .ZN(HWDATA[19]) );
  OAI222_X4 U266 ( .A1(n6875), .A2(n670), .B1(n3956), .B2(n3874), .C1(n4172), 
        .C2(n3876), .ZN(HWDATA[12]) );
  OAI22_X4 U267 ( .A1(n222), .A2(n1693), .B1(n7641), .B2(n946), .ZN(HADDR[14])
         );
  OAI22_X4 U268 ( .A1(n7487), .A2(n941), .B1(n955), .B2(n1529), .ZN(HADDR[31])
         );
  OAI22_X4 U269 ( .A1(n4275), .A2(n3878), .B1(n6900), .B2(n3872), .ZN(
        HWDATA[6]) );
  NOR3_X4 U270 ( .A1(n3426), .A2(n632), .A3(n263), .ZN(n2252) );
  NOR3_X4 U271 ( .A1(n3402), .A2(n2150), .A3(n307), .ZN(n2230) );
  NOR3_X4 U272 ( .A1(n3415), .A2(n635), .A3(n362), .ZN(n2311) );
  OAI22_X4 U273 ( .A1(n952), .A2(n1769), .B1(n7407), .B2(n950), .ZN(HADDR[9])
         );
  OAI222_X4 U274 ( .A1(n6907), .A2(n670), .B1(n4078), .B2(n4906), .C1(n3648), 
        .C2(n2692), .ZN(HWDATA[21]) );
  OAI222_X4 U276 ( .A1(n6756), .A2(n670), .B1(n3773), .B2(n3874), .C1(n2817), 
        .C2(n3876), .ZN(HWDATA[11]) );
  OAI22_X4 U277 ( .A1(n222), .A2(n1709), .B1(n7447), .B2(n946), .ZN(HADDR[13])
         );
  OAI22_X4 U278 ( .A1(n4180), .A2(n3878), .B1(n6889), .B2(n3872), .ZN(
        HWDATA[7]) );
  NOR3_X4 U279 ( .A1(n3427), .A2(n632), .A3(n358), .ZN(n2228) );
  NOR3_X4 U280 ( .A1(n3393), .A2(n2150), .A3(n297), .ZN(n2343) );
  NOR3_X4 U281 ( .A1(n3414), .A2(n635), .A3(n325), .ZN(n2323) );
  OAI22_X4 U282 ( .A1(n952), .A2(n1793), .B1(n7424), .B2(n950), .ZN(HADDR[4])
         );
  OAI222_X4 U283 ( .A1(n6905), .A2(n670), .B1(n3873), .B2(n4906), .C1(n3278), 
        .C2(n2692), .ZN(HWDATA[17]) );
  AOI22_X4 U284 ( .A1(n1774), .A2(n941), .B1(n955), .B2(n7406), .ZN(HADDR[8])
         );
  OAI222_X4 U285 ( .A1(n6750), .A2(n670), .B1(n3881), .B2(n3874), .C1(n3608), 
        .C2(n3876), .ZN(HWDATA[10]) );
  OAI22_X4 U286 ( .A1(n222), .A2(n1718), .B1(n7450), .B2(n946), .ZN(HADDR[12])
         );
  OAI22_X4 U287 ( .A1(n3881), .A2(n3878), .B1(n7491), .B2(n3012), .ZN(
        HWDATA[2]) );
  AOI22_X4 U288 ( .A1(n950), .A2(n1573), .B1(n222), .B2(n7430), .ZN(HADDR[29])
         );
  NOR3_X4 U289 ( .A1(n3403), .A2(n2150), .A3(n312), .ZN(n2314) );
  NOR3_X4 U290 ( .A1(n3430), .A2(n635), .A3(n337), .ZN(n2274) );
  NOR3_X4 U291 ( .A1(n3413), .A2(n632), .A3(n246), .ZN(n2284) );
  OAI222_X4 U292 ( .A1(n6741), .A2(n670), .B1(n4275), .B2(n4906), .C1(n2728), 
        .C2(n2692), .ZN(HWDATA[22]) );
  OAI221_X4 U293 ( .B1(n3873), .B2(n3874), .C1(n6915), .C2(n3872), .A(n4919), 
        .ZN(HWDATA[25]) );
  AOI22_X4 U294 ( .A1(n1738), .A2(n941), .B1(n955), .B2(n7631), .ZN(HADDR[11])
         );
  INV_X1 U295 ( .A(n3141), .ZN(n382) );
  OAI22_X4 U296 ( .A1(n7426), .A2(n3892), .B1(n222), .B2(n2959), .ZN(HADDR[1])
         );
  OAI211_X4 U297 ( .C1(n5245), .C2(n7378), .A(n5246), .B(n5247), .ZN(LOCKUP)
         );
  OAI22_X4 U298 ( .A1(n222), .A2(n1681), .B1(n7437), .B2(n946), .ZN(HADDR[15])
         );
  OAI22_X4 U299 ( .A1(n7306), .A2(n4016), .B1(n7293), .B2(n7315), .ZN(SWDO) );
  NOR2_X4 U300 ( .A1(n2107), .A2(n2121), .ZN(HMASTER) );
  OAI22_X4 U301 ( .A1(n3885), .A2(n3878), .B1(n7491), .B2(n1832), .ZN(
        HWDATA[0]) );
  NOR3_X4 U302 ( .A1(n3417), .A2(n635), .A3(n368), .ZN(n2327) );
  NOR3_X4 U303 ( .A1(n3399), .A2(n2150), .A3(n292), .ZN(n2276) );
  NOR3_X4 U304 ( .A1(n3431), .A2(n632), .A3(n252), .ZN(n2278) );
  NOR3_X4 U305 ( .A1(n3800), .A2(n7374), .A3(n2072), .ZN(TXEV) );
  OAI222_X4 U306 ( .A1(n6912), .A2(n670), .B1(n4180), .B2(n4906), .C1(n3780), 
        .C2(n2692), .ZN(HWDATA[23]) );
  OAI221_X4 U307 ( .B1(n3956), .B2(n3874), .C1(n6882), .C2(n3872), .A(n4849), 
        .ZN(HWDATA[28]) );
  CLKBUF_X1 U308 ( .A(n8379), .Z(HSIZE[0]) );
  NAND2_X1 U309 ( .A1(n3898), .A2(n941), .ZN(n3896) );
  OAI221_X1 U310 ( .B1(n3796), .B2(n3900), .C1(n1801), .C2(n661), .A(n4114), 
        .ZN(\eq_3147/A[1] ) );
  NOR2_X1 U311 ( .A1(n6503), .A2(n3369), .ZN(n5280) );
  NOR2_X1 U312 ( .A1(n3968), .A2(vis_ipsr_o[0]), .ZN(n5798) );
  INV_X1 U313 ( .A(n761), .ZN(n757) );
  INV_X1 U314 ( .A(n768), .ZN(n764) );
  INV_X1 U315 ( .A(n739), .ZN(n737) );
  INV_X1 U316 ( .A(n780), .ZN(n776) );
  INV_X1 U317 ( .A(n686), .ZN(n684) );
  INV_X1 U318 ( .A(n695), .ZN(n691) );
  BUF_X1 U319 ( .A(n210), .Z(n934) );
  INV_X1 U320 ( .A(n234), .ZN(n762) );
  BUF_X1 U321 ( .A(n3851), .Z(n460) );
  INV_X1 U322 ( .A(n4440), .ZN(n2720) );
  INV_X1 U323 ( .A(n499), .ZN(n2603) );
  BUF_X1 U324 ( .A(n678), .Z(n680) );
  BUF_X1 U325 ( .A(n678), .Z(n679) );
  INV_X1 U326 ( .A(n5459), .ZN(n2787) );
  INV_X1 U327 ( .A(n838), .ZN(n2090) );
  NOR2_X1 U328 ( .A1(n3760), .A2(n4193), .ZN(n1661) );
  NOR2_X1 U329 ( .A1(n3068), .A2(n3107), .ZN(n3309) );
  OAI21_X1 U330 ( .B1(n3347), .B2(n3103), .A(n3089), .ZN(n3346) );
  INV_X1 U331 ( .A(n4415), .ZN(n2710) );
  AND2_X1 U332 ( .A1(n2569), .A2(n462), .ZN(n210) );
  INV_X1 U333 ( .A(n5473), .ZN(n3089) );
  NAND3_X1 U334 ( .A1(n5568), .A2(n5569), .A3(n5570), .ZN(n5561) );
  INV_X1 U335 ( .A(n4653), .ZN(n2724) );
  AND2_X1 U336 ( .A1(n5567), .A2(n5600), .ZN(n4343) );
  NAND2_X1 U337 ( .A1(n4343), .A2(n5575), .ZN(n4440) );
  INV_X1 U338 ( .A(n4490), .ZN(n2718) );
  NOR2_X1 U339 ( .A1(n2607), .A2(n4693), .ZN(n499) );
  INV_X1 U340 ( .A(n4148), .ZN(n2717) );
  INV_X1 U341 ( .A(n3565), .ZN(n3851) );
  INV_X1 U342 ( .A(n4347), .ZN(n2716) );
  INV_X1 U343 ( .A(n4150), .ZN(n2721) );
  INV_X1 U344 ( .A(n1628), .ZN(n2547) );
  INV_X1 U345 ( .A(n5567), .ZN(n2725) );
  INV_X1 U346 ( .A(n4173), .ZN(n650) );
  INV_X1 U347 ( .A(n4173), .ZN(n654) );
  INV_X1 U348 ( .A(n1620), .ZN(n4193) );
  NOR3_X1 U349 ( .A1(n516), .A2(n4237), .A3(n4246), .ZN(n3562) );
  INV_X1 U350 ( .A(n5013), .ZN(n3858) );
  NOR2_X1 U351 ( .A1(n3828), .A2(n4237), .ZN(n2880) );
  INV_X1 U352 ( .A(n4094), .ZN(n3805) );
  INV_X1 U353 ( .A(n416), .ZN(n3836) );
  INV_X1 U354 ( .A(Nxkbx6[32]), .ZN(n1544) );
  NAND2_X1 U355 ( .A1(n3749), .A2(n3726), .ZN(n4303) );
  INV_X1 U356 ( .A(n1463), .ZN(n4642) );
  INV_X1 U357 ( .A(n1565), .ZN(n3830) );
  INV_X1 U358 ( .A(n4583), .ZN(n3833) );
  INV_X1 U359 ( .A(n474), .ZN(n4738) );
  INV_X1 U360 ( .A(n1950), .ZN(n4598) );
  INV_X1 U361 ( .A(n3466), .ZN(n4591) );
  INV_X1 U362 ( .A(n3058), .ZN(n2512) );
  INV_X1 U363 ( .A(n511), .ZN(n2575) );
  NAND2_X1 U364 ( .A1(n1986), .A2(n941), .ZN(HPROT_0) );
  INV_X1 U365 ( .A(n222), .ZN(n941) );
  INV_X1 U366 ( .A(n955), .ZN(n946) );
  INV_X1 U367 ( .A(n222), .ZN(n950) );
  AOI22_X1 U368 ( .A1(n4790), .A2(n2782), .B1(n6169), .B2(n2783), .ZN(n6160)
         );
  INV_X1 U369 ( .A(n6170), .ZN(n2782) );
  INV_X1 U370 ( .A(n1763), .ZN(n2607) );
  INV_X1 U371 ( .A(n4790), .ZN(n2783) );
  INV_X1 U372 ( .A(n1902), .ZN(n4608) );
  INV_X1 U373 ( .A(n80), .ZN(n4693) );
  INV_X1 U374 ( .A(n1626), .ZN(n4205) );
  NOR2_X1 U375 ( .A1(n2788), .A2(n3290), .ZN(n5459) );
  INV_X1 U376 ( .A(n5314), .ZN(n3014) );
  NOR2_X1 U377 ( .A1(n2965), .A2(n741), .ZN(n838) );
  INV_X1 U378 ( .A(n5149), .ZN(n2150) );
  INV_X1 U379 ( .A(n1938), .ZN(n4749) );
  OAI21_X1 U380 ( .B1(n2594), .B2(n3836), .A(n4616), .ZN(n462) );
  NOR2_X1 U381 ( .A1(n4738), .A2(n4237), .ZN(n3511) );
  INV_X1 U382 ( .A(n415), .ZN(n3746) );
  INV_X1 U383 ( .A(n3211), .ZN(n3628) );
  INV_X1 U384 ( .A(n808), .ZN(n3766) );
  NOR3_X1 U385 ( .A1(n3831), .A2(n4507), .A3(n4610), .ZN(n4093) );
  INV_X1 U386 ( .A(n1478), .ZN(n3838) );
  INV_X1 U387 ( .A(n4068), .ZN(n2617) );
  INV_X1 U388 ( .A(n483), .ZN(n4756) );
  INV_X1 U389 ( .A(n2116), .ZN(n3855) );
  INV_X1 U390 ( .A(n514), .ZN(n3737) );
  INV_X1 U391 ( .A(n428), .ZN(n4616) );
  INV_X1 U392 ( .A(n2571), .ZN(n4203) );
  INV_X1 U393 ( .A(n1627), .ZN(n3760) );
  INV_X1 U394 ( .A(n275), .ZN(n2513) );
  INV_X1 U395 ( .A(n890), .ZN(n885) );
  NOR2_X1 U396 ( .A1(n1911), .A2(n2594), .ZN(n2894) );
  OAI21_X1 U397 ( .B1(n5677), .B2(n5564), .A(n5568), .ZN(n4415) );
  INV_X1 U398 ( .A(n5391), .ZN(n3108) );
  NOR2_X1 U399 ( .A1(n3081), .A2(n4571), .ZN(n3308) );
  BUF_X1 U400 ( .A(n212), .Z(n931) );
  BUF_X1 U401 ( .A(n3347), .Z(n459) );
  BUF_X1 U402 ( .A(n2569), .Z(n458) );
  NAND2_X1 U403 ( .A1(n3309), .A2(n5564), .ZN(n5568) );
  INV_X1 U404 ( .A(n5661), .ZN(n3080) );
  AOI21_X1 U405 ( .B1(n3832), .B2(n4569), .A(n3308), .ZN(n5661) );
  INV_X1 U406 ( .A(n4565), .ZN(n3068) );
  INV_X1 U407 ( .A(n5657), .ZN(n3078) );
  INV_X1 U408 ( .A(n4571), .ZN(n3832) );
  INV_X1 U409 ( .A(n3353), .ZN(n3107) );
  NAND2_X1 U410 ( .A1(n3091), .A2(n5494), .ZN(n5473) );
  NAND3_X1 U411 ( .A1(n3347), .A2(n3358), .A3(n3108), .ZN(n5494) );
  INV_X1 U412 ( .A(n5274), .ZN(n3103) );
  INV_X1 U413 ( .A(n970), .ZN(n2000) );
  OAI22_X1 U414 ( .A1(n2722), .A2(n3068), .B1(n5677), .B2(n5564), .ZN(n4346)
         );
  OAI21_X1 U415 ( .B1(n2722), .B2(n5657), .A(n5576), .ZN(n4347) );
  NOR2_X1 U416 ( .A1(n5570), .A2(n4571), .ZN(n4653) );
  NOR3_X1 U417 ( .A1(n4205), .A2(n4628), .A3(n3855), .ZN(n3565) );
  INV_X1 U418 ( .A(n734), .ZN(n733) );
  INV_X1 U419 ( .A(n701), .ZN(n696) );
  INV_X1 U420 ( .A(n788), .ZN(n794) );
  INV_X1 U421 ( .A(n788), .ZN(n791) );
  INV_X1 U422 ( .A(n5564), .ZN(n2722) );
  NOR2_X1 U423 ( .A1(n4688), .A2(n2572), .ZN(n1628) );
  NAND2_X1 U424 ( .A1(n5600), .A2(n5601), .ZN(n4150) );
  NOR2_X1 U425 ( .A1(n4738), .A2(n3749), .ZN(n3170) );
  NAND3_X1 U426 ( .A1(n5013), .A2(n1620), .A3(n2722), .ZN(n5575) );
  NAND2_X1 U427 ( .A1(n5576), .A2(n5567), .ZN(n4148) );
  NAND2_X1 U428 ( .A1(n4569), .A2(n5564), .ZN(n5570) );
  NOR2_X1 U429 ( .A1(n2266), .A2(n878), .ZN(n1704) );
  INV_X1 U430 ( .A(n1064), .ZN(n2965) );
  INV_X1 U431 ( .A(n519), .ZN(n3547) );
  NAND2_X1 U432 ( .A1(n514), .A2(n2722), .ZN(n5600) );
  NAND2_X1 U433 ( .A1(n3308), .A2(n5564), .ZN(n5567) );
  INV_X1 U434 ( .A(n2495), .ZN(n2527) );
  INV_X1 U435 ( .A(n1504), .ZN(n3835) );
  OR2_X1 U436 ( .A1(n5601), .A2(n3107), .ZN(n5569) );
  NOR2_X1 U437 ( .A1(n3466), .A2(n3764), .ZN(n3465) );
  NAND2_X1 U438 ( .A1(n5576), .A2(n5569), .ZN(n4490) );
  INV_X1 U439 ( .A(n3165), .ZN(n4222) );
  AND2_X1 U440 ( .A1(n2371), .A2(n2268), .ZN(n2756) );
  INV_X1 U441 ( .A(n496), .ZN(n4602) );
  INV_X1 U442 ( .A(n1624), .ZN(n3761) );
  NOR2_X1 U443 ( .A1(n4631), .A2(n1911), .ZN(n1909) );
  INV_X1 U444 ( .A(n509), .ZN(n4215) );
  INV_X1 U445 ( .A(n2561), .ZN(n1974) );
  INV_X1 U446 ( .A(n692), .ZN(n3762) );
  NOR2_X1 U447 ( .A1(n491), .A2(n477), .ZN(n1902) );
  NOR2_X1 U448 ( .A1(n482), .A2(n267), .ZN(n5013) );
  INV_X1 U449 ( .A(n87), .ZN(n4237) );
  INV_X1 U450 ( .A(n1539), .ZN(n3714) );
  NOR2_X1 U451 ( .A1(n482), .A2(n228), .ZN(n808) );
  INV_X1 U452 ( .A(n1642), .ZN(n3804) );
  INV_X1 U453 ( .A(n3189), .ZN(n3831) );
  NOR2_X1 U454 ( .A1(n254), .A2(n503), .ZN(n1463) );
  NAND2_X1 U455 ( .A1(n493), .A2(n517), .ZN(n3828) );
  INV_X1 U456 ( .A(n1520), .ZN(n3860) );
  INV_X1 U457 ( .A(n693), .ZN(n3749) );
  NOR2_X1 U458 ( .A1(n491), .A2(n267), .ZN(n3466) );
  NOR2_X1 U459 ( .A1(n3831), .A2(n517), .ZN(n1565) );
  NOR2_X1 U460 ( .A1(n4628), .A2(n477), .ZN(n428) );
  INV_X1 U461 ( .A(n493), .ZN(n3764) );
  INV_X1 U462 ( .A(n1663), .ZN(n4229) );
  INV_X1 U463 ( .A(n5253), .ZN(n4628) );
  NOR2_X1 U464 ( .A1(n503), .A2(n482), .ZN(n416) );
  NOR2_X1 U465 ( .A1(n482), .A2(n7355), .ZN(n4583) );
  INV_X1 U466 ( .A(n2743), .ZN(n3730) );
  BUF_X1 U467 ( .A(n5272), .Z(n468) );
  NAND2_X1 U468 ( .A1(n7355), .A2(n272), .ZN(n1528) );
  NOR2_X1 U469 ( .A1(n4193), .A2(n517), .ZN(n3829) );
  NOR2_X1 U470 ( .A1(n3831), .A2(n477), .ZN(n4094) );
  INV_X1 U471 ( .A(n1454), .ZN(n4232) );
  OAI22_X1 U472 ( .A1(n7355), .A2(n3836), .B1(n265), .B2(n3837), .ZN(n5764) );
  INV_X1 U473 ( .A(n4581), .ZN(n4246) );
  INV_X1 U474 ( .A(n52), .ZN(n3837) );
  INV_X1 U475 ( .A(n3561), .ZN(n3800) );
  NAND2_X1 U476 ( .A1(n1748), .A2(n225), .ZN(n3232) );
  INV_X1 U477 ( .A(n63), .ZN(n3788) );
  INV_X1 U478 ( .A(n5775), .ZN(n4650) );
  INV_X1 U479 ( .A(n3509), .ZN(n3732) );
  INV_X1 U480 ( .A(n2742), .ZN(n4202) );
  INV_X1 U481 ( .A(n4298), .ZN(n4631) );
  NAND2_X1 U482 ( .A1(n2743), .A2(n265), .ZN(n5755) );
  INV_X1 U483 ( .A(n1951), .ZN(n3726) );
  INV_X1 U484 ( .A(n4582), .ZN(n4611) );
  INV_X1 U485 ( .A(n4096), .ZN(n4245) );
  INV_X1 U486 ( .A(n5745), .ZN(n4244) );
  INV_X1 U487 ( .A(Nxkbx6[31]), .ZN(n1551) );
  INV_X1 U488 ( .A(n62), .ZN(n3713) );
  INV_X1 U489 ( .A(n2881), .ZN(n2591) );
  INV_X1 U490 ( .A(n1724), .ZN(n4199) );
  INV_X1 U491 ( .A(n5566), .ZN(n4196) );
  INV_X1 U492 ( .A(n230), .ZN(n875) );
  INV_X1 U493 ( .A(n82), .ZN(n2572) );
  INV_X1 U494 ( .A(n230), .ZN(n878) );
  INV_X1 U495 ( .A(n229), .ZN(n640) );
  NOR2_X1 U496 ( .A1(n505), .A2(n875), .ZN(n80) );
  NOR2_X1 U497 ( .A1(n4688), .A2(n7381), .ZN(n1538) );
  INV_X1 U498 ( .A(n1442), .ZN(n4688) );
  NOR2_X1 U499 ( .A1(n4688), .A2(n517), .ZN(n4092) );
  NAND2_X1 U500 ( .A1(n1520), .A2(n493), .ZN(n2873) );
  NOR2_X1 U501 ( .A1(n538), .A2(n482), .ZN(n1504) );
  INV_X1 U502 ( .A(n1462), .ZN(n2594) );
  NOR2_X1 U503 ( .A1(n254), .A2(n482), .ZN(n1478) );
  INV_X1 U504 ( .A(n1457), .ZN(n3623) );
  AOI21_X1 U505 ( .B1(n505), .B2(n513), .A(n1615), .ZN(n3058) );
  NOR2_X1 U506 ( .A1(n521), .A2(n505), .ZN(n4133) );
  NOR2_X1 U507 ( .A1(n503), .A2(n491), .ZN(n1950) );
  NAND2_X1 U508 ( .A1(n3266), .A2(n82), .ZN(n511) );
  NAND3_X1 U509 ( .A1(n1442), .A2(n7381), .A3(n493), .ZN(n3722) );
  INV_X1 U510 ( .A(n1540), .ZN(n4633) );
  INV_X1 U511 ( .A(n1748), .ZN(n4195) );
  INV_X1 U512 ( .A(n1563), .ZN(n4194) );
  AOI21_X1 U513 ( .B1(n230), .B2(n2575), .A(n3134), .ZN(n2611) );
  NOR3_X1 U514 ( .A1(n3858), .A2(n225), .A3(n4598), .ZN(n3134) );
  NAND2_X1 U515 ( .A1(n2743), .A2(n266), .ZN(n4128) );
  INV_X1 U516 ( .A(n2071), .ZN(n3790) );
  INV_X1 U517 ( .A(Nxkbx6[16]), .ZN(n1692) );
  INV_X1 U518 ( .A(Nxkbx6[24]), .ZN(n1614) );
  OAI22_X1 U519 ( .A1(n5316), .A2(n6172), .B1(n6173), .B2(n6174), .ZN(n4790)
         );
  OAI22_X1 U520 ( .A1(n5309), .A2(n6171), .B1(n6169), .B2(n6170), .ZN(n6174)
         );
  AOI22_X1 U521 ( .A1(n2786), .A2(n6166), .B1(n6169), .B2(n6170), .ZN(n6173)
         );
  INV_X1 U522 ( .A(n6165), .ZN(n2786) );
  NOR2_X1 U523 ( .A1(n2608), .A2(n517), .ZN(n1763) );
  NOR2_X1 U524 ( .A1(n4608), .A2(n517), .ZN(n496) );
  NOR2_X1 U525 ( .A1(n4229), .A2(n517), .ZN(n1626) );
  OAI22_X1 U526 ( .A1(n5309), .A2(n2790), .B1(n3287), .B2(n2788), .ZN(n6170)
         );
  AND2_X1 U527 ( .A1(n5602), .A2(n5656), .ZN(n4349) );
  OAI21_X1 U528 ( .B1(n3078), .B2(n4565), .A(n5564), .ZN(n5656) );
  INV_X1 U529 ( .A(n6193), .ZN(n3290) );
  NOR2_X1 U530 ( .A1(n3015), .A2(n3016), .ZN(n5314) );
  BUF_X1 U531 ( .A(n3901), .Z(n661) );
  NAND3_X1 U532 ( .A1(n267), .A2(n1620), .A3(n1567), .ZN(n3729) );
  INV_X1 U533 ( .A(n131), .ZN(n1537) );
  AOI22_X1 U534 ( .A1(n6165), .A2(n4790), .B1(n6166), .B2(n2783), .ZN(n6157)
         );
  BUF_X1 U535 ( .A(n3900), .Z(n664) );
  NAND2_X1 U536 ( .A1(n1455), .A2(n1442), .ZN(n3221) );
  AOI21_X1 U537 ( .B1(n254), .B2(n693), .A(n2903), .ZN(n4073) );
  INV_X1 U538 ( .A(n72), .ZN(n2529) );
  INV_X1 U539 ( .A(n5309), .ZN(n2788) );
  INV_X1 U540 ( .A(n5316), .ZN(n3015) );
  NAND3_X1 U541 ( .A1(n5253), .A2(n1457), .A3(n1748), .ZN(n1524) );
  INV_X1 U542 ( .A(n1567), .ZN(n2608) );
  INV_X1 U543 ( .A(n1952), .ZN(n2528) );
  BUF_X1 U544 ( .A(n955), .Z(n952) );
  INV_X1 U545 ( .A(n6198), .ZN(n3287) );
  INV_X1 U546 ( .A(n407), .ZN(n1805) );
  INV_X1 U547 ( .A(n3891), .ZN(n2121) );
  INV_X1 U548 ( .A(n3660), .ZN(n3954) );
  BUF_X1 U549 ( .A(n222), .Z(n955) );
  INV_X1 U550 ( .A(n1532), .ZN(n2516) );
  INV_X1 U551 ( .A(Nxkbx6[6]), .ZN(n1790) );
  INV_X1 U552 ( .A(n1124), .ZN(n2086) );
  INV_X1 U553 ( .A(n1125), .ZN(n2092) );
  AOI21_X1 U554 ( .B1(n210), .B2(n2150), .A(n213), .ZN(n273) );
  INV_X1 U555 ( .A(n884), .ZN(n2082) );
  AOI211_X1 U556 ( .C1(n7375), .C2(n1748), .A(n4583), .B(n63), .ZN(n3897) );
  NOR2_X1 U557 ( .A1(n2608), .A2(n503), .ZN(n1761) );
  NOR2_X1 U558 ( .A1(n878), .A2(n7381), .ZN(n3211) );
  NOR2_X1 U559 ( .A1(n477), .A2(n521), .ZN(n1624) );
  NOR2_X1 U560 ( .A1(n477), .A2(n517), .ZN(n1938) );
  NOR2_X1 U561 ( .A1(n3749), .A2(n267), .ZN(n514) );
  INV_X1 U562 ( .A(n2915), .ZN(n4610) );
  NOR2_X1 U563 ( .A1(n3749), .A2(n477), .ZN(n415) );
  NOR3_X1 U564 ( .A1(n2783), .A2(n5309), .A3(n6171), .ZN(n6161) );
  AOI22_X1 U565 ( .A1(n3048), .A2(n3015), .B1(n6179), .B2(n5316), .ZN(n6169)
         );
  INV_X1 U566 ( .A(n6180), .ZN(n3048) );
  NOR2_X1 U567 ( .A1(n477), .A2(n505), .ZN(n483) );
  OAI211_X1 U568 ( .C1(n4088), .C2(n4591), .A(n4089), .B(n4090), .ZN(n4068) );
  AOI22_X1 U569 ( .A1(n4095), .A2(n265), .B1(n4096), .B2(n230), .ZN(n4088) );
  OAI21_X1 U570 ( .B1(n4093), .B2(n4094), .A(n693), .ZN(n4089) );
  AOI211_X1 U571 ( .C1(n4091), .C2(n4092), .A(n483), .B(n1649), .ZN(n4090) );
  INV_X1 U572 ( .A(n37), .ZN(n2524) );
  NOR2_X1 U573 ( .A1(n491), .A2(n521), .ZN(n2563) );
  NOR2_X1 U574 ( .A1(n4749), .A2(n521), .ZN(n1627) );
  NOR2_X1 U575 ( .A1(n4229), .A2(n491), .ZN(n2571) );
  NAND2_X1 U576 ( .A1(n2163), .A2(n796), .ZN(n746) );
  NAND2_X1 U577 ( .A1(n3897), .A2(n2693), .ZN(n2439) );
  INV_X1 U578 ( .A(n433), .ZN(n4507) );
  NOR3_X1 U579 ( .A1(n3855), .A2(n1994), .A3(n3746), .ZN(n4079) );
  INV_X1 U581 ( .A(n1584), .ZN(n2698) );
  NOR2_X1 U582 ( .A1(n878), .A2(n482), .ZN(n2116) );
  NOR2_X1 U583 ( .A1(n4203), .A2(n3173), .ZN(n1649) );
  INV_X1 U584 ( .A(n202), .ZN(n1986) );
  INV_X1 U585 ( .A(n1751), .ZN(n2275) );
  INV_X1 U586 ( .A(n429), .ZN(n3709) );
  NAND3_X1 U587 ( .A1(n5601), .A2(n5568), .A3(n5602), .ZN(n5149) );
  INV_X1 U588 ( .A(n877), .ZN(n2096) );
  INV_X1 U589 ( .A(n1674), .ZN(n1926) );
  INV_X1 U590 ( .A(n4084), .ZN(n3787) );
  NAND2_X1 U591 ( .A1(n491), .A2(n3838), .ZN(n5240) );
  OAI21_X1 U592 ( .B1(n4507), .B2(n3173), .A(n4097), .ZN(n4095) );
  NAND3_X1 U593 ( .A1(n230), .A2(n516), .A3(n524), .ZN(n4097) );
  NAND4_X1 U594 ( .A1(n1718), .A2(n1671), .A3(n1656), .A4(n1652), .ZN(n140) );
  INV_X1 U595 ( .A(n1908), .ZN(n4732) );
  INV_X1 U596 ( .A(n752), .ZN(n2189) );
  INV_X1 U597 ( .A(n4789), .ZN(n2212) );
  INV_X1 U598 ( .A(n6199), .ZN(n2790) );
  NAND2_X1 U599 ( .A1(n3788), .A2(n84), .ZN(n4082) );
  NOR3_X1 U600 ( .A1(n3110), .A2(n3305), .A3(n3111), .ZN(n4565) );
  INV_X1 U601 ( .A(n233), .ZN(n906) );
  INV_X1 U602 ( .A(n631), .ZN(n629) );
  INV_X1 U603 ( .A(n239), .ZN(n881) );
  INV_X1 U604 ( .A(n399), .ZN(n784) );
  INV_X1 U605 ( .A(n399), .ZN(n783) );
  NAND2_X1 U606 ( .A1(n3475), .A2(n883), .ZN(n735) );
  NAND2_X1 U607 ( .A1(n3475), .A2(n883), .ZN(n456) );
  AOI221_X1 U608 ( .B1(n2420), .B2(n3308), .C1(n3349), .C2(n4565), .A(n2361), 
        .ZN(n3459) );
  INV_X1 U609 ( .A(n3315), .ZN(n2420) );
  INV_X1 U610 ( .A(n4567), .ZN(n2361) );
  AOI221_X1 U611 ( .B1(n3078), .B2(n2364), .C1(n4568), .C2(n4569), .A(n4570), 
        .ZN(n4567) );
  INV_X1 U612 ( .A(n1080), .ZN(n2094) );
  NAND3_X1 U613 ( .A1(n693), .A2(n906), .A3(n677), .ZN(n675) );
  NOR2_X1 U614 ( .A1(n461), .A2(n3058), .ZN(n275) );
  INV_X1 U615 ( .A(n241), .ZN(n1849) );
  NOR3_X1 U616 ( .A1(n2512), .A2(n461), .A3(n462), .ZN(n212) );
  NOR2_X1 U617 ( .A1(n521), .A2(n5274), .ZN(n4762) );
  NOR2_X1 U618 ( .A1(n516), .A2(n3189), .ZN(n4571) );
  NOR2_X1 U619 ( .A1(n4550), .A2(n3305), .ZN(n4569) );
  INV_X1 U620 ( .A(n4690), .ZN(n3104) );
  INV_X1 U621 ( .A(n6041), .ZN(n3111) );
  NOR2_X1 U622 ( .A1(n3108), .A2(n3105), .ZN(n5274) );
  INV_X1 U623 ( .A(n182), .ZN(n1847) );
  INV_X1 U624 ( .A(n2496), .ZN(n4685) );
  NAND2_X1 U625 ( .A1(n3108), .A2(n3105), .ZN(n5675) );
  OAI21_X1 U626 ( .B1(n5274), .B2(n5275), .A(n5276), .ZN(n5271) );
  NAND3_X1 U627 ( .A1(n459), .A2(n631), .A3(n3089), .ZN(n5276) );
  AOI21_X1 U628 ( .B1(n3091), .B2(n629), .A(n3089), .ZN(n5275) );
  NAND2_X1 U629 ( .A1(n1454), .A2(n7375), .ZN(n1911) );
  NOR2_X1 U630 ( .A1(n6536), .A2(n6533), .ZN(n6527) );
  NOR2_X1 U631 ( .A1(n2001), .A2(n2002), .ZN(n970) );
  NAND2_X1 U632 ( .A1(n732), .A2(n840), .ZN(n858) );
  NAND2_X1 U633 ( .A1(n3354), .A2(n3832), .ZN(n5657) );
  INV_X1 U634 ( .A(n1643), .ZN(n4818) );
  AOI22_X1 U635 ( .A1(n4543), .A2(n4544), .B1(n3111), .B2(n3315), .ZN(n4542)
         );
  OAI21_X1 U636 ( .B1(n2364), .B2(n3111), .A(n3110), .ZN(n4543) );
  OR3_X1 U637 ( .A1(n3111), .A2(n3110), .A3(n4547), .ZN(n4544) );
  NAND3_X1 U638 ( .A1(n412), .A2(n1452), .A3(N701), .ZN(n2904) );
  NAND3_X1 U639 ( .A1(n3108), .A2(n4734), .A3(n4762), .ZN(n4736) );
  INV_X1 U640 ( .A(n2408), .ZN(n1927) );
  NOR2_X1 U641 ( .A1(n4549), .A2(n4550), .ZN(n4541) );
  NAND2_X1 U642 ( .A1(n516), .A2(n6033), .ZN(n3353) );
  INV_X1 U643 ( .A(n4458), .ZN(n3763) );
  NOR2_X1 U644 ( .A1(n3056), .A2(n5316), .ZN(n5320) );
  INV_X1 U645 ( .A(n3374), .ZN(n2364) );
  INV_X1 U646 ( .A(n4549), .ZN(n2391) );
  NAND2_X1 U647 ( .A1(n3832), .A2(n6033), .ZN(n5391) );
  NOR2_X1 U648 ( .A1(n4571), .A2(n4549), .ZN(n4568) );
  INV_X1 U649 ( .A(n513), .ZN(n2509) );
  INV_X1 U650 ( .A(n461), .ZN(n2569) );
  INV_X1 U651 ( .A(n409), .ZN(n1979) );
  NOR2_X1 U652 ( .A1(n5253), .A2(n87), .ZN(n6544) );
  INV_X1 U653 ( .A(n4734), .ZN(n3347) );
  INV_X1 U654 ( .A(n1166), .ZN(n2004) );
  INV_X1 U655 ( .A(n5987), .ZN(n3081) );
  NAND2_X1 U656 ( .A1(n5172), .A2(n4609), .ZN(n2237) );
  NAND2_X1 U657 ( .A1(n5172), .A2(n4748), .ZN(n2289) );
  AND2_X1 U658 ( .A1(n2710), .A2(n6424), .ZN(n5572) );
  NAND3_X1 U659 ( .A1(n2722), .A2(n538), .A3(n4133), .ZN(n6424) );
  INV_X1 U660 ( .A(n3294), .ZN(n2609) );
  INV_X1 U661 ( .A(n840), .ZN(n2001) );
  INV_X1 U662 ( .A(n5495), .ZN(n3091) );
  INV_X1 U663 ( .A(n4733), .ZN(n3102) );
  OAI21_X1 U664 ( .B1(n4734), .B2(n4735), .A(n4736), .ZN(n4733) );
  INV_X1 U665 ( .A(n1747), .ZN(n2506) );
  INV_X1 U666 ( .A(n4758), .ZN(n3101) );
  OAI211_X1 U667 ( .C1(n4735), .C2(n4759), .A(n4760), .B(n4736), .ZN(n4758) );
  NAND2_X1 U668 ( .A1(n459), .A2(n631), .ZN(n4759) );
  NAND3_X1 U669 ( .A1(n3108), .A2(n629), .A3(n4762), .ZN(n4760) );
  INV_X1 U670 ( .A(n3920), .ZN(n1812) );
  NAND2_X1 U671 ( .A1(n1166), .A2(n732), .ZN(n1165) );
  INV_X1 U672 ( .A(n5988), .ZN(n3072) );
  OAI21_X1 U673 ( .B1(n4569), .B2(n3354), .A(n3353), .ZN(n5988) );
  NAND2_X1 U674 ( .A1(n840), .A2(n2096), .ZN(n1120) );
  NAND2_X1 U675 ( .A1(n4609), .A2(n4401), .ZN(n2285) );
  INV_X1 U676 ( .A(n2902), .ZN(n2125) );
  AOI211_X1 U677 ( .C1(n429), .C2(n1563), .A(n2903), .B(n2904), .ZN(n2902) );
  INV_X1 U678 ( .A(n5318), .ZN(n3060) );
  INV_X1 U679 ( .A(n183), .ZN(n2133) );
  OAI221_X1 U680 ( .B1(n3232), .B2(n3855), .C1(n2529), .C2(n4610), .A(n3222), 
        .ZN(n2495) );
  NOR2_X1 U681 ( .A1(n3749), .A2(n3765), .ZN(n99) );
  INV_X1 U682 ( .A(n233), .ZN(n897) );
  NOR2_X1 U683 ( .A1(n914), .A2(n1342), .ZN(n1064) );
  INV_X1 U684 ( .A(n226), .ZN(n672) );
  INV_X1 U685 ( .A(n4717), .ZN(n3106) );
  NOR2_X1 U686 ( .A1(n3548), .A2(n7381), .ZN(n519) );
  NAND2_X1 U687 ( .A1(n4250), .A2(n6453), .ZN(n5564) );
  NAND3_X1 U688 ( .A1(n4507), .A2(n2726), .A3(n477), .ZN(n6453) );
  NAND3_X1 U689 ( .A1(n1520), .A2(n516), .A3(n1950), .ZN(n504) );
  OAI221_X1 U690 ( .B1(n4651), .B2(n2071), .C1(n272), .C2(n2072), .A(n2067), 
        .ZN(n1957) );
  AOI21_X1 U691 ( .B1(n2529), .B2(n237), .A(n4298), .ZN(n1924) );
  NAND2_X1 U692 ( .A1(n2722), .A2(n493), .ZN(n5576) );
  NAND2_X1 U693 ( .A1(n270), .A2(n7514), .ZN(n93) );
  NOR2_X1 U694 ( .A1(n4229), .A2(n267), .ZN(n3165) );
  NOR2_X1 U695 ( .A1(n4738), .A2(n521), .ZN(n497) );
  NOR2_X1 U696 ( .A1(n2243), .A2(n270), .ZN(n2916) );
  NAND2_X1 U697 ( .A1(n90), .A2(n7514), .ZN(n2371) );
  NAND2_X1 U698 ( .A1(n267), .A2(n493), .ZN(n2755) );
  NAND2_X1 U699 ( .A1(n1563), .A2(n272), .ZN(n412) );
  NOR3_X1 U700 ( .A1(n3749), .A2(n524), .A3(n266), .ZN(n5565) );
  BUF_X1 U701 ( .A(n537), .Z(n928) );
  AOI21_X1 U702 ( .B1(n4628), .B2(n4611), .A(n524), .ZN(n5677) );
  BUF_X1 U703 ( .A(n3582), .Z(n674) );
  NAND2_X1 U704 ( .A1(n1908), .A2(n90), .ZN(n2377) );
  OAI21_X1 U705 ( .B1(n5037), .B2(n1923), .A(n3122), .ZN(n3270) );
  INV_X1 U706 ( .A(n90), .ZN(n2273) );
  NAND2_X1 U707 ( .A1(n228), .A2(n265), .ZN(n692) );
  NAND2_X1 U708 ( .A1(n3141), .A2(n913), .ZN(n551) );
  NAND2_X1 U709 ( .A1(n3354), .A2(n5564), .ZN(n5601) );
  AOI22_X1 U710 ( .A1(n63), .A2(n37), .B1(n1951), .B2(n1952), .ZN(n1940) );
  NOR2_X1 U711 ( .A1(n460), .A2(n2357), .ZN(n2354) );
  NOR2_X1 U712 ( .A1(n460), .A2(n3660), .ZN(n2602) );
  AOI21_X1 U713 ( .B1(n4245), .B2(n3173), .A(n2529), .ZN(n3172) );
  NAND2_X1 U714 ( .A1(n3565), .A2(n3983), .ZN(n2831) );
  INV_X1 U715 ( .A(n417), .ZN(n2726) );
  NAND2_X1 U716 ( .A1(n3511), .A2(n429), .ZN(n3568) );
  NAND2_X1 U717 ( .A1(n4222), .A2(n447), .ZN(n509) );
  INV_X1 U718 ( .A(n2899), .ZN(n3122) );
  NOR2_X1 U719 ( .A1(n482), .A2(n1975), .ZN(n1562) );
  INV_X1 U720 ( .A(n2073), .ZN(n2519) );
  INV_X1 U721 ( .A(n88), .ZN(n1958) );
  INV_X1 U722 ( .A(n2560), .ZN(n4651) );
  NAND2_X1 U723 ( .A1(n3097), .A2(n2273), .ZN(n1697) );
  INV_X1 U724 ( .A(n1511), .ZN(n2697) );
  INV_X1 U725 ( .A(n1488), .ZN(n1925) );
  NAND2_X1 U726 ( .A1(n3266), .A2(n225), .ZN(n2911) );
  INV_X1 U727 ( .A(n1918), .ZN(n2268) );
  INV_X1 U728 ( .A(n1342), .ZN(n2964) );
  INV_X1 U729 ( .A(n4254), .ZN(n2550) );
  INV_X1 U730 ( .A(n2488), .ZN(n2254) );
  OR4_X1 U731 ( .A1(n2072), .A2(n3860), .A3(n272), .A4(n875), .ZN(n3715) );
  INV_X1 U732 ( .A(n5220), .ZN(n4190) );
  INV_X1 U733 ( .A(n4317), .ZN(n1923) );
  INV_X1 U734 ( .A(n2941), .ZN(n2610) );
  INV_X1 U735 ( .A(n4256), .ZN(n2549) );
  INV_X1 U736 ( .A(n2067), .ZN(n3786) );
  INV_X1 U737 ( .A(n3181), .ZN(n4566) );
  NAND2_X1 U738 ( .A1(n674), .A2(n3258), .ZN(n3671) );
  INV_X1 U739 ( .A(n6534), .ZN(n2714) );
  INV_X1 U740 ( .A(n5776), .ZN(n4250) );
  NAND2_X1 U741 ( .A1(n3582), .A2(n2477), .ZN(n3619) );
  INV_X1 U742 ( .A(n1588), .ZN(n2266) );
  INV_X1 U743 ( .A(n4231), .ZN(n3727) );
  OR2_X1 U744 ( .A1(n3851), .A2(n457), .ZN(n698) );
  INV_X1 U745 ( .A(n3001), .ZN(n3697) );
  INV_X1 U746 ( .A(n2492), .ZN(n2247) );
  INV_X1 U747 ( .A(n5574), .ZN(n3768) );
  INV_X1 U748 ( .A(n98), .ZN(n2508) );
  INV_X1 U749 ( .A(n28), .ZN(n1936) );
  INV_X1 U750 ( .A(n2306), .ZN(n3843) );
  INV_X1 U751 ( .A(n2103), .ZN(n800) );
  INV_X1 U752 ( .A(n389), .ZN(n892) );
  INV_X1 U753 ( .A(n389), .ZN(n894) );
  NOR3_X1 U754 ( .A1(n1563), .A2(n1462), .A3(n509), .ZN(n2414) );
  NAND3_X1 U755 ( .A1(n3221), .A2(n4651), .A3(n3222), .ZN(n1705) );
  OAI21_X1 U756 ( .B1(n474), .B2(n415), .A(n7375), .ZN(n2567) );
  OAI21_X1 U757 ( .B1(n237), .B2(n3788), .A(n4685), .ZN(n1699) );
  NAND4_X1 U758 ( .A1(n3189), .A2(n7355), .A3(n1455), .A4(n230), .ZN(n3182) );
  INV_X1 U759 ( .A(n1455), .ZN(n2515) );
  NAND3_X1 U760 ( .A1(n7355), .A2(n1620), .A3(n875), .ZN(n3220) );
  NOR2_X1 U761 ( .A1(n1975), .A2(n878), .ZN(n2561) );
  NOR2_X1 U762 ( .A1(n482), .A2(n4195), .ZN(n1621) );
  INV_X1 U763 ( .A(n1505), .ZN(n3705) );
  INV_X1 U764 ( .A(n1760), .ZN(n4564) );
  INV_X1 U765 ( .A(n2767), .ZN(n2614) );
  INV_X1 U766 ( .A(n1586), .ZN(n2246) );
  NOR2_X1 U767 ( .A1(n508), .A2(n7375), .ZN(n1520) );
  NOR2_X1 U768 ( .A1(n4263), .A2(n485), .ZN(n1642) );
  NOR2_X1 U769 ( .A1(n523), .A2(n482), .ZN(n1539) );
  NOR2_X1 U770 ( .A1(n522), .A2(n538), .ZN(n693) );
  NOR2_X1 U771 ( .A1(n529), .A2(n521), .ZN(n82) );
  INV_X1 U772 ( .A(n4259), .ZN(n2730) );
  NOR2_X1 U773 ( .A1(n477), .A2(n7282), .ZN(n1663) );
  NOR2_X2 U774 ( .A1(n526), .A2(n7374), .ZN(n1462) );
  NOR2_X1 U775 ( .A1(n508), .A2(n536), .ZN(n1454) );
  NOR2_X1 U776 ( .A1(n485), .A2(n7373), .ZN(n3189) );
  INV_X1 U777 ( .A(n486), .ZN(n482) );
  INV_X1 U778 ( .A(n7374), .ZN(n491) );
  INV_X1 U779 ( .A(n7282), .ZN(n538) );
  INV_X1 U780 ( .A(n502), .ZN(n503) );
  INV_X1 U781 ( .A(n523), .ZN(n521) );
  INV_X1 U782 ( .A(n508), .ZN(n505) );
  INV_X1 U783 ( .A(n479), .ZN(n477) );
  NOR2_X1 U784 ( .A1(n254), .A2(n536), .ZN(n1748) );
  NOR2_X1 U785 ( .A1(n522), .A2(n267), .ZN(n2743) );
  NOR2_X1 U786 ( .A1(n463), .A2(n482), .ZN(n52) );
  NOR2_X1 U787 ( .A1(n479), .A2(n7374), .ZN(n4298) );
  NOR2_X1 U788 ( .A1(n503), .A2(n7374), .ZN(n5253) );
  AOI222_X1 U789 ( .A1(n529), .A2(n4096), .B1(n5013), .B2(n4581), .C1(n5253), 
        .C2(n1663), .ZN(n4127) );
  NOR2_X1 U790 ( .A1(n503), .A2(n485), .ZN(n63) );
  NOR2_X1 U791 ( .A1(n463), .A2(n7373), .ZN(n4581) );
  NOR2_X1 U792 ( .A1(n491), .A2(n7282), .ZN(n87) );
  NOR2_X1 U793 ( .A1(n485), .A2(n505), .ZN(n3561) );
  NOR2_X1 U794 ( .A1(n3860), .A2(n522), .ZN(n1951) );
  NOR2_X1 U795 ( .A1(n503), .A2(n536), .ZN(n2742) );
  BUF_X1 U796 ( .A(n4868), .Z(n581) );
  NAND2_X1 U797 ( .A1(n1539), .A2(n4263), .ZN(n3173) );
  BUF_X1 U798 ( .A(n4856), .Z(n628) );
  BUF_X1 U799 ( .A(n4860), .Z(n623) );
  BUF_X1 U800 ( .A(n5999), .Z(n565) );
  BUF_X1 U801 ( .A(n6004), .Z(n550) );
  NOR2_X1 U802 ( .A1(n4265), .A2(n7282), .ZN(n1724) );
  NOR2_X1 U803 ( .A1(n492), .A2(n505), .ZN(n4582) );
  NOR2_X1 U804 ( .A1(n503), .A2(n463), .ZN(n4096) );
  NOR2_X1 U805 ( .A1(n502), .A2(n505), .ZN(n5775) );
  BUF_X1 U806 ( .A(n4176), .Z(n646) );
  NOR2_X1 U807 ( .A1(n508), .A2(n522), .ZN(n3509) );
  BUF_X1 U808 ( .A(n3789), .Z(n671) );
  BUF_X1 U809 ( .A(n4864), .Z(n599) );
  BUF_X1 U810 ( .A(n4862), .Z(n615) );
  BUF_X1 U811 ( .A(n4858), .Z(n627) );
  BUF_X1 U812 ( .A(n4872), .Z(n576) );
  BUF_X1 U813 ( .A(n4867), .Z(n582) );
  BUF_X1 U814 ( .A(n4875), .Z(n572) );
  INV_X1 U815 ( .A(\eq_3147/A[26] ), .ZN(n1580) );
  NOR2_X1 U816 ( .A1(n3714), .A2(n7373), .ZN(n62) );
  INV_X1 U817 ( .A(n201), .ZN(n1573) );
  NOR3_X1 U818 ( .A1(n522), .A2(n5253), .A3(n63), .ZN(n5750) );
  NOR2_X1 U819 ( .A1(n3858), .A2(n526), .ZN(n2881) );
  NOR2_X1 U820 ( .A1(n4650), .A2(n536), .ZN(n5566) );
  NOR2_X1 U821 ( .A1(n463), .A2(n492), .ZN(n5745) );
  INV_X1 U822 ( .A(\eq_3147/A[25] ), .ZN(n1582) );
  INV_X1 U823 ( .A(n200), .ZN(n1545) );
  AOI21_X1 U824 ( .B1(n5760), .B2(n808), .A(n5745), .ZN(n5759) );
  NOR2_X1 U825 ( .A1(n4202), .A2(n4265), .ZN(n5760) );
  NAND2_X1 U826 ( .A1(n267), .A2(n7373), .ZN(n2754) );
  NAND2_X1 U827 ( .A1(n492), .A2(n485), .ZN(n2071) );
  INV_X1 U828 ( .A(n4288), .ZN(n2473) );
  NOR2_X1 U829 ( .A1(n671), .A2(n2334), .ZN(Idfpw6[25]) );
  NOR2_X1 U830 ( .A1(n671), .A2(n2328), .ZN(Idfpw6[26]) );
  NOR2_X1 U831 ( .A1(n671), .A2(n2324), .ZN(Idfpw6[27]) );
  INV_X1 U832 ( .A(n4503), .ZN(n2338) );
  INV_X1 U833 ( .A(n5018), .ZN(n5272) );
  BUF_X1 U834 ( .A(n4173), .Z(n660) );
  BUF_X1 U835 ( .A(n7355), .Z(n517) );
  NOR2_X1 U836 ( .A1(n4512), .A2(n524), .ZN(n417) );
  INV_X1 U837 ( .A(n4258), .ZN(n2545) );
  NOR2_X1 U838 ( .A1(n476), .A2(n875), .ZN(n1457) );
  NOR2_X1 U839 ( .A1(n4738), .A2(n536), .ZN(n1563) );
  NOR2_X1 U840 ( .A1(n508), .A2(n491), .ZN(n2915) );
  NOR2_X1 U841 ( .A1(n479), .A2(n875), .ZN(n1442) );
  NOR2_X1 U842 ( .A1(n529), .A2(n7373), .ZN(n513) );
  NOR3_X1 U843 ( .A1(n2572), .A2(n485), .A3(n479), .ZN(n5219) );
  INV_X1 U844 ( .A(n526), .ZN(n524) );
  NOR2_X1 U845 ( .A1(n4512), .A2(n875), .ZN(n433) );
  AOI21_X1 U846 ( .B1(n505), .B2(n7375), .A(n2915), .ZN(n5211) );
  INV_X1 U847 ( .A(n4092), .ZN(n4687) );
  NOR2_X1 U848 ( .A1(n523), .A2(n485), .ZN(n429) );
  NOR2_X1 U849 ( .A1(n2594), .A2(n7373), .ZN(n1615) );
  NOR2_X1 U850 ( .A1(n477), .A2(n492), .ZN(n1540) );
  NOR2_X1 U851 ( .A1(n508), .A2(n538), .ZN(n5220) );
  NOR3_X1 U852 ( .A1(n4202), .A2(n7375), .A3(n4265), .ZN(n3266) );
  NOR2_X1 U853 ( .A1(n3285), .A2(n354), .ZN(n4354) );
  BUF_X1 U854 ( .A(n4861), .Z(n617) );
  BUF_X1 U855 ( .A(n6004), .Z(n547) );
  BUF_X1 U856 ( .A(n4863), .Z(n602) );
  NOR3_X1 U857 ( .A1(n3623), .A2(n228), .A3(n4243), .ZN(n5217) );
  INV_X1 U858 ( .A(\eq_3147/A[22] ), .ZN(n1606) );
  NOR3_X1 U859 ( .A1(n3837), .A2(n517), .A3(n479), .ZN(n5207) );
  NAND2_X1 U860 ( .A1(n492), .A2(n516), .ZN(n84) );
  INV_X1 U861 ( .A(\eq_3147/A[16] ), .ZN(n1652) );
  NAND4_X1 U862 ( .A1(n1565), .A2(n87), .A3(n508), .A4(n4263), .ZN(n4130) );
  INV_X1 U863 ( .A(\eq_3147/A[15] ), .ZN(n1656) );
  INV_X1 U864 ( .A(\eq_3147/A[14] ), .ZN(n1671) );
  INV_X1 U865 ( .A(\eq_3147/A[23] ), .ZN(n1603) );
  INV_X1 U866 ( .A(\eq_3147/A[21] ), .ZN(n1610) );
  INV_X1 U867 ( .A(\eq_3147/A[17] ), .ZN(n1639) );
  INV_X1 U868 ( .A(\eq_3147/A[18] ), .ZN(n1633) );
  INV_X1 U869 ( .A(\eq_3147/A[24] ), .ZN(n1596) );
  INV_X1 U870 ( .A(\eq_3147/A[19] ), .ZN(n1631) );
  INV_X1 U871 ( .A(\eq_3147/A[20] ), .ZN(n1616) );
  NAND4_X1 U872 ( .A1(n1680), .A2(n1669), .A3(n3390), .A4(n3391), .ZN(n3387)
         );
  INV_X1 U873 ( .A(n3403), .ZN(n1680) );
  INV_X1 U874 ( .A(n3402), .ZN(n1669) );
  NOR3_X1 U875 ( .A1(n3399), .A2(n3400), .A3(n3401), .ZN(n3390) );
  NAND4_X1 U876 ( .A1(n1716), .A2(n1782), .A3(n3406), .A4(n3407), .ZN(n3386)
         );
  INV_X1 U877 ( .A(n3417), .ZN(n1782) );
  INV_X1 U878 ( .A(n3418), .ZN(n1716) );
  NOR3_X1 U879 ( .A1(n3414), .A2(n3415), .A3(n3416), .ZN(n3406) );
  INV_X1 U880 ( .A(\eq_3147/A[13] ), .ZN(n1681) );
  AOI21_X1 U882 ( .B1(n1464), .B2(n3548), .A(n4688), .ZN(n5218) );
  NAND2_X1 U883 ( .A1(n2512), .A2(n3059), .ZN(n3285) );
  INV_X1 U884 ( .A(n4290), .ZN(n2468) );
  INV_X1 U885 ( .A(n4291), .ZN(n2322) );
  INV_X1 U886 ( .A(n2376), .ZN(n3548) );
  INV_X1 U887 ( .A(n5251), .ZN(n4271) );
  NOR2_X1 U888 ( .A1(n680), .A2(n2459), .ZN(Mifpw6[0]) );
  NOR2_X1 U889 ( .A1(n679), .A2(n5278), .ZN(Tgfpw6[6]) );
  NOR2_X1 U890 ( .A1(n679), .A2(n5277), .ZN(Tgfpw6[5]) );
  NOR2_X1 U891 ( .A1(n2611), .A2(n5282), .ZN(Tgfpw6[4]) );
  NOR2_X1 U892 ( .A1(n2611), .A2(n4351), .ZN(Tgfpw6[1]) );
  NOR2_X1 U893 ( .A1(n680), .A2(n2458), .ZN(Mifpw6[1]) );
  NOR2_X1 U894 ( .A1(n679), .A2(n2460), .ZN(Mifpw6[3]) );
  NOR2_X1 U895 ( .A1(n679), .A2(n2355), .ZN(Mifpw6[4]) );
  NOR2_X1 U896 ( .A1(n679), .A2(n2347), .ZN(Mifpw6[5]) );
  NOR2_X1 U897 ( .A1(n679), .A2(n2462), .ZN(Mifpw6[2]) );
  NOR2_X1 U898 ( .A1(n2611), .A2(n5273), .ZN(Tgfpw6[7]) );
  NOR2_X1 U899 ( .A1(n6208), .A2(n6209), .ZN(n6259) );
  AOI22_X1 U900 ( .A1(n6192), .A2(n6189), .B1(n6208), .B2(n6209), .ZN(n6258)
         );
  OR3_X1 U901 ( .A1(n632), .A2(Affpw6[28]), .A3(n2301), .ZN(n5106) );
  OR3_X1 U902 ( .A1(n632), .A2(Affpw6[4]), .A3(n3438), .ZN(n5712) );
  OAI22_X1 U903 ( .A1(n6196), .A2(n6197), .B1(n2790), .B2(n6198), .ZN(n6195)
         );
  OAI22_X1 U904 ( .A1(n6192), .A2(n6193), .B1(n3656), .B2(n3290), .ZN(n6196)
         );
  OAI21_X1 U905 ( .B1(n3287), .B2(n6199), .A(n6190), .ZN(n6197) );
  NOR2_X2 U906 ( .A1(n269), .A2(n3412), .ZN(n2335) );
  NOR2_X2 U907 ( .A1(n232), .A2(n1574), .ZN(n2213) );
  INV_X1 U908 ( .A(n3420), .ZN(n1574) );
  NOR2_X1 U909 ( .A1(n678), .A2(n2370), .ZN(Mifpw6[9]) );
  NOR2_X1 U910 ( .A1(n678), .A2(n2387), .ZN(Mifpw6[11]) );
  NOR2_X1 U911 ( .A1(n4693), .A2(n529), .ZN(n37) );
  NOR2_X1 U912 ( .A1(n678), .A2(n2411), .ZN(Mifpw6[12]) );
  NOR2_X1 U913 ( .A1(n680), .A2(n2406), .ZN(Mifpw6[13]) );
  NAND2_X1 U914 ( .A1(n5694), .A2(n2545), .ZN(n4332) );
  NOR2_X1 U915 ( .A1(n680), .A2(n2403), .ZN(Mifpw6[14]) );
  NAND2_X1 U916 ( .A1(n2730), .A2(n4258), .ZN(n4334) );
  NOR2_X1 U917 ( .A1(n479), .A2(n526), .ZN(n1567) );
  NOR2_X1 U918 ( .A1(n4047), .A2(n2107), .ZN(n3898) );
  OAI22_X1 U919 ( .A1(n4431), .A2(n6311), .B1(n3926), .B2(n3925), .ZN(n6307)
         );
  NOR4_X1 U920 ( .A1(n5812), .A2(n5813), .A3(n3984), .A4(n3983), .ZN(n5806) );
  INV_X1 U921 ( .A(n3558), .ZN(n3984) );
  NAND4_X1 U922 ( .A1(n3449), .A2(n3660), .A3(n3958), .A4(n3612), .ZN(n5812)
         );
  NAND3_X1 U923 ( .A1(n2800), .A2(n3742), .A3(n2685), .ZN(n5813) );
  AOI22_X1 U924 ( .A1(n6193), .A2(n3654), .B1(n6208), .B2(n3290), .ZN(n6198)
         );
  INV_X1 U925 ( .A(n6209), .ZN(n3654) );
  NOR2_X1 U926 ( .A1(n2529), .A2(n4512), .ZN(n1952) );
  NOR4_X1 U927 ( .A1(n522), .A2(n4610), .A3(n1572), .A4(n1571), .ZN(n5230) );
  INV_X1 U928 ( .A(n5693), .ZN(n2544) );
  OAI22_X1 U929 ( .A1(n2730), .A2(n4332), .B1(n2545), .B2(n5694), .ZN(n5693)
         );
  NOR2_X1 U930 ( .A1(n2792), .A2(n2797), .ZN(n5310) );
  AOI22_X1 U931 ( .A1(n3897), .A2(n3898), .B1(n4085), .B2(n1811), .ZN(n407) );
  OR2_X1 U932 ( .A1(n3898), .A2(n1808), .ZN(n4085) );
  NOR3_X1 U933 ( .A1(n4237), .A2(n485), .A3(n5214), .ZN(n5231) );
  INV_X1 U934 ( .A(n5778), .ZN(n2148) );
  OAI21_X1 U935 ( .B1(n5558), .B2(n5779), .A(n5560), .ZN(n5778) );
  NOR4_X1 U936 ( .A1(n3309), .A2(n3072), .A3(n5987), .A4(n2722), .ZN(n5779) );
  INV_X1 U937 ( .A(n5557), .ZN(n2158) );
  OAI21_X1 U938 ( .B1(n5558), .B2(n5559), .A(n5560), .ZN(n5557) );
  NOR3_X1 U939 ( .A1(n5561), .A2(n2725), .A3(n5563), .ZN(n5559) );
  NOR3_X1 U940 ( .A1(n5564), .A2(n5565), .A3(n5566), .ZN(n5563) );
  OAI221_X1 U941 ( .B1(n2429), .B2(n2711), .C1(n4343), .C2(n2389), .A(n4671), 
        .ZN(n252) );
  INV_X1 U942 ( .A(n4346), .ZN(n2711) );
  AOI221_X1 U943 ( .B1(n2350), .B2(n4347), .C1(n4653), .C2(n2383), .A(n4349), 
        .ZN(n4671) );
  NOR3_X1 U944 ( .A1(n503), .A2(n3123), .A3(n2607), .ZN(n1745) );
  OAI221_X1 U945 ( .B1(n3329), .B2(n4153), .C1(n439), .C2(n1604), .A(n4493), 
        .ZN(n3426) );
  AOI211_X1 U946 ( .C1(n4494), .C2(Qbfpw6[25]), .A(Affpw6[25]), .B(n4495), 
        .ZN(n4493) );
  OAI22_X1 U947 ( .A1(n2550), .A2(n2334), .B1(n4446), .B2(n4497), .ZN(n4494)
         );
  NOR3_X1 U948 ( .A1(n2334), .A2(Qbfpw6[25]), .A3(n2549), .ZN(n4495) );
  OAI221_X1 U949 ( .B1(n6189), .B2(n2787), .C1(n5309), .C2(n6190), .A(n6191), 
        .ZN(n6165) );
  NAND3_X1 U950 ( .A1(n3290), .A2(n6192), .A3(n5309), .ZN(n6191) );
  OAI222_X1 U951 ( .A1(n2537), .A2(n1544), .B1(D5epw6), .B2(n2281), .C1(
        Nxkbx6[32]), .C2(Idfpw6[31]), .ZN(n2934) );
  NOR2_X1 U952 ( .A1(n6118), .A2(n6311), .ZN(n5318) );
  NOR2_X1 U953 ( .A1(n4688), .A2(n526), .ZN(n72) );
  NOR2_X1 U954 ( .A1(n2219), .A2(n2226), .ZN(n5453) );
  AOI22_X1 U955 ( .A1(n6118), .A2(n6305), .B1(n3924), .B2(n3056), .ZN(n6180)
         );
  INV_X1 U956 ( .A(n6307), .ZN(n3924) );
  NAND4_X1 U957 ( .A1(n5804), .A2(n5805), .A3(n5806), .A4(n5807), .ZN(n5260)
         );
  NOR4_X1 U958 ( .A1(n5817), .A2(n5818), .A3(n3959), .A4(n3975), .ZN(n5804) );
  NOR4_X1 U959 ( .A1(n5815), .A2(n5816), .A3(n3961), .A4(n3978), .ZN(n5805) );
  NOR4_X1 U960 ( .A1(n5808), .A2(n5809), .A3(n3989), .A4(n3935), .ZN(n5807) );
  OAI21_X1 U961 ( .B1(n5633), .B2(n5634), .A(n242), .ZN(n3901) );
  NAND4_X1 U962 ( .A1(n5653), .A2(n3732), .A3(n4193), .A4(n4263), .ZN(n5633)
         );
  OAI221_X1 U963 ( .B1(n7282), .B2(n3714), .C1(n7355), .C2(n3836), .A(n5651), 
        .ZN(n5634) );
  NAND3_X1 U964 ( .A1(n237), .A2(n7375), .A3(n2563), .ZN(n5653) );
  NAND2_X1 U965 ( .A1(n462), .A2(n3059), .ZN(n1978) );
  NAND2_X1 U966 ( .A1(n5868), .A2(n5255), .ZN(n2357) );
  OAI21_X1 U967 ( .B1(n3047), .B2(n6314), .A(n6118), .ZN(n6185) );
  INV_X1 U968 ( .A(n6315), .ZN(n3047) );
  OAI21_X1 U969 ( .B1(n6181), .B2(n3014), .A(n6182), .ZN(n6166) );
  OAI211_X1 U970 ( .C1(n3015), .C2(n3017), .A(n3014), .B(n6184), .ZN(n6182) );
  INV_X1 U971 ( .A(n6187), .ZN(n3017) );
  NAND3_X1 U972 ( .A1(n3015), .A2(n6185), .A3(n6186), .ZN(n6184) );
  OAI21_X1 U973 ( .B1(n5643), .B2(n3714), .A(n4756), .ZN(n2903) );
  AOI21_X1 U974 ( .B1(n1902), .B2(n3550), .A(n496), .ZN(n5643) );
  NAND2_X1 U975 ( .A1(n5255), .A2(n5244), .ZN(n457) );
  INV_X1 U976 ( .A(n6311), .ZN(n3925) );
  NAND2_X1 U977 ( .A1(n5889), .A2(n5255), .ZN(n3660) );
  OAI22_X1 U978 ( .A1(n6181), .A2(n3016), .B1(n6187), .B2(n6115), .ZN(n6308)
         );
  NOR2_X1 U979 ( .A1(n3221), .A2(n4512), .ZN(n1532) );
  NAND2_X1 U980 ( .A1(n909), .A2(n3844), .ZN(n131) );
  NAND4_X1 U981 ( .A1(n1805), .A2(n1580), .A3(n2121), .A4(n3847), .ZN(n3844)
         );
  NOR2_X1 U982 ( .A1(n3848), .A2(n1979), .ZN(n3847) );
  INV_X1 U983 ( .A(\eq_3147/A[10] ), .ZN(n1718) );
  INV_X1 U984 ( .A(\eq_3147/A[12] ), .ZN(n1693) );
  INV_X1 U985 ( .A(\eq_3147/A[11] ), .ZN(n1709) );
  INV_X1 U986 ( .A(\eq_3147/A[7] ), .ZN(n1769) );
  INV_X1 U987 ( .A(\eq_3147/A[2] ), .ZN(n1793) );
  INV_X1 U988 ( .A(n6143), .ZN(n2792) );
  INV_X1 U989 ( .A(\eq_3147/A[3] ), .ZN(n1788) );
  OAI211_X1 U990 ( .C1(n2528), .C2(n4598), .A(n4073), .B(n5639), .ZN(n5638) );
  AOI221_X1 U991 ( .B1(n4084), .B2(n37), .C1(n5640), .C2(n4263), .A(n5641), 
        .ZN(n5639) );
  NOR3_X1 U992 ( .A1(n2594), .A2(n267), .A3(n516), .ZN(n5641) );
  OAI211_X1 U993 ( .C1(n492), .C2(n2873), .A(n2516), .B(n4204), .ZN(n5640) );
  NAND4_X1 U994 ( .A1(n2824), .A2(n2426), .A3(n4121), .A4(n2472), .ZN(n5815)
         );
  NAND4_X1 U995 ( .A1(n2357), .A2(n3644), .A3(n3649), .A4(n2526), .ZN(n5817)
         );
  NAND4_X1 U996 ( .A1(n2536), .A2(n3862), .A3(n4843), .A4(n3639), .ZN(n5808)
         );
  INV_X1 U997 ( .A(\eq_3147/A[9] ), .ZN(n1738) );
  INV_X1 U998 ( .A(\eq_3147/A[8] ), .ZN(n1766) );
  INV_X1 U999 ( .A(\eq_3147/A[6] ), .ZN(n1774) );
  INV_X1 U1000 ( .A(\eq_3147/A[5] ), .ZN(n1780) );
  INV_X1 U1001 ( .A(\eq_3147/A[4] ), .ZN(n1785) );
  INV_X1 U1002 ( .A(n6118), .ZN(n3056) );
  INV_X1 U1003 ( .A(n5838), .ZN(n3983) );
  INV_X1 U1004 ( .A(n4497), .ZN(n2334) );
  INV_X1 U1005 ( .A(n2806), .ZN(n3551) );
  INV_X1 U1006 ( .A(\eq_3147/A[1] ), .ZN(n1798) );
  NAND3_X1 U1007 ( .A1(n242), .A2(n4521), .A3(n5199), .ZN(n3891) );
  INV_X1 U1008 ( .A(n5457), .ZN(n2219) );
  INV_X1 U1009 ( .A(n5303), .ZN(n3659) );
  NAND4_X1 U1010 ( .A1(n1610), .A2(n1606), .A3(n149), .A4(n150), .ZN(n139) );
  NOR4_X1 U1011 ( .A1(\eq_3147/A[20] ), .A2(\eq_3147/A[19] ), .A3(
        \eq_3147/A[18] ), .A4(\eq_3147/A[17] ), .ZN(n150) );
  NOR3_X1 U1012 ( .A1(\eq_3147/A[23] ), .A2(\eq_3147/A[25] ), .A3(
        \eq_3147/A[24] ), .ZN(n149) );
  AOI22_X1 U1013 ( .A1(n6115), .A2(n6301), .B1(n6172), .B2(n6302), .ZN(n5316)
         );
  OAI22_X1 U1014 ( .A1(n6303), .A2(n6180), .B1(n6304), .B2(n6179), .ZN(n6302)
         );
  AND2_X1 U1015 ( .A1(n6179), .A2(n6304), .ZN(n6303) );
  NAND3_X1 U1016 ( .A1(n6308), .A2(n6185), .A3(n6186), .ZN(n6304) );
  INV_X1 U1017 ( .A(n6115), .ZN(n3016) );
  INV_X1 U1018 ( .A(n3579), .ZN(n3959) );
  INV_X1 U1019 ( .A(n4039), .ZN(n3975) );
  INV_X1 U1020 ( .A(n5648), .ZN(n3566) );
  NOR2_X1 U1021 ( .A1(n678), .A2(n2384), .ZN(Mifpw6[10]) );
  AND3_X1 U1022 ( .A1(n4271), .A2(n2548), .A3(n5199), .ZN(n3283) );
  NAND3_X1 U1023 ( .A1(n3597), .A2(n3778), .A3(n1636), .ZN(n5816) );
  INV_X1 U1024 ( .A(n111), .ZN(n1527) );
  INV_X1 U1025 ( .A(n124), .ZN(n1526) );
  OR2_X1 U1026 ( .A1(n669), .A2(n5626), .ZN(n3900) );
  AOI211_X1 U1027 ( .C1(n1624), .C2(n7375), .A(n5627), .B(n5628), .ZN(n5626)
         );
  OAI222_X1 U1028 ( .A1(n508), .A2(n3828), .B1(n272), .B2(n2873), .C1(n7373), 
        .C2(n3737), .ZN(n5627) );
  INV_X1 U1029 ( .A(n3199), .ZN(n3989) );
  INV_X1 U1030 ( .A(n3742), .ZN(n3986) );
  INV_X1 U1031 ( .A(n466), .ZN(n1811) );
  INV_X1 U1032 ( .A(n3677), .ZN(n3978) );
  INV_X1 U1033 ( .A(n3639), .ZN(n3973) );
  INV_X1 U1034 ( .A(n3644), .ZN(n3977) );
  INV_X1 U1035 ( .A(n3958), .ZN(n3971) );
  INV_X1 U1036 ( .A(n3612), .ZN(n3985) );
  INV_X1 U1037 ( .A(n4013), .ZN(n3939) );
  INV_X1 U1038 ( .A(n2536), .ZN(n3934) );
  INV_X1 U1039 ( .A(n3597), .ZN(n3951) );
  INV_X1 U1040 ( .A(n3624), .ZN(n3955) );
  INV_X1 U1041 ( .A(n4472), .ZN(n3961) );
  INV_X1 U1042 ( .A(n3542), .ZN(n3935) );
  INV_X1 U1043 ( .A(n3649), .ZN(n3946) );
  INV_X1 U1044 ( .A(n6205), .ZN(n2794) );
  INV_X1 U1045 ( .A(n3862), .ZN(n3987) );
  AND2_X1 U1046 ( .A1(n5658), .A2(n5560), .ZN(n5602) );
  OAI22_X1 U1047 ( .A1(n2722), .A2(n3080), .B1(n5659), .B2(n5564), .ZN(n5658)
         );
  AOI211_X1 U1048 ( .C1(n5013), .C2(n265), .A(n5558), .B(n5660), .ZN(n5659) );
  NOR3_X1 U1049 ( .A1(n4193), .A2(n225), .A3(n7375), .ZN(n5660) );
  INV_X1 U1050 ( .A(n6350), .ZN(n3063) );
  NAND4_X1 U1051 ( .A1(n2752), .A2(n2606), .A3(n5238), .A4(n5239), .ZN(n5235)
         );
  AOI221_X1 U1052 ( .B1(n1763), .B2(n3466), .C1(n1761), .C2(n5240), .A(n5241), 
        .ZN(n5239) );
  INV_X1 U1053 ( .A(n1745), .ZN(n2606) );
  OR3_X1 U1054 ( .A1(n4610), .A2(n522), .A3(n1572), .ZN(n5238) );
  OR3_X1 U1055 ( .A1(n3426), .A2(n3427), .A3(n3428), .ZN(n3423) );
  NAND2_X1 U1056 ( .A1(n4013), .A2(n3624), .ZN(n5818) );
  INV_X1 U1057 ( .A(n6316), .ZN(n3635) );
  NOR3_X1 U1059 ( .A1(n4633), .A2(n4512), .A3(n265), .ZN(n5635) );
  INV_X1 U1060 ( .A(n4235), .ZN(n4204) );
  NOR2_X1 U1061 ( .A1(n2611), .A2(n2360), .ZN(Mifpw6[6]) );
  INV_X1 U1062 ( .A(n5803), .ZN(n2216) );
  NOR2_X1 U1063 ( .A1(n2611), .A2(n2365), .ZN(Mifpw6[7]) );
  NOR2_X1 U1064 ( .A1(n678), .A2(n2367), .ZN(Mifpw6[8]) );
  INV_X1 U1065 ( .A(n839), .ZN(n2088) );
  NOR2_X1 U1066 ( .A1(n2164), .A2(n792), .ZN(n763) );
  NOR2_X2 U1067 ( .A1(n319), .A2(n3400), .ZN(n2248) );
  NOR2_X2 U1068 ( .A1(n375), .A2(n3428), .ZN(n2255) );
  NOR2_X1 U1069 ( .A1(n2699), .A2(n475), .ZN(n1584) );
  INV_X1 U1070 ( .A(n449), .ZN(n2124) );
  NOR2_X1 U1071 ( .A1(n1006), .A2(n741), .ZN(n884) );
  NOR2_X1 U1072 ( .A1(n1023), .A2(n741), .ZN(n877) );
  NOR2_X1 U1073 ( .A1(n475), .A2(n2124), .ZN(n1674) );
  NOR2_X1 U1074 ( .A1(n680), .A2(n2413), .ZN(Mifpw6[15]) );
  NAND4_X1 U1075 ( .A1(n2522), .A2(n4073), .A3(n4074), .A4(n4075), .ZN(n202)
         );
  AOI22_X1 U1076 ( .A1(n37), .A2(n4082), .B1(n496), .B2(n1730), .ZN(n4074) );
  NOR4_X1 U1077 ( .A1(n4076), .A2(n4077), .A3(n3767), .A4(n4079), .ZN(n4075)
         );
  INV_X1 U1078 ( .A(n1931), .ZN(n2522) );
  INV_X1 U1079 ( .A(n798), .ZN(n2167) );
  NOR2_X1 U1080 ( .A1(n680), .A2(n2397), .ZN(Mifpw6[16]) );
  INV_X1 U1081 ( .A(n3050), .ZN(n1815) );
  AOI222_X1 U1082 ( .A1(n269), .A2(n99), .B1(n462), .B2(n3051), .C1(n2512), 
        .C2(Nxkbx6[1]), .ZN(n3050) );
  NOR2_X1 U1083 ( .A1(n680), .A2(n2392), .ZN(Mifpw6[17]) );
  NOR2_X1 U1084 ( .A1(n5063), .A2(n270), .ZN(n1908) );
  NOR2_X1 U1086 ( .A1(n470), .A2(n2277), .ZN(n1751) );
  AND3_X1 U1087 ( .A1(n3395), .A2(n5149), .A3(n282), .ZN(n2325) );
  NOR2_X1 U1088 ( .A1(n5457), .A2(n2224), .ZN(n4789) );
  NOR3_X1 U1089 ( .A1(n4265), .A2(n4232), .A3(n2509), .ZN(n1749) );
  NOR2_X1 U1090 ( .A1(n680), .A2(n2390), .ZN(Mifpw6[18]) );
  AOI22_X1 U1091 ( .A1(n5652), .A2(n516), .B1(n493), .B2(n508), .ZN(n5651) );
  NAND2_X1 U1092 ( .A1(n492), .A2(n4650), .ZN(n5652) );
  INV_X1 U1093 ( .A(n806), .ZN(n2163) );
  INV_X1 U1094 ( .A(n4851), .ZN(n2692) );
  AOI22_X1 U1095 ( .A1(n6115), .A2(n6316), .B1(n3018), .B2(n3016), .ZN(n6179)
         );
  NOR2_X1 U1096 ( .A1(n680), .A2(n2400), .ZN(Mifpw6[19]) );
  AND2_X1 U1097 ( .A1(n2140), .A2(n3433), .ZN(n2288) );
  OAI22_X1 U1098 ( .A1(n2524), .A2(n3787), .B1(n2528), .B2(n4083), .ZN(n1931)
         );
  NAND2_X1 U1099 ( .A1(n1620), .A2(n492), .ZN(n4083) );
  NOR2_X1 U1100 ( .A1(n990), .A2(n741), .ZN(n1125) );
  INV_X1 U1101 ( .A(n1685), .ZN(n2699) );
  NOR2_X1 U1102 ( .A1(n741), .A2(n1009), .ZN(n1124) );
  NOR2_X1 U1103 ( .A1(n265), .A2(n485), .ZN(n4084) );
  NOR2_X1 U1104 ( .A1(n680), .A2(n2440), .ZN(Mifpw6[20]) );
  NAND3_X1 U1105 ( .A1(n4789), .A2(n4790), .A3(n4791), .ZN(n756) );
  AOI22_X1 U1106 ( .A1(n6143), .A2(n6205), .B1(n6206), .B2(n2792), .ZN(n6199)
         );
  NOR2_X1 U1107 ( .A1(n230), .A2(n479), .ZN(n2496) );
  NAND3_X1 U1108 ( .A1(n3897), .A2(n466), .A3(n3898), .ZN(n3920) );
  NAND3_X1 U1109 ( .A1(n485), .A2(n491), .A3(n1626), .ZN(n2752) );
  NOR2_X1 U1110 ( .A1(n680), .A2(n2438), .ZN(Mifpw6[21]) );
  NOR2_X1 U1111 ( .A1(n4512), .A2(n492), .ZN(n1723) );
  INV_X1 U1112 ( .A(n473), .ZN(n2260) );
  NOR3_X1 U1113 ( .A1(n4610), .A2(n486), .A3(n479), .ZN(n5249) );
  NOR3_X1 U1114 ( .A1(n3800), .A2(n529), .A3(n265), .ZN(n5241) );
  OAI21_X1 U1115 ( .B1(n5974), .B2(n2212), .A(n4791), .ZN(n752) );
  AOI22_X1 U1116 ( .A1(n2783), .A2(n5316), .B1(n5309), .B2(n4790), .ZN(n5974)
         );
  NOR2_X1 U1117 ( .A1(n680), .A2(n2437), .ZN(Mifpw6[22]) );
  NAND3_X1 U1118 ( .A1(n4789), .A2(n2783), .A3(n4791), .ZN(n754) );
  OAI22_X1 U1119 ( .A1(n3788), .A2(n4738), .B1(n4265), .B2(n2873), .ZN(n5232)
         );
  NAND2_X1 U1120 ( .A1(n792), .A2(n798), .ZN(n796) );
  NOR2_X1 U1121 ( .A1(n680), .A2(n2442), .ZN(Mifpw6[23]) );
  INV_X1 U1122 ( .A(n6127), .ZN(n3019) );
  INV_X1 U1123 ( .A(n856), .ZN(n2098) );
  INV_X1 U1124 ( .A(n2395), .ZN(n3895) );
  INV_X1 U1125 ( .A(n1672), .ZN(n1945) );
  INV_X1 U1126 ( .A(n4047), .ZN(n2693) );
  NAND2_X1 U1127 ( .A1(n5310), .A2(n6211), .ZN(n6171) );
  OR2_X1 U1128 ( .A1(n5214), .A2(n265), .ZN(n2072) );
  AOI21_X1 U1129 ( .B1(n2107), .B2(n1986), .A(n3891), .ZN(n3889) );
  INV_X1 U1130 ( .A(n2952), .ZN(n3682) );
  NAND2_X1 U1131 ( .A1(n7373), .A2(n516), .ZN(n3055) );
  INV_X1 U1132 ( .A(n4350), .ZN(n2138) );
  NAND2_X1 U1133 ( .A1(n6318), .A2(n6118), .ZN(n6172) );
  NOR2_X1 U1134 ( .A1(n4512), .A2(n3714), .ZN(n4091) );
  OR2_X1 U1135 ( .A1(n985), .A2(n741), .ZN(n727) );
  OR2_X1 U1136 ( .A1(n989), .A2(n741), .ZN(n728) );
  INV_X1 U1137 ( .A(n501), .ZN(n3686) );
  INV_X1 U1138 ( .A(n379), .ZN(n2145) );
  INV_X1 U1139 ( .A(n453), .ZN(n2139) );
  INV_X1 U1140 ( .A(n1571), .ZN(n1994) );
  INV_X1 U1141 ( .A(n3051), .ZN(n2140) );
  AND3_X1 U1142 ( .A1(n1723), .A2(n7282), .A3(n474), .ZN(n4077) );
  INV_X1 U1143 ( .A(n6375), .ZN(n3272) );
  AND2_X1 U1144 ( .A1(n6261), .A2(n3659), .ZN(n6194) );
  INV_X1 U1145 ( .A(n6366), .ZN(n3018) );
  INV_X1 U1146 ( .A(n4081), .ZN(n2517) );
  INV_X1 U1147 ( .A(n6189), .ZN(n3656) );
  INV_X1 U1149 ( .A(Nxkbx6[1]), .ZN(n1814) );
  INV_X1 U1150 ( .A(n6277), .ZN(n3866) );
  INV_X1 U1151 ( .A(n259), .ZN(n2130) );
  AOI21_X1 U1152 ( .B1(n906), .B2(n3765), .A(n963), .ZN(n677) );
  INV_X1 U1153 ( .A(n3327), .ZN(n3105) );
  NOR2_X1 U1154 ( .A1(n963), .A2(n477), .ZN(n1643) );
  NOR3_X1 U1155 ( .A1(n3111), .A2(n3305), .A3(n4556), .ZN(n3354) );
  INV_X1 U1156 ( .A(n1966), .ZN(HALTED) );
  OR3_X1 U1157 ( .A1(n3382), .A2(n3327), .A3(n3383), .ZN(n3376) );
  OR3_X1 U1158 ( .A1(n3380), .A2(n3105), .A3(n3381), .ZN(n3377) );
  AOI22_X1 U1159 ( .A1(n6127), .A2(n3274), .B1(n3024), .B2(n3019), .ZN(n6114)
         );
  NOR3_X1 U1161 ( .A1(n6118), .A2(n3928), .A3(n3925), .ZN(n6117) );
  OAI22_X1 U1162 ( .A1(n4432), .A2(n3060), .B1(n3056), .B2(n6123), .ZN(n6116)
         );
  OAI21_X1 U1163 ( .B1(n4137), .B2(n4119), .A(n1361), .ZN(n720) );
  OAI22_X1 U1164 ( .A1(n3105), .A2(n3326), .B1(n3327), .B2(n3340), .ZN(n3315)
         );
  INV_X1 U1165 ( .A(n731), .ZN(n729) );
  INV_X1 U1166 ( .A(n731), .ZN(n722) );
  OAI221_X1 U1167 ( .B1(n5280), .B2(n5675), .C1(n3108), .C2(n3358), .A(n4762), 
        .ZN(n4735) );
  INV_X1 U1168 ( .A(n398), .ZN(n872) );
  AOI22_X1 U1169 ( .A1(n3327), .A2(n2366), .B1(n3105), .B2(n2402), .ZN(n3359)
         );
  OAI21_X1 U1170 ( .B1(n3166), .B2(n3167), .A(N701), .ZN(n2408) );
  OAI211_X1 U1171 ( .C1(n3714), .C2(n4602), .A(n3168), .B(n3169), .ZN(n3167)
         );
  NAND4_X1 U1172 ( .A1(n3182), .A2(n3183), .A3(n3184), .A4(n3185), .ZN(n3166)
         );
  AOI211_X1 U1173 ( .C1(n3170), .C2(n875), .A(n3171), .B(n3172), .ZN(n3169) );
  NOR2_X1 U1174 ( .A1(n5174), .A2(n2582), .ZN(n4748) );
  OAI21_X1 U1175 ( .B1(n3327), .B2(n3378), .A(n3087), .ZN(n3338) );
  INV_X1 U1176 ( .A(n5271), .ZN(n3087) );
  OAI21_X1 U1177 ( .B1(n3327), .B2(n4731), .A(n3102), .ZN(n3342) );
  OAI21_X1 U1178 ( .B1(n3327), .B2(n5674), .A(n4735), .ZN(n3336) );
  OAI22_X1 U1179 ( .A1(n3327), .A2(n3381), .B1(n3105), .B2(n5395), .ZN(n3373)
         );
  OAI22_X1 U1180 ( .A1(n3323), .A2(n3327), .B1(n3105), .B2(n3361), .ZN(n4549)
         );
  AOI211_X1 U1181 ( .C1(HALTED), .C2(n876), .A(n877), .B(n2000), .ZN(n867) );
  OAI21_X1 U1182 ( .B1(n3327), .B2(n3339), .A(n3101), .ZN(n3344) );
  OAI22_X1 U1183 ( .A1(n3105), .A2(n3360), .B1(n3327), .B2(n3325), .ZN(n3314)
         );
  INV_X1 U1185 ( .A(n1361), .ZN(n1998) );
  OAI211_X1 U1186 ( .C1(n524), .C2(n6545), .A(n2072), .B(n6546), .ZN(n6529) );
  AOI222_X1 U1187 ( .A1(n1520), .A2(n7373), .B1(n52), .B2(n265), .C1(n5253), 
        .C2(n463), .ZN(n6545) );
  AOI22_X1 U1188 ( .A1(n1642), .A2(n2743), .B1(n4582), .B2(n1539), .ZN(n6546)
         );
  OAI22_X1 U1190 ( .A1(n3327), .A2(n3380), .B1(n3105), .B2(n5674), .ZN(n4547)
         );
  INV_X1 U1191 ( .A(n354), .ZN(n3712) );
  OAI22_X1 U1192 ( .A1(n3327), .A2(n3368), .B1(n3105), .B2(n3382), .ZN(n3374)
         );
  OAI21_X1 U1193 ( .B1(n228), .B2(n4616), .A(n5923), .ZN(n4458) );
  NAND3_X1 U1194 ( .A1(n1520), .A2(n7282), .A3(n4092), .ZN(n5923) );
  NOR2_X1 U1195 ( .A1(n3369), .A2(n3351), .ZN(n4734) );
  NAND4_X1 U1196 ( .A1(n5280), .A2(n6041), .A3(n3327), .A4(n4556), .ZN(n6033)
         );
  NAND4_X1 U1197 ( .A1(n6539), .A2(n1911), .A3(n6540), .A4(n6541), .ZN(n6530)
         );
  OAI211_X1 U1198 ( .C1(n493), .C2(n491), .A(n1528), .B(n6544), .ZN(n6539) );
  AOI221_X1 U1199 ( .B1(n2915), .B2(n482), .C1(n1642), .C2(n523), .A(n5738), 
        .ZN(n6541) );
  AOI22_X1 U1200 ( .A1(n6543), .A2(n4263), .B1(n1462), .B2(n1463), .ZN(n6540)
         );
  NOR4_X1 U1202 ( .A1(n344), .A2(n2632), .A3(n2676), .A4(n2671), .ZN(n4846) );
  NOR2_X1 U1203 ( .A1(n963), .A2(n1986), .ZN(n409) );
  NOR4_X1 U1204 ( .A1(n3078), .A2(n4565), .A3(n3080), .A4(n2444), .ZN(n4570)
         );
  NOR2_X1 U1205 ( .A1(n5622), .A2(n2464), .ZN(n4401) );
  NOR3_X1 U1206 ( .A1(n6041), .A2(n3305), .A3(n4556), .ZN(n5987) );
  OAI221_X1 U1207 ( .B1(n2428), .B2(n3342), .C1(n2425), .C2(n3344), .A(n3345), 
        .ZN(n3331) );
  INV_X1 U1208 ( .A(n3318), .ZN(n2425) );
  AOI221_X1 U1209 ( .B1(n3346), .B2(n2349), .C1(n3105), .C2(n3348), .A(n3349), 
        .ZN(n3345) );
  NAND4_X1 U1210 ( .A1(n3344), .A2(n3336), .A3(n3342), .A4(n3338), .ZN(n3348)
         );
  OAI211_X1 U1211 ( .C1(n7375), .C2(n3746), .A(n6567), .B(n6568), .ZN(n6534)
         );
  NAND4_X1 U1212 ( .A1(n417), .A2(n3509), .A3(n266), .A4(n4263), .ZN(n6567) );
  NAND4_X1 U1213 ( .A1(n2915), .A2(n517), .A3(n433), .A4(n225), .ZN(n6568) );
  NOR2_X1 U1214 ( .A1(n2595), .A2(n2464), .ZN(n5172) );
  NAND4_X1 U1215 ( .A1(n5919), .A2(n5920), .A3(n6531), .A4(n6532), .ZN(n5174)
         );
  AND2_X1 U1216 ( .A1(N701), .A2(n5921), .ZN(n6532) );
  INV_X1 U1217 ( .A(n5392), .ZN(n2418) );
  OAI22_X1 U1218 ( .A1(n3105), .A2(n3328), .B1(n3327), .B2(n5393), .ZN(n5392)
         );
  AOI21_X1 U1219 ( .B1(n2610), .B2(n97), .A(n961), .ZN(n3294) );
  AND2_X1 U1220 ( .A1(n1410), .A2(n3488), .ZN(n715) );
  XOR2_X1 U1221 ( .A(n384), .B(n4561), .Z(n6041) );
  NOR2_X1 U1222 ( .A1(n517), .A2(n4559), .ZN(n384) );
  NOR2_X1 U1223 ( .A1(n988), .A2(n741), .ZN(n1080) );
  AOI211_X1 U1224 ( .C1(n1567), .C2(n536), .A(n2592), .B(n2593), .ZN(n2555) );
  OAI22_X1 U1225 ( .A1(n3835), .A2(n4602), .B1(n3714), .B2(n4205), .ZN(n2592)
         );
  OAI22_X1 U1226 ( .A1(n2444), .A2(n5992), .B1(n3086), .B2(n5994), .ZN(n3333)
         );
  AOI22_X1 U1227 ( .A1(n5393), .A2(n3327), .B1(n3105), .B2(n5395), .ZN(n5994)
         );
  INV_X1 U1228 ( .A(n5992), .ZN(n3086) );
  NAND2_X1 U1229 ( .A1(n4762), .A2(n5675), .ZN(n5992) );
  NAND4_X1 U1230 ( .A1(N701), .A2(n3514), .A3(n3515), .A4(n3122), .ZN(n2593)
         );
  NAND3_X1 U1231 ( .A1(n4512), .A2(n491), .A3(n7375), .ZN(n3514) );
  NOR2_X1 U1232 ( .A1(n3831), .A2(n526), .ZN(n1747) );
  INV_X1 U1233 ( .A(n4397), .ZN(n2703) );
  BUF_X1 U1234 ( .A(n1861), .Z(n866) );
  OAI221_X1 U1235 ( .B1(n4552), .B2(n3111), .C1(n4550), .C2(n3314), .A(n4553), 
        .ZN(n4551) );
  NAND3_X1 U1236 ( .A1(n3111), .A2(n3110), .A3(n2418), .ZN(n4553) );
  AOI22_X1 U1237 ( .A1(n2346), .A2(n4556), .B1(n3359), .B2(n3110), .ZN(n4552)
         );
  INV_X1 U1238 ( .A(n3373), .ZN(n2346) );
  BUF_X1 U1239 ( .A(n3872), .Z(n670) );
  INV_X1 U1240 ( .A(n1376), .ZN(n2118) );
  AOI22_X1 U1241 ( .A1(n2444), .A2(n5947), .B1(n3096), .B2(n4547), .ZN(n3349)
         );
  INV_X1 U1242 ( .A(n5947), .ZN(n3096) );
  AOI21_X1 U1243 ( .B1(n3358), .B2(n3108), .A(n5495), .ZN(n5947) );
  AOI21_X1 U1244 ( .B1(n524), .B2(n3712), .A(n961), .ZN(n1982) );
  NOR3_X1 U1245 ( .A1(n3828), .A2(n529), .A3(n4610), .ZN(n4359) );
  OAI211_X1 U1246 ( .C1(n3358), .C2(n3103), .A(n5675), .B(n523), .ZN(n5495) );
  NAND3_X1 U1247 ( .A1(n6485), .A2(n3351), .A3(n3112), .ZN(n6447) );
  INV_X1 U1248 ( .A(n1050), .ZN(n2002) );
  NOR3_X1 U1249 ( .A1(n2506), .A2(n4237), .A3(n4265), .ZN(n4360) );
  NAND2_X1 U1250 ( .A1(N701), .A2(n3059), .ZN(n461) );
  OAI21_X1 U1251 ( .B1(n522), .B2(n4738), .A(n4685), .ZN(n2870) );
  INV_X1 U1252 ( .A(n4556), .ZN(n3110) );
  OAI21_X1 U1253 ( .B1(n7282), .B2(n2591), .A(n3055), .ZN(n6533) );
  OAI22_X1 U1254 ( .A1(n2433), .A2(n3336), .B1(n2449), .B2(n3338), .ZN(n3332)
         );
  INV_X1 U1255 ( .A(n3340), .ZN(n2433) );
  INV_X1 U1256 ( .A(n3339), .ZN(n2449) );
  NAND2_X1 U1257 ( .A1(n883), .A2(n999), .ZN(n732) );
  OAI22_X1 U1258 ( .A1(n2549), .A2(N3epw6), .B1(n2550), .B2(n4422), .ZN(n4421)
         );
  OAI22_X1 U1259 ( .A1(n2549), .A2(U3epw6), .B1(n2550), .B2(n5608), .ZN(n5607)
         );
  OAI22_X1 U1260 ( .A1(n2549), .A2(I4epw6), .B1(n2550), .B2(n4600), .ZN(n4599)
         );
  OAI22_X1 U1261 ( .A1(n2549), .A2(B4epw6), .B1(n2550), .B2(n4660), .ZN(n4659)
         );
  OAI22_X1 U1262 ( .A1(n2549), .A2(L2epw6), .B1(n2550), .B2(n4480), .ZN(n4479)
         );
  OAI22_X1 U1263 ( .A1(n2549), .A2(Z2epw6), .B1(n2550), .B2(n5072), .ZN(n5071)
         );
  NOR2_X1 U1264 ( .A1(n6143), .A2(n3117), .ZN(n5311) );
  OAI22_X1 U1265 ( .A1(n505), .A2(n3831), .B1(n479), .B2(n4591), .ZN(n6543) );
  AND2_X1 U1266 ( .A1(n732), .A2(n1050), .ZN(n901) );
  INV_X1 U1267 ( .A(n909), .ZN(n2102) );
  NOR2_X1 U1268 ( .A1(n679), .A2(n2419), .ZN(Mifpw6[24]) );
  NAND2_X1 U1269 ( .A1(n3111), .A2(n4556), .ZN(n4550) );
  NAND2_X1 U1270 ( .A1(n1293), .A2(n4119), .ZN(n1166) );
  OAI211_X1 U1271 ( .C1(n3304), .C2(n3305), .A(n3306), .B(n3307), .ZN(n3303)
         );
  OAI21_X1 U1272 ( .B1(n3309), .B2(n3080), .A(n3330), .ZN(n3306) );
  NOR4_X1 U1273 ( .A1(n3331), .A2(n3332), .A3(n3333), .A4(n3334), .ZN(n3304)
         );
  OAI211_X1 U1274 ( .C1(n210), .C2(n275), .A(n3054), .B(n2548), .ZN(n3053) );
  NAND3_X1 U1275 ( .A1(n3055), .A2(n3836), .A3(n3057), .ZN(n3054) );
  AOI22_X1 U1276 ( .A1(n521), .A2(n477), .B1(n508), .B2(n516), .ZN(n3057) );
  NAND3_X1 U1277 ( .A1(n3350), .A2(n2444), .A3(n3352), .ZN(n3302) );
  NAND3_X1 U1278 ( .A1(n3330), .A2(n3353), .A3(n3354), .ZN(n3352) );
  NAND3_X1 U1279 ( .A1(n3373), .A2(n3374), .A3(n3375), .ZN(n3370) );
  NAND3_X1 U1280 ( .A1(n6531), .A2(n2607), .A3(N701), .ZN(n6536) );
  NAND3_X1 U1281 ( .A1(n5426), .A2(n2543), .A3(n4446), .ZN(n5425) );
  INV_X1 U1282 ( .A(Qbfpw6[30]), .ZN(n2543) );
  AND2_X1 U1283 ( .A1(n2582), .A2(n5174), .ZN(n4609) );
  NAND2_X1 U1284 ( .A1(n1107), .A2(n4119), .ZN(n840) );
  NAND3_X1 U1285 ( .A1(n872), .A2(n2977), .A3(n1887), .ZN(n1858) );
  NOR2_X1 U1286 ( .A1(n679), .A2(n2427), .ZN(Mifpw6[25]) );
  OAI21_X1 U1287 ( .B1(n99), .B2(n3049), .A(N701), .ZN(n3052) );
  AND3_X1 U1288 ( .A1(n3712), .A2(n1376), .A3(n1431), .ZN(n1410) );
  INV_X1 U1289 ( .A(n6498), .ZN(n3369) );
  INV_X1 U1290 ( .A(D5epw6), .ZN(n2537) );
  NAND2_X1 U1291 ( .A1(n203), .A2(n202), .ZN(n4064) );
  INV_X1 U1292 ( .A(n1916), .ZN(n1837) );
  NAND2_X1 U1293 ( .A1(n1361), .A2(n720), .ZN(n719) );
  NAND3_X1 U1294 ( .A1(n3314), .A2(n3315), .A3(n3316), .ZN(n3311) );
  OR3_X1 U1295 ( .A1(n3326), .A2(n3327), .A3(n3328), .ZN(n3317) );
  OR3_X1 U1296 ( .A1(n3323), .A2(n3105), .A3(n3325), .ZN(n3320) );
  INV_X1 U1297 ( .A(n5127), .ZN(n2345) );
  OAI21_X1 U1298 ( .B1(N701), .B2(n405), .A(n406), .ZN(n7825) );
  AOI21_X1 U1299 ( .B1(n4157), .B2(n410), .A(n4512), .ZN(n405) );
  NAND3_X1 U1300 ( .A1(n407), .A2(n242), .A3(n409), .ZN(n406) );
  NAND4_X1 U1301 ( .A1(n411), .A2(n412), .A3(n413), .A4(n414), .ZN(n410) );
  NAND2_X1 U1302 ( .A1(n3355), .A2(n3356), .ZN(n3330) );
  AOI211_X1 U1303 ( .C1(n3362), .C2(n3327), .A(n3363), .B(n3364), .ZN(n3355)
         );
  AOI211_X1 U1304 ( .C1(n3105), .C2(n3357), .A(n2391), .B(n3359), .ZN(n3356)
         );
  OR4_X1 U1305 ( .A1(n3365), .A2(n3366), .A3(n3367), .A4(n3368), .ZN(n3362) );
  INV_X1 U1306 ( .A(n5280), .ZN(n3358) );
  INV_X1 U1307 ( .A(n5553), .ZN(n2398) );
  INV_X1 U1308 ( .A(n4837), .ZN(n2385) );
  INV_X1 U1309 ( .A(n4412), .ZN(n2350) );
  NOR2_X1 U1310 ( .A1(n679), .A2(n2432), .ZN(Mifpw6[26]) );
  INV_X1 U1311 ( .A(n5487), .ZN(n2349) );
  AOI22_X1 U1312 ( .A1(n3379), .A2(n3105), .B1(n3327), .B2(n4731), .ZN(n5487)
         );
  INV_X1 U1313 ( .A(n5622), .ZN(n2595) );
  INV_X1 U1314 ( .A(n1694), .ZN(n1885) );
  NAND3_X1 U1315 ( .A1(n4256), .A2(n2538), .A3(n2293), .ZN(n4809) );
  BUF_X1 U1316 ( .A(n399), .Z(n787) );
  NOR2_X1 U1317 ( .A1(n679), .A2(n2447), .ZN(Mifpw6[31]) );
  OR4_X1 U1318 ( .A1(n3322), .A2(n3321), .A3(n3360), .A4(n3361), .ZN(n3357) );
  INV_X1 U1319 ( .A(n4416), .ZN(n2389) );
  INV_X1 U1320 ( .A(n4654), .ZN(n2415) );
  NAND3_X1 U1321 ( .A1(n5919), .A2(n5920), .A3(n5921), .ZN(n5918) );
  NOR2_X1 U1322 ( .A1(n679), .A2(n2436), .ZN(Mifpw6[27]) );
  INV_X1 U1323 ( .A(n3319), .ZN(n2428) );
  NAND2_X1 U1324 ( .A1(n4521), .A2(n6542), .ZN(n5738) );
  NAND3_X1 U1325 ( .A1(n1567), .A2(n875), .A3(n2915), .ZN(n6542) );
  NAND2_X1 U1326 ( .A1(n4400), .A2(n4401), .ZN(n2210) );
  NAND2_X1 U1327 ( .A1(n4612), .A2(n4748), .ZN(n2214) );
  NAND2_X1 U1328 ( .A1(n4612), .A2(n4400), .ZN(n2231) );
  INV_X1 U1329 ( .A(n3367), .ZN(n2402) );
  NAND2_X1 U1330 ( .A1(n4407), .A2(n4400), .ZN(n2253) );
  NAND2_X1 U1331 ( .A1(n4407), .A2(n5087), .ZN(n2229) );
  NAND2_X1 U1332 ( .A1(n4407), .A2(n4748), .ZN(n2348) );
  INV_X1 U1333 ( .A(n2152), .ZN(n1989) );
  INV_X1 U1334 ( .A(n3383), .ZN(n2366) );
  INV_X1 U1335 ( .A(Qbfpw6[29]), .ZN(n2538) );
  NAND2_X1 U1336 ( .A1(n5172), .A2(n5087), .ZN(n2362) );
  NAND2_X1 U1337 ( .A1(n5172), .A2(n4400), .ZN(n2249) );
  INV_X1 U1338 ( .A(Qbfpw6[24]), .ZN(n2541) );
  NOR2_X1 U1339 ( .A1(n679), .A2(n2457), .ZN(Mifpw6[28]) );
  OR2_X1 U1340 ( .A1(n6498), .A2(n3351), .ZN(n387) );
  AOI21_X1 U1341 ( .B1(n7373), .B2(n961), .A(n3490), .ZN(Jrohu6) );
  AND4_X1 U1342 ( .A1(n3491), .A2(n3492), .A3(n3493), .A4(n3494), .ZN(n3490)
         );
  AOI211_X1 U1343 ( .C1(n1674), .C2(n3500), .A(n3501), .B(n3502), .ZN(n3493)
         );
  AOI221_X1 U1345 ( .B1(n1747), .B2(n514), .C1(n3786), .C2(n1974), .A(n3506), 
        .ZN(n3492) );
  NAND2_X1 U1346 ( .A1(n4609), .A2(n4612), .ZN(n2315) );
  NAND2_X1 U1347 ( .A1(n5087), .A2(n4612), .ZN(n2218) );
  NAND2_X1 U1348 ( .A1(n4609), .A2(n4407), .ZN(n2344) );
  NOR2_X1 U1349 ( .A1(n679), .A2(n2456), .ZN(Mifpw6[29]) );
  NOR2_X1 U1350 ( .A1(n679), .A2(n2451), .ZN(Mifpw6[30]) );
  AND3_X1 U1351 ( .A1(n1812), .A2(n2297), .A3(Ntkbx6[0]), .ZN(Gwhhu6) );
  AND3_X1 U1352 ( .A1(n1812), .A2(n2264), .A3(Nvkbx6[0]), .ZN(Ufkhu6) );
  INV_X1 U1353 ( .A(n4730), .ZN(n2866) );
  NOR2_X1 U1354 ( .A1(n3623), .A2(n2277), .ZN(n90) );
  OAI21_X1 U1355 ( .B1(n426), .B2(n267), .A(n6474), .ZN(n6473) );
  NAND3_X1 U1356 ( .A1(n417), .A2(n463), .A3(n267), .ZN(n6474) );
  INV_X1 U1357 ( .A(n4729), .ZN(n2852) );
  NOR2_X1 U1358 ( .A1(n397), .A2(n4123), .ZN(n183) );
  NOR2_X1 U1359 ( .A1(n3522), .A2(n875), .ZN(n1918) );
  NAND2_X1 U1360 ( .A1(n878), .A2(n536), .ZN(n1722) );
  AOI21_X1 U1361 ( .B1(n72), .B2(n7375), .A(n1628), .ZN(n1721) );
  NAND2_X1 U1362 ( .A1(n3189), .A2(n82), .ZN(n3724) );
  OAI22_X1 U1363 ( .A1(n6559), .A2(n516), .B1(n3737), .B2(n4658), .ZN(n6558)
         );
  INV_X1 U1364 ( .A(n1519), .ZN(n4658) );
  AOI21_X1 U1365 ( .B1(n4231), .B2(n80), .A(n6561), .ZN(n6559) );
  INV_X1 U1366 ( .A(n542), .ZN(n3190) );
  INV_X1 U1367 ( .A(n236), .ZN(n908) );
  INV_X1 U1368 ( .A(n243), .ZN(n632) );
  INV_X1 U1369 ( .A(n243), .ZN(n635) );
  NOR3_X1 U1370 ( .A1(n508), .A2(n479), .A3(n5564), .ZN(n6040) );
  INV_X1 U1371 ( .A(n4153), .ZN(n2551) );
  INV_X1 U1372 ( .A(n4788), .ZN(n2973) );
  NOR3_X1 U1373 ( .A1(n476), .A2(n2124), .A3(n2694), .ZN(n4317) );
  NOR2_X1 U1374 ( .A1(n4572), .A2(n5047), .ZN(n1594) );
  NOR2_X1 U1375 ( .A1(n3082), .A2(n228), .ZN(n3305) );
  INV_X1 U1376 ( .A(n2184), .ZN(n3141) );
  INV_X1 U1378 ( .A(n5387), .ZN(n3725) );
  NOR2_X1 U1379 ( .A1(n523), .A2(n463), .ZN(n1505) );
  NOR2_X1 U1380 ( .A1(n2856), .A2(n2852), .ZN(n4723) );
  NOR2_X1 U1381 ( .A1(n2694), .A2(n1926), .ZN(n1488) );
  INV_X1 U1382 ( .A(n4446), .ZN(n2745) );
  AOI222_X1 U1383 ( .A1(n415), .A2(n416), .B1(n417), .B2(n418), .C1(n419), 
        .C2(n463), .ZN(n414) );
  OAI21_X1 U1384 ( .B1(n508), .B2(n4265), .A(n426), .ZN(n418) );
  OAI22_X1 U1385 ( .A1(n523), .A2(n4203), .B1(n4688), .B2(n3726), .ZN(n419) );
  NAND2_X1 U1386 ( .A1(n5716), .A2(n5426), .ZN(n4254) );
  OAI221_X1 U1387 ( .B1(n4298), .B2(n3464), .C1(n1454), .C2(n516), .A(n267), 
        .ZN(n5716) );
  NOR4_X1 U1388 ( .A1(n4512), .A2(n4628), .A3(n4685), .A4(n3838), .ZN(n6552)
         );
  OAI22_X1 U1389 ( .A1(n3804), .A2(n4631), .B1(n524), .B2(n3461), .ZN(n2941)
         );
  NOR4_X1 U1390 ( .A1(n3462), .A2(n3463), .A3(n1505), .A4(n3464), .ZN(n3461)
         );
  OAI222_X1 U1391 ( .A1(n463), .A2(n4202), .B1(n538), .B2(n4246), .C1(n4237), 
        .C2(n3858), .ZN(n3462) );
  OAI22_X1 U1392 ( .A1(n7374), .A2(n2755), .B1(n7355), .B2(n3465), .ZN(n3463)
         );
  INV_X1 U1393 ( .A(n2202), .ZN(n2975) );
  NOR2_X1 U1394 ( .A1(n1458), .A2(n479), .ZN(n2875) );
  NOR2_X1 U1395 ( .A1(n2699), .A2(n476), .ZN(n1511) );
  NAND2_X1 U1396 ( .A1(n474), .A2(n508), .ZN(n447) );
  NOR2_X1 U1397 ( .A1(n4512), .A2(n1967), .ZN(n88) );
  NOR4_X1 U1398 ( .A1(n2898), .A2(n3495), .A3(n3496), .A4(n3497), .ZN(n3494)
         );
  NOR4_X1 U1399 ( .A1(n536), .A2(n267), .A3(n529), .A4(n4263), .ZN(n3495) );
  AOI211_X1 U1400 ( .C1(n2243), .C2(n3499), .A(n1967), .B(n270), .ZN(n3496) );
  AOI221_X1 U1401 ( .B1(n2572), .B2(n3498), .C1(n3860), .C2(n692), .A(n7373), 
        .ZN(n3497) );
  AOI221_X1 U1402 ( .B1(n1567), .B2(n1568), .C1(n82), .C2(n1569), .A(n1570), 
        .ZN(n1560) );
  OAI21_X1 U1403 ( .B1(n3831), .B2(n4190), .A(n3833), .ZN(n1569) );
  NOR3_X1 U1404 ( .A1(n1571), .A2(n3714), .A3(n1572), .ZN(n1570) );
  OAI21_X1 U1405 ( .B1(n3550), .B2(n4237), .A(n4263), .ZN(n1568) );
  NAND2_X1 U1406 ( .A1(n493), .A2(n3563), .ZN(n2073) );
  OAI221_X1 U1407 ( .B1(n4246), .B2(n3835), .C1(n3730), .C2(n3804), .A(n4577), 
        .ZN(n2935) );
  NAND4_X1 U1408 ( .A1(n4578), .A2(n2755), .A3(n4265), .A4(n529), .ZN(n4577)
         );
  OAI221_X1 U1409 ( .B1(n517), .B2(n493), .C1(n272), .C2(n3858), .A(n84), .ZN(
        n4578) );
  NOR3_X1 U1410 ( .A1(n503), .A2(n4688), .A3(n1458), .ZN(n3175) );
  NAND3_X1 U1411 ( .A1(n474), .A2(n3550), .A3(n3790), .ZN(n3187) );
  NAND3_X1 U1412 ( .A1(n449), .A2(n523), .A3(n1563), .ZN(n1452) );
  NAND2_X1 U1413 ( .A1(n1539), .A2(n7373), .ZN(n426) );
  NAND3_X1 U1414 ( .A1(n1345), .A2(n1277), .A3(n3439), .ZN(n914) );
  NAND3_X1 U1415 ( .A1(n429), .A2(n2915), .A3(n4106), .ZN(n1436) );
  NOR3_X1 U1416 ( .A1(n516), .A2(n4263), .A3(n4193), .ZN(n4106) );
  NOR4_X1 U1417 ( .A1(n1712), .A2(n1713), .A3(n1714), .A4(n1715), .ZN(n1711)
         );
  NOR3_X1 U1418 ( .A1(n3787), .A2(n1723), .A3(n4738), .ZN(n1712) );
  AOI21_X1 U1419 ( .B1(n2246), .B2(n1720), .A(n3623), .ZN(n1714) );
  NOR2_X1 U1420 ( .A1(n4318), .A2(n464), .ZN(n3181) );
  AOI22_X1 U1421 ( .A1(n1951), .A2(n1902), .B1(n7282), .B2(n483), .ZN(n3222)
         );
  NAND2_X1 U1422 ( .A1(n1856), .A2(n2969), .ZN(n1342) );
  NOR2_X1 U1423 ( .A1(n878), .A2(n7373), .ZN(n1519) );
  NAND2_X1 U1424 ( .A1(n5426), .A2(n2732), .ZN(n4256) );
  NOR2_X1 U1425 ( .A1(n508), .A2(n228), .ZN(n5574) );
  NOR2_X1 U1426 ( .A1(n463), .A2(n517), .ZN(n3464) );
  NOR2_X1 U1427 ( .A1(n2935), .A2(n2936), .ZN(n98) );
  NOR2_X1 U1428 ( .A1(n2394), .A2(n2395), .ZN(n1351) );
  NOR2_X1 U1429 ( .A1(n475), .A2(n4572), .ZN(n1760) );
  NOR2_X1 U1430 ( .A1(n2260), .A2(n475), .ZN(n1586) );
  NOR2_X1 U1431 ( .A1(n2267), .A2(n524), .ZN(n1588) );
  NAND3_X1 U1432 ( .A1(n1672), .A2(n7381), .A3(n473), .ZN(n3271) );
  NOR2_X1 U1433 ( .A1(n463), .A2(n479), .ZN(n5776) );
  NOR2_X1 U1434 ( .A1(n1939), .A2(n476), .ZN(n28) );
  INV_X1 U1435 ( .A(n1587), .ZN(n5037) );
  AOI22_X1 U1436 ( .A1(n2857), .A2(n2477), .B1(n3728), .B2(n3113), .ZN(n1634)
         );
  OAI21_X1 U1437 ( .B1(n3729), .B2(n485), .A(n3715), .ZN(n3728) );
  INV_X1 U1438 ( .A(n518), .ZN(n2243) );
  BUF_X1 U1439 ( .A(n2085), .Z(n815) );
  BUF_X1 U1440 ( .A(n2081), .Z(n836) );
  BUF_X1 U1441 ( .A(n2077), .Z(n855) );
  BUF_X1 U1442 ( .A(n2079), .Z(n848) );
  AOI21_X1 U1443 ( .B1(n1457), .B2(n518), .A(n1704), .ZN(n2498) );
  XNOR2_X1 U1444 ( .A(n2994), .B(n2993), .ZN(n2991) );
  NOR2_X1 U1445 ( .A1(n3238), .A2(n3239), .ZN(n2504) );
  AOI21_X1 U1446 ( .B1(n3238), .B2(n3239), .A(n2504), .ZN(n3237) );
  AOI21_X1 U1447 ( .B1(n1563), .B2(n1975), .A(n1654), .ZN(n1651) );
  NOR3_X1 U1448 ( .A1(n1572), .A2(n272), .A3(n230), .ZN(n1654) );
  NAND4_X1 U1449 ( .A1(n2371), .A2(n2378), .A3(n3251), .A4(n3252), .ZN(n2488)
         );
  NAND3_X1 U1450 ( .A1(n3211), .A2(n473), .A3(n1762), .ZN(n3251) );
  AOI22_X1 U1451 ( .A1(n90), .A2(n4188), .B1(n1462), .B2(n1442), .ZN(n3252) );
  XNOR2_X1 U1452 ( .A(n2991), .B(n3699), .ZN(n3239) );
  INV_X1 U1453 ( .A(n2933), .ZN(n5002) );
  NOR3_X1 U1454 ( .A1(n4246), .A2(n3123), .A3(n529), .ZN(n1746) );
  NOR2_X1 U1455 ( .A1(n2818), .A2(n356), .ZN(n2305) );
  AOI21_X1 U1456 ( .B1(n4240), .B2(n4580), .A(n7374), .ZN(n4576) );
  INV_X1 U1457 ( .A(n3464), .ZN(n4240) );
  OAI21_X1 U1458 ( .B1(n1520), .B2(n228), .A(n4581), .ZN(n4580) );
  NOR3_X1 U1459 ( .A1(n4598), .A2(n4512), .A3(n479), .ZN(n6566) );
  NOR2_X1 U1460 ( .A1(n477), .A2(n7373), .ZN(n2560) );
  OAI22_X1 U1461 ( .A1(n5063), .A2(n2260), .B1(n2256), .B2(n5002), .ZN(n2579)
         );
  INV_X1 U1462 ( .A(n1009), .ZN(n2961) );
  NOR2_X1 U1463 ( .A1(n3831), .A2(n522), .ZN(n4231) );
  OAI22_X1 U1464 ( .A1(n7375), .A2(n2528), .B1(n7374), .B2(n4749), .ZN(n4236)
         );
  NOR2_X1 U1465 ( .A1(n4738), .A2(n502), .ZN(n717) );
  INV_X1 U1466 ( .A(n810), .ZN(n3765) );
  INV_X1 U1467 ( .A(n2194), .ZN(n2985) );
  NOR2_X1 U1468 ( .A1(n4685), .A2(n3123), .ZN(n2899) );
  INV_X1 U1469 ( .A(n2665), .ZN(n3133) );
  NOR2_X1 U1470 ( .A1(n3746), .A2(n463), .ZN(n1653) );
  INV_X1 U1471 ( .A(n3510), .ZN(n1975) );
  INV_X1 U1472 ( .A(n2196), .ZN(n2884) );
  NAND3_X1 U1473 ( .A1(n7375), .A2(n522), .A3(n496), .ZN(n495) );
  NOR2_X1 U1474 ( .A1(n460), .A2(n3742), .ZN(n3038) );
  NOR2_X1 U1475 ( .A1(n460), .A2(n2426), .ZN(n2424) );
  NOR2_X1 U1476 ( .A1(n460), .A2(n2685), .ZN(n2683) );
  NOR2_X1 U1477 ( .A1(n460), .A2(n2800), .ZN(n2798) );
  NOR2_X1 U1478 ( .A1(n3851), .A2(n2536), .ZN(n2534) );
  NOR2_X1 U1479 ( .A1(n460), .A2(n455), .ZN(n2306) );
  NOR2_X1 U1480 ( .A1(n3851), .A2(n4013), .ZN(n2672) );
  NOR2_X1 U1481 ( .A1(n460), .A2(n3862), .ZN(n3859) );
  NOR2_X1 U1482 ( .A1(n3851), .A2(n3579), .ZN(n2245) );
  NOR2_X1 U1483 ( .A1(n460), .A2(n2472), .ZN(n2469) );
  NOR2_X1 U1484 ( .A1(n460), .A2(n3958), .ZN(n3751) );
  OAI211_X1 U1485 ( .C1(n2577), .C2(n476), .A(n1672), .B(n3188), .ZN(n3184) );
  NOR2_X1 U1486 ( .A1(n3851), .A2(n3199), .ZN(n3196) );
  NOR2_X1 U1487 ( .A1(n460), .A2(n3778), .ZN(n3756) );
  NOR2_X1 U1488 ( .A1(n460), .A2(n3558), .ZN(n3555) );
  NOR2_X1 U1489 ( .A1(n3851), .A2(n4843), .ZN(n3927) );
  INV_X1 U1490 ( .A(n1835), .ZN(n2477) );
  NOR2_X1 U1491 ( .A1(n3851), .A2(n2526), .ZN(n2523) );
  NOR2_X1 U1492 ( .A1(n3851), .A2(n4121), .ZN(n4021) );
  INV_X1 U1493 ( .A(n1345), .ZN(n4324) );
  NOR2_X1 U1494 ( .A1(n3851), .A2(n4276), .ZN(n3665) );
  NOR2_X1 U1495 ( .A1(n3851), .A2(n3639), .ZN(n3090) );
  NOR2_X1 U1496 ( .A1(n460), .A2(n3677), .ZN(n3157) );
  NOR2_X1 U1497 ( .A1(n3851), .A2(n3644), .ZN(n2259) );
  NOR2_X1 U1498 ( .A1(n3851), .A2(n2824), .ZN(n2821) );
  NOR2_X1 U1499 ( .A1(n3851), .A2(n3612), .ZN(n2223) );
  NOR2_X1 U1500 ( .A1(n3851), .A2(n3542), .ZN(n3539) );
  NOR2_X1 U1501 ( .A1(n3851), .A2(n3597), .ZN(n2968) );
  NOR2_X1 U1502 ( .A1(n460), .A2(n4039), .ZN(n3627) );
  NOR2_X1 U1503 ( .A1(n3851), .A2(n3624), .ZN(n2463) );
  NOR2_X1 U1504 ( .A1(n3851), .A2(n3649), .ZN(n3487) );
  NOR2_X1 U1505 ( .A1(n3851), .A2(n4472), .ZN(n3613) );
  NAND2_X1 U1506 ( .A1(n3211), .A2(n3250), .ZN(n2492) );
  OAI21_X1 U1507 ( .B1(n475), .B2(n2694), .A(n2256), .ZN(n3250) );
  AOI22_X1 U1508 ( .A1(n3697), .A2(n2503), .B1(n2504), .B2(n2505), .ZN(n2491)
         );
  NAND3_X1 U1509 ( .A1(n4559), .A2(n3082), .A3(n4561), .ZN(n4536) );
  INV_X1 U1510 ( .A(n2198), .ZN(n2978) );
  NAND4_X1 U1511 ( .A1(n2911), .A2(n2912), .A3(n2913), .A4(n2914), .ZN(n2910)
         );
  AOI22_X1 U1512 ( .A1(n513), .A2(n693), .B1(n1761), .B2(n2915), .ZN(n2914) );
  NAND3_X1 U1513 ( .A1(n1672), .A2(n476), .A3(n2916), .ZN(n2913) );
  INV_X1 U1514 ( .A(n4439), .ZN(n2715) );
  INV_X1 U1515 ( .A(n2193), .ZN(n2882) );
  OAI21_X1 U1516 ( .B1(n1586), .B2(n518), .A(n28), .ZN(n1935) );
  NAND2_X1 U1517 ( .A1(n3511), .A2(n485), .ZN(n2067) );
  INV_X1 U1518 ( .A(n2053), .ZN(n3144) );
  NAND2_X1 U1519 ( .A1(n913), .A2(n3156), .ZN(n537) );
  INV_X1 U1520 ( .A(n1762), .ZN(n4186) );
  INV_X1 U1521 ( .A(n2200), .ZN(n2886) );
  INV_X1 U1522 ( .A(n700), .ZN(n3258) );
  INV_X1 U1523 ( .A(n1512), .ZN(n1939) );
  NOR2_X1 U1524 ( .A1(n3550), .A2(n503), .ZN(n1625) );
  INV_X1 U1525 ( .A(n2199), .ZN(n2988) );
  INV_X1 U1526 ( .A(n1284), .ZN(n4306) );
  NAND2_X1 U1527 ( .A1(n3170), .A2(n1571), .ZN(n3183) );
  AND2_X1 U1528 ( .A1(n5544), .A2(n1856), .ZN(n3582) );
  INV_X1 U1529 ( .A(n2704), .ZN(n3200) );
  INV_X1 U1530 ( .A(n3049), .ZN(n3066) );
  INV_X1 U1531 ( .A(n4342), .ZN(n2702) );
  INV_X1 U1532 ( .A(n1683), .ZN(n4555) );
  AND3_X1 U1533 ( .A1(n2378), .A2(n3209), .A3(n3210), .ZN(n3097) );
  AOI22_X1 U1534 ( .A1(n2916), .A2(n3211), .B1(n1462), .B2(n230), .ZN(n3210)
         );
  INV_X1 U1535 ( .A(n455), .ZN(n3952) );
  NAND2_X1 U1536 ( .A1(n3582), .A2(n3010), .ZN(n3541) );
  INV_X1 U1537 ( .A(n905), .ZN(n3010) );
  INV_X1 U1538 ( .A(n1894), .ZN(n2998) );
  NAND3_X1 U1539 ( .A1(n2911), .A2(n4756), .A3(n3265), .ZN(n3264) );
  NAND3_X1 U1540 ( .A1(n473), .A2(n7381), .A3(n1456), .ZN(n3265) );
  INV_X1 U1541 ( .A(n3188), .ZN(n2250) );
  INV_X1 U1542 ( .A(n3321), .ZN(n2388) );
  INV_X1 U1543 ( .A(n3366), .ZN(n2368) );
  NAND3_X1 U1544 ( .A1(n6563), .A2(n3740), .A3(n6565), .ZN(n6556) );
  AOI21_X1 U1545 ( .B1(n5776), .B2(n516), .A(n6566), .ZN(n6565) );
  INV_X1 U1546 ( .A(n3170), .ZN(n3740) );
  NAND3_X1 U1547 ( .A1(n87), .A2(n523), .A3(n4092), .ZN(n6563) );
  NAND2_X1 U1548 ( .A1(n3236), .A2(n3237), .ZN(n3001) );
  INV_X1 U1549 ( .A(n2046), .ZN(n3142) );
  AND2_X1 U1550 ( .A1(n5668), .A2(n2969), .ZN(n4781) );
  INV_X1 U1551 ( .A(n2842), .ZN(n2244) );
  INV_X1 U1552 ( .A(n70), .ZN(n1934) );
  INV_X1 U1553 ( .A(n3363), .ZN(n2396) );
  INV_X1 U1554 ( .A(n4835), .ZN(n3981) );
  INV_X1 U1555 ( .A(n530), .ZN(n3158) );
  INV_X1 U1556 ( .A(n3372), .ZN(n2358) );
  INV_X1 U1557 ( .A(n57), .ZN(n3556) );
  INV_X1 U1558 ( .A(n4243), .ZN(n4668) );
  NAND2_X1 U1559 ( .A1(n7355), .A2(n57), .ZN(n4230) );
  INV_X1 U1560 ( .A(Idfpw6[31]), .ZN(n2281) );
  INV_X1 U1561 ( .A(n4309), .ZN(n2122) );
  OAI221_X1 U1562 ( .B1(n2607), .B2(n4310), .C1(n2608), .C2(n3173), .A(n3183), 
        .ZN(n4309) );
  NAND2_X1 U1563 ( .A1(n228), .A2(n7373), .ZN(n4310) );
  AND4_X1 U1564 ( .A1(n4756), .A2(n1452), .A3(n3186), .A4(n3187), .ZN(n3185)
         );
  INV_X1 U1565 ( .A(n1638), .ZN(n2857) );
  INV_X1 U1566 ( .A(n2586), .ZN(n3701) );
  OAI21_X1 U1567 ( .B1(n4572), .B2(n1739), .A(n79), .ZN(n2586) );
  OAI221_X1 U1568 ( .B1(n7514), .B2(n3271), .C1(n4749), .C2(n426), .A(n2126), 
        .ZN(n3255) );
  INV_X1 U1569 ( .A(n3273), .ZN(n2126) );
  OAI221_X1 U1570 ( .B1(n1470), .B2(n2608), .C1(n3275), .C2(n3684), .A(n2912), 
        .ZN(n3273) );
  OR2_X1 U1571 ( .A1(n449), .A2(n3186), .ZN(n3275) );
  INV_X1 U1572 ( .A(n2738), .ZN(n3630) );
  INV_X1 U1573 ( .A(n4304), .ZN(n1910) );
  BUF_X1 U1574 ( .A(n2155), .Z(n788) );
  INV_X1 U1575 ( .A(n244), .ZN(n913) );
  INV_X1 U1576 ( .A(n244), .ZN(n917) );
  INV_X1 U1577 ( .A(n247), .ZN(n847) );
  INV_X1 U1578 ( .A(n247), .ZN(n841) );
  INV_X1 U1579 ( .A(n249), .ZN(n833) );
  INV_X1 U1580 ( .A(n249), .ZN(n830) );
  INV_X1 U1581 ( .A(n250), .ZN(n863) );
  INV_X1 U1582 ( .A(n253), .ZN(n854) );
  INV_X1 U1583 ( .A(n253), .ZN(n850) );
  INV_X1 U1584 ( .A(n250), .ZN(n857) );
  NAND4_X1 U1585 ( .A1(n1455), .A2(n477), .A3(n4263), .A4(n265), .ZN(n2912) );
  NOR3_X1 U1586 ( .A1(n516), .A2(n502), .A3(n1458), .ZN(n1475) );
  NOR4_X1 U1587 ( .A1(n524), .A2(n7514), .A3(n3625), .A4(n4186), .ZN(n2763) );
  OAI21_X1 U1588 ( .B1(n1685), .B2(n470), .A(n2454), .ZN(n2412) );
  BUF_X1 U1589 ( .A(n703), .Z(n891) );
  NOR2_X1 U1590 ( .A1(n2267), .A2(n2699), .ZN(n1737) );
  NAND4_X1 U1591 ( .A1(n1748), .A2(n502), .A3(n1462), .A4(n4242), .ZN(n2907)
         );
  NOR2_X1 U1592 ( .A1(n4189), .A2(n4668), .ZN(n4242) );
  NOR2_X1 U1593 ( .A1(n470), .A2(n270), .ZN(n2577) );
  NAND2_X1 U1594 ( .A1(n693), .A2(n485), .ZN(n1470) );
  BUF_X1 U1595 ( .A(n2087), .Z(n803) );
  NAND3_X1 U1596 ( .A1(n3561), .A2(n523), .A3(n3562), .ZN(n1959) );
  NOR3_X1 U1597 ( .A1(n2594), .A2(n416), .A3(n479), .ZN(n3502) );
  INV_X1 U1598 ( .A(n988), .ZN(n3476) );
  NOR3_X1 U1599 ( .A1(n1503), .A2(n1504), .A3(n1505), .ZN(n1502) );
  OAI22_X1 U1600 ( .A1(n4265), .A2(n3788), .B1(n4195), .B2(n3709), .ZN(n1503)
         );
  NOR3_X1 U1601 ( .A1(n3768), .A2(n486), .A3(n4237), .ZN(n1912) );
  NAND3_X1 U1602 ( .A1(n80), .A2(n81), .A3(n82), .ZN(n68) );
  NAND4_X1 U1603 ( .A1(n3787), .A2(n266), .A3(n84), .A4(n85), .ZN(n81) );
  AOI22_X1 U1604 ( .A1(n536), .A2(n1975), .B1(n87), .B2(n485), .ZN(n85) );
  NAND3_X1 U1605 ( .A1(n479), .A2(n485), .A3(n493), .ZN(n2746) );
  NOR2_X1 U1606 ( .A1(n476), .A2(n225), .ZN(n2767) );
  INV_X1 U1607 ( .A(n609), .ZN(n3202) );
  INV_X1 U1608 ( .A(n990), .ZN(n3474) );
  NAND2_X1 U1609 ( .A1(n1763), .A2(n2753), .ZN(n2750) );
  OAI211_X1 U1610 ( .C1(n3123), .C2(n2754), .A(n3727), .B(n2755), .ZN(n2753)
         );
  AOI21_X1 U1611 ( .B1(n1519), .B2(n536), .A(n1536), .ZN(n1535) );
  NOR3_X1 U1612 ( .A1(n4188), .A2(n3628), .A3(n4195), .ZN(n1536) );
  NAND2_X1 U1613 ( .A1(n1685), .A2(n475), .ZN(n444) );
  NAND4_X1 U1614 ( .A1(n2877), .A2(n3122), .A3(n2878), .A4(n2879), .ZN(n2871)
         );
  NAND3_X1 U1615 ( .A1(n474), .A2(n492), .A3(n429), .ZN(n2878) );
  NAND3_X1 U1616 ( .A1(n237), .A2(n536), .A3(n1615), .ZN(n2877) );
  AOI22_X1 U1617 ( .A1(n2880), .A2(n2881), .B1(n1505), .B2(n1938), .ZN(n2879)
         );
  BUF_X1 U1618 ( .A(n2083), .Z(n828) );
  INV_X1 U1619 ( .A(n1004), .ZN(n3475) );
  AOI21_X1 U1620 ( .B1(n2739), .B2(n1620), .A(n1462), .ZN(n2737) );
  NOR2_X1 U1621 ( .A1(n485), .A2(n2572), .ZN(n2739) );
  OAI21_X1 U1622 ( .B1(n470), .B2(n4188), .A(n90), .ZN(n3098) );
  NAND3_X1 U1623 ( .A1(n88), .A2(n89), .A3(n90), .ZN(n66) );
  OAI22_X1 U1624 ( .A1(n4566), .A2(n4725), .B1(n4572), .B2(n93), .ZN(n89) );
  OAI21_X1 U1625 ( .B1(n1474), .B2(n1475), .A(n230), .ZN(n1473) );
  NOR3_X1 U1626 ( .A1(n2607), .A2(n485), .A3(n508), .ZN(n1474) );
  OAI21_X1 U1627 ( .B1(n427), .B2(n428), .A(n429), .ZN(n413) );
  NOR3_X1 U1628 ( .A1(n4642), .A2(n4237), .A3(n479), .ZN(n427) );
  NOR2_X1 U1629 ( .A1(n270), .A2(n4672), .ZN(n1941) );
  AND2_X1 U1630 ( .A1(n1854), .A2(n1856), .ZN(n389) );
  NOR2_X1 U1631 ( .A1(n5063), .A2(n4564), .ZN(n2589) );
  NAND3_X1 U1632 ( .A1(n476), .A2(n529), .A3(n7514), .ZN(n3499) );
  INV_X1 U1633 ( .A(n2123), .ZN(n2967) );
  NAND2_X1 U1634 ( .A1(n2699), .A2(n2277), .ZN(n2454) );
  INV_X1 U1635 ( .A(n2434), .ZN(n3904) );
  INV_X1 U1636 ( .A(n591), .ZN(n3204) );
  INV_X1 U1637 ( .A(n1073), .ZN(n3480) );
  NOR2_X1 U1638 ( .A1(n529), .A2(n523), .ZN(n1564) );
  INV_X1 U1639 ( .A(n999), .ZN(n2136) );
  NAND2_X1 U1640 ( .A1(n4330), .A2(n4301), .ZN(n1275) );
  INV_X1 U1641 ( .A(n1701), .ZN(n2258) );
  INV_X1 U1642 ( .A(n657), .ZN(n3219) );
  INV_X1 U1643 ( .A(n1272), .ZN(n3441) );
  OR3_X1 U1644 ( .A1(n878), .A2(n270), .A3(n2381), .ZN(n4321) );
  INV_X1 U1645 ( .A(n639), .ZN(n3192) );
  NAND2_X1 U1646 ( .A1(n2107), .A2(n1986), .ZN(n3887) );
  OAI211_X1 U1647 ( .C1(\eq_3147/A[26] ), .C2(n3848), .A(n1805), .B(n3889), 
        .ZN(n3888) );
  INV_X1 U1648 ( .A(n2153), .ZN(n1530) );
  INV_X1 U1649 ( .A(HADDR[29]), .ZN(n1553) );
  OAI21_X1 U1650 ( .B1(n5756), .B2(n5757), .A(n2731), .ZN(n4259) );
  OAI222_X1 U1651 ( .A1(n7355), .A2(n4631), .B1(n4232), .B2(n3830), .C1(n4193), 
        .C2(n3800), .ZN(n5757) );
  OAI221_X1 U1652 ( .B1(n228), .B2(n3804), .C1(n228), .C2(n5758), .A(n5759), 
        .ZN(n5756) );
  AOI22_X1 U1653 ( .A1(n2071), .A2(n516), .B1(n1454), .B2(n1463), .ZN(n5758)
         );
  OAI221_X1 U1654 ( .B1(n1590), .B2(n661), .C1(n2324), .C2(n3900), .A(n3909), 
        .ZN(\eq_3147/A[25] ) );
  NAND2_X1 U1655 ( .A1(N5fpw6[26]), .A2(n669), .ZN(n3909) );
  INV_X1 U1656 ( .A(n435), .ZN(n4265) );
  OR2_X1 U1657 ( .A1(HADDR[29]), .A2(HADDR[30]), .ZN(HPROT[2]) );
  OAI221_X1 U1658 ( .B1(n3802), .B2(n664), .C1(n1581), .C2(n661), .A(n3963), 
        .ZN(\eq_3147/A[26] ) );
  NAND2_X1 U1659 ( .A1(N5fpw6[27]), .A2(n667), .ZN(n3963) );
  NOR4_X1 U1660 ( .A1(n5304), .A2(n2466), .A3(n5307), .A4(n5302), .ZN(n6004)
         );
  OAI221_X1 U1661 ( .B1(n3801), .B2(n664), .C1(n1575), .C2(n661), .A(n4026), 
        .ZN(n201) );
  NAND2_X1 U1662 ( .A1(N5fpw6[28]), .A2(n667), .ZN(n4026) );
  OAI221_X1 U1663 ( .B1(n3798), .B2(n3900), .C1(n1551), .C2(n661), .A(n3906), 
        .ZN(n200) );
  NAND2_X1 U1664 ( .A1(N5fpw6[29]), .A2(n669), .ZN(n3906) );
  BUF_X1 U1665 ( .A(n6007), .Z(n540) );
  OAI21_X1 U1666 ( .B1(n5748), .B2(n5749), .A(n2731), .ZN(n4452) );
  OAI22_X1 U1667 ( .A1(n5750), .A2(n4229), .B1(n4265), .B2(n5751), .ZN(n5749)
         );
  NAND2_X1 U1668 ( .A1(n4298), .A2(n228), .ZN(n5751) );
  NAND2_X1 U1669 ( .A1(n5722), .A2(n5728), .ZN(n4291) );
  INV_X1 U1670 ( .A(n4424), .ZN(n2757) );
  NAND3_X1 U1671 ( .A1(n1462), .A2(n2731), .A3(n3561), .ZN(n4451) );
  NAND2_X1 U1672 ( .A1(n5724), .A2(n5728), .ZN(n4288) );
  BUF_X1 U1673 ( .A(n4873), .Z(n575) );
  NAND2_X1 U1674 ( .A1(n5722), .A2(n5723), .ZN(n4503) );
  OAI222_X1 U1675 ( .A1(n627), .A2(n3774), .B1(n625), .B2(n5928), .C1(n623), 
        .C2(n6260), .ZN(n4992) );
  OAI222_X1 U1676 ( .A1(n4858), .A2(n4272), .B1(n4859), .B2(n5976), .C1(n623), 
        .C2(n6249), .ZN(n4977) );
  BUF_X1 U1677 ( .A(n4876), .Z(n569) );
  BUF_X1 U1678 ( .A(n4870), .Z(n578) );
  BUF_X1 U1679 ( .A(n4263), .Z(n463) );
  NOR2_X1 U1680 ( .A1(n5313), .A2(n5312), .ZN(n5910) );
  AOI22_X1 U1681 ( .A1(n200), .A2(n1573), .B1(n201), .B2(n199), .ZN(n2153) );
  BUF_X1 U1682 ( .A(n4859), .Z(n625) );
  BUF_X1 U1683 ( .A(n6001), .Z(n564) );
  BUF_X1 U1684 ( .A(n6006), .Z(n541) );
  BUF_X1 U1685 ( .A(n6002), .Z(n563) );
  BUF_X1 U1686 ( .A(n6003), .Z(n561) );
  OAI21_X1 U1687 ( .B1(n474), .B2(n435), .A(n505), .ZN(n5734) );
  NOR2_X1 U1688 ( .A1(n3789), .A2(n3822), .ZN(Idfpw6[0]) );
  OAI22_X1 U1689 ( .A1(n5018), .A2(n8088), .B1(n623), .B2(n6176), .ZN(n5909)
         );
  OAI22_X1 U1690 ( .A1(n5018), .A2(n8078), .B1(n623), .B2(n6219), .ZN(n5017)
         );
  OAI22_X1 U1691 ( .A1(n572), .A2(n7800), .B1(n569), .B2(n5484), .ZN(n6513) );
  OAI22_X1 U1692 ( .A1(n572), .A2(n7748), .B1(n569), .B2(n5506), .ZN(n6451) );
  OAI22_X1 U1693 ( .A1(n572), .A2(n7760), .B1(n569), .B2(n5468), .ZN(n6519) );
  OAI22_X1 U1694 ( .A1(n572), .A2(n7809), .B1(n569), .B2(n5562), .ZN(n6491) );
  NAND3_X1 U1695 ( .A1(n200), .A2(n201), .A3(n199), .ZN(n3848) );
  OAI22_X1 U1696 ( .A1(n8127), .A2(n646), .B1(n8055), .B2(n4291), .ZN(n4391)
         );
  NAND3_X1 U1697 ( .A1(n5769), .A2(n4394), .A3(n5770), .ZN(n4858) );
  INV_X1 U1698 ( .A(n4821), .ZN(n3773) );
  OAI22_X1 U1699 ( .A1(n5730), .A2(n564), .B1(n6628), .B2(n563), .ZN(n6014) );
  OAI22_X1 U1700 ( .A1(n5673), .A2(n564), .B1(n6686), .B2(n563), .ZN(n6000) );
  OAI22_X1 U1701 ( .A1(n5642), .A2(n564), .B1(n6642), .B2(n563), .ZN(n6018) );
  NAND3_X1 U1702 ( .A1(n5304), .A2(n5302), .A3(n5722), .ZN(n4176) );
  INV_X1 U1703 ( .A(n199), .ZN(n1529) );
  NAND2_X1 U1704 ( .A1(n5770), .A2(n5911), .ZN(n5018) );
  NAND2_X1 U1705 ( .A1(n5741), .A2(n2731), .ZN(n4258) );
  OAI211_X1 U1706 ( .C1(n4232), .C2(n4244), .A(n4127), .B(n5742), .ZN(n5741)
         );
  AOI21_X1 U1707 ( .B1(n7282), .B2(n5743), .A(n5744), .ZN(n5742) );
  OAI21_X1 U1708 ( .B1(n4263), .B2(n4611), .A(n3805), .ZN(n5743) );
  INV_X1 U1709 ( .A(n4386), .ZN(Qbfpw6_0) );
  NAND2_X1 U1710 ( .A1(n5770), .A2(n5910), .ZN(n4860) );
  INV_X1 U1711 ( .A(n5492), .ZN(n2462) );
  INV_X1 U1712 ( .A(n4502), .ZN(n2336) );
  BUF_X1 U1713 ( .A(n529), .Z(n526) );
  INV_X1 U1714 ( .A(n4833), .ZN(n2546) );
  NAND2_X1 U1715 ( .A1(n5913), .A2(n6517), .ZN(n4875) );
  INV_X1 U1716 ( .A(n4255), .ZN(Qbfpw6_1) );
  NOR2_X1 U1717 ( .A1(n671), .A2(n3811), .ZN(Idfpw6[1]) );
  INV_X1 U1718 ( .A(n4824), .ZN(Qbfpw6_3) );
  NOR2_X1 U1719 ( .A1(n3789), .A2(n3796), .ZN(Idfpw6[3]) );
  INV_X1 U1720 ( .A(n5715), .ZN(Qbfpw6_4) );
  NOR2_X1 U1721 ( .A1(n3789), .A2(n3795), .ZN(Idfpw6[4]) );
  INV_X1 U1722 ( .A(n5094), .ZN(Qbfpw6_5) );
  NOR2_X1 U1723 ( .A1(n3789), .A2(n3794), .ZN(Idfpw6[5]) );
  NOR2_X1 U1724 ( .A1(n3789), .A2(n3793), .ZN(Idfpw6[6]) );
  INV_X1 U1725 ( .A(n4511), .ZN(E2epw6) );
  NOR2_X1 U1726 ( .A1(n3789), .A2(n3792), .ZN(Idfpw6[7]) );
  NOR2_X1 U1727 ( .A1(n3789), .A2(n3791), .ZN(Idfpw6[8]) );
  NOR2_X1 U1728 ( .A1(n671), .A2(n2326), .ZN(Idfpw6[9]) );
  INV_X1 U1729 ( .A(n4741), .ZN(Qbfpw6_10) );
  NOR2_X1 U1730 ( .A1(n671), .A2(n3821), .ZN(Idfpw6[10]) );
  NOR2_X1 U1731 ( .A1(n671), .A2(n3820), .ZN(Idfpw6[11]) );
  NOR2_X1 U1732 ( .A1(n671), .A2(n3819), .ZN(Idfpw6[12]) );
  NOR2_X1 U1733 ( .A1(n671), .A2(n3818), .ZN(Idfpw6[13]) );
  NOR2_X1 U1734 ( .A1(n3789), .A2(n3817), .ZN(Idfpw6[14]) );
  INV_X1 U1735 ( .A(n4480), .ZN(L2epw6) );
  NOR2_X1 U1736 ( .A1(n3789), .A2(n3816), .ZN(Idfpw6[15]) );
  INV_X1 U1737 ( .A(n5072), .ZN(Z2epw6) );
  NOR2_X1 U1738 ( .A1(n3789), .A2(n3815), .ZN(Idfpw6[16]) );
  NOR2_X1 U1739 ( .A1(n671), .A2(n3814), .ZN(Idfpw6[17]) );
  INV_X1 U1740 ( .A(n4422), .ZN(N3epw6) );
  NOR2_X1 U1741 ( .A1(n671), .A2(n3813), .ZN(Idfpw6[18]) );
  INV_X1 U1742 ( .A(n5608), .ZN(U3epw6) );
  NOR2_X1 U1743 ( .A1(n671), .A2(n3812), .ZN(Idfpw6[19]) );
  INV_X1 U1744 ( .A(n4660), .ZN(B4epw6) );
  NOR2_X1 U1745 ( .A1(n671), .A2(n3810), .ZN(Idfpw6[20]) );
  INV_X1 U1746 ( .A(n4600), .ZN(I4epw6) );
  NOR2_X1 U1747 ( .A1(n671), .A2(n3809), .ZN(Idfpw6[21]) );
  NOR2_X1 U1748 ( .A1(n671), .A2(n3808), .ZN(Idfpw6[22]) );
  INV_X1 U1749 ( .A(n4162), .ZN(Qbfpw6[23]) );
  NOR2_X1 U1750 ( .A1(n671), .A2(n3807), .ZN(Idfpw6[23]) );
  NOR2_X1 U1751 ( .A1(n671), .A2(n3806), .ZN(Idfpw6[24]) );
  NOR2_X1 U1752 ( .A1(n3789), .A2(n3802), .ZN(Idfpw6[28]) );
  NOR2_X1 U1753 ( .A1(n3789), .A2(n3801), .ZN(Idfpw6[29]) );
  NOR2_X1 U1754 ( .A1(n3789), .A2(n3798), .ZN(Idfpw6[30]) );
  AND2_X1 U1755 ( .A1(n2546), .A2(n4627), .ZN(n4260) );
  NAND3_X1 U1756 ( .A1(n508), .A2(n2731), .A3(n3562), .ZN(n4627) );
  INV_X1 U1757 ( .A(n5281), .ZN(n2458) );
  BUF_X1 U1758 ( .A(n7374), .Z(n492) );
  AND2_X1 U1759 ( .A1(n5770), .A2(n5913), .ZN(n4864) );
  AND2_X1 U1760 ( .A1(n5769), .A2(n6517), .ZN(n4867) );
  AND2_X1 U1761 ( .A1(n5911), .A2(n6517), .ZN(n4872) );
  AND2_X1 U1762 ( .A1(n5910), .A2(n6517), .ZN(n4868) );
  AND2_X1 U1763 ( .A1(n5912), .A2(n5769), .ZN(n4863) );
  AND2_X1 U1764 ( .A1(n6523), .A2(n2466), .ZN(n5999) );
  AND2_X1 U1765 ( .A1(n5912), .A2(n5911), .ZN(n4861) );
  AND2_X1 U1766 ( .A1(n5912), .A2(n5913), .ZN(n4862) );
  AND2_X1 U1767 ( .A1(n5912), .A2(n5910), .ZN(n4856) );
  INV_X1 U1768 ( .A(n2709), .ZN(n2330) );
  AND4_X1 U1769 ( .A1(n3823), .A2(n3824), .A3(n3825), .A4(n3826), .ZN(n3789)
         );
  NAND3_X1 U1770 ( .A1(n82), .A2(n272), .A3(n1454), .ZN(n3824) );
  OAI21_X1 U1771 ( .B1(n435), .B2(n3790), .A(n477), .ZN(n3823) );
  AOI221_X1 U1772 ( .B1(n1902), .B2(n7282), .C1(n3561), .C2(n265), .A(n3829), 
        .ZN(n3825) );
  INV_X1 U1773 ( .A(n5724), .ZN(n2470) );
  INV_X1 U1774 ( .A(n5019), .ZN(n4351) );
  OAI21_X1 U1775 ( .B1(n3831), .B2(n4633), .A(n5922), .ZN(n354) );
  NAND3_X1 U1776 ( .A1(n1663), .A2(n522), .A3(n2562), .ZN(n5922) );
  OAI221_X1 U1777 ( .B1(n3810), .B2(n3900), .C1(n1637), .C2(n3901), .A(n3914), 
        .ZN(\eq_3147/A[18] ) );
  NAND2_X1 U1778 ( .A1(N5fpw6[19]), .A2(n667), .ZN(n3914) );
  INV_X1 U1779 ( .A(Nxkbx6[21]), .ZN(n1637) );
  OAI221_X1 U1780 ( .B1(n2328), .B2(n664), .C1(n1597), .C2(n661), .A(n3945), 
        .ZN(\eq_3147/A[24] ) );
  NAND2_X1 U1781 ( .A1(N5fpw6[25]), .A2(n667), .ZN(n3945) );
  OAI221_X1 U1782 ( .B1(n3809), .B2(n664), .C1(n1632), .C2(n3901), .A(n3976), 
        .ZN(\eq_3147/A[19] ) );
  NAND2_X1 U1783 ( .A1(N5fpw6[20]), .A2(n667), .ZN(n3976) );
  INV_X1 U1784 ( .A(Nxkbx6[22]), .ZN(n1632) );
  OAI221_X1 U1785 ( .B1(n3808), .B2(n3900), .C1(n1618), .C2(n661), .A(n5064), 
        .ZN(\eq_3147/A[20] ) );
  NAND2_X1 U1786 ( .A1(N5fpw6[21]), .A2(n667), .ZN(n5064) );
  INV_X1 U1787 ( .A(Nxkbx6[23]), .ZN(n1618) );
  NOR3_X2 U1788 ( .A1(n5304), .A2(n5302), .A3(n2470), .ZN(n4290) );
  OAI221_X1 U1789 ( .B1(n3807), .B2(n3900), .C1(n1614), .C2(n3901), .A(n3912), 
        .ZN(\eq_3147/A[21] ) );
  NAND2_X1 U1790 ( .A1(N5fpw6[22]), .A2(n667), .ZN(n3912) );
  OAI221_X1 U1791 ( .B1(n1657), .B2(n661), .C1(n3814), .C2(n3900), .A(n5625), 
        .ZN(\eq_3147/A[15] ) );
  NAND2_X1 U1792 ( .A1(N5fpw6[16]), .A2(n667), .ZN(n5625) );
  INV_X1 U1793 ( .A(Nxkbx6[18]), .ZN(n1657) );
  OAI221_X1 U1794 ( .B1(n2334), .B2(n3900), .C1(n1604), .C2(n661), .A(n3910), 
        .ZN(\eq_3147/A[23] ) );
  NAND2_X1 U1795 ( .A1(N5fpw6[24]), .A2(n667), .ZN(n3910) );
  OAI221_X1 U1796 ( .B1(n3816), .B2(n664), .C1(n1692), .C2(n3901), .A(n3917), 
        .ZN(\eq_3147/A[13] ) );
  NAND2_X1 U1797 ( .A1(N5fpw6[14]), .A2(n667), .ZN(n3917) );
  NOR2_X1 U1798 ( .A1(n2611), .A2(n2612), .ZN(Tgfpw6[9]) );
  AOI221_X1 U1799 ( .B1(n4424), .B2(n4637), .C1(n2730), .C2(n4425), .A(n4426), 
        .ZN(n4423) );
  AOI221_X1 U1800 ( .B1(n4424), .B2(n5070), .C1(n2730), .C2(n4471), .A(n4426), 
        .ZN(n4481) );
  AOI221_X1 U1801 ( .B1(n4424), .B2(n5074), .C1(n2730), .C2(n4909), .A(n4426), 
        .ZN(n5073) );
  NOR2_X1 U1802 ( .A1(n2611), .A2(n2641), .ZN(Tgfpw6[11]) );
  OAI221_X1 U1803 ( .B1(n3806), .B2(n664), .C1(n1608), .C2(n661), .A(n4051), 
        .ZN(\eq_3147/A[22] ) );
  NAND2_X1 U1804 ( .A1(N5fpw6[23]), .A2(n667), .ZN(n4051) );
  NOR4_X1 U1805 ( .A1(Affpw6[29]), .A2(n635), .A3(n4803), .A4(n4804), .ZN(
        n3420) );
  OAI21_X1 U1806 ( .B1(n2538), .B2(n4808), .A(n4809), .ZN(n4803) );
  OAI222_X1 U1807 ( .A1(n2729), .A2(n2702), .B1(n3032), .B2(n4153), .C1(n439), 
        .C2(n1575), .ZN(n4804) );
  AOI22_X1 U1808 ( .A1(n2293), .A2(n4254), .B1(n4253), .B2(n3801), .ZN(n4808)
         );
  NOR2_X1 U1809 ( .A1(n2611), .A2(n2640), .ZN(Tgfpw6[12]) );
  NOR2_X1 U1810 ( .A1(n678), .A2(n2639), .ZN(Tgfpw6[13]) );
  BUF_X1 U1811 ( .A(n4871), .Z(n577) );
  NOR2_X1 U1812 ( .A1(n679), .A2(n2638), .ZN(Tgfpw6[14]) );
  NOR2_X1 U1813 ( .A1(n678), .A2(n2637), .ZN(Tgfpw6[15]) );
  OAI211_X1 U1814 ( .C1(n2926), .C2(n2927), .A(n2928), .B(n2929), .ZN(n2925)
         );
  NOR2_X1 U1815 ( .A1(n2933), .A2(n1752), .ZN(n2926) );
  OAI221_X1 U1816 ( .B1(n1752), .B2(n472), .C1(n2507), .C2(n1523), .A(n2945), 
        .ZN(n2928) );
  NAND4_X1 U1817 ( .A1(n3433), .A2(n3434), .A3(n3435), .A4(n3436), .ZN(n3384)
         );
  NOR3_X1 U1818 ( .A1(n3440), .A2(n2298), .A3(n3442), .ZN(n3435) );
  NOR4_X1 U1819 ( .A1(n3437), .A2(Affpw6[2]), .A3(Affpw6[5]), .A4(Affpw6[4]), 
        .ZN(n3436) );
  OR3_X1 U1820 ( .A1(n3438), .A2(Affpw6[28]), .A3(n2301), .ZN(n3437) );
  NOR2_X1 U1821 ( .A1(n678), .A2(n2635), .ZN(Tgfpw6[17]) );
  OAI221_X1 U1822 ( .B1(n3602), .B2(n4153), .C1(n4154), .C2(n1590), .A(n5690), 
        .ZN(n3413) );
  AOI211_X1 U1823 ( .C1(n5691), .C2(Qbfpw6[27]), .A(Affpw6[27]), .B(n5692), 
        .ZN(n5690) );
  OAI22_X1 U1824 ( .A1(n2550), .A2(n2324), .B1(n4446), .B2(n5695), .ZN(n5691)
         );
  NOR3_X1 U1825 ( .A1(n2324), .A2(Qbfpw6[27]), .A3(n2549), .ZN(n5692) );
  NOR2_X1 U1826 ( .A1(n679), .A2(n2634), .ZN(Tgfpw6[18]) );
  XNOR2_X1 U1827 ( .A(n2545), .B(n5589), .ZN(C1epw6) );
  AOI221_X1 U1828 ( .B1(n4424), .B2(n470), .C1(n2730), .C2(n4938), .A(n4426), 
        .ZN(n5589) );
  XNOR2_X1 U1829 ( .A(n2545), .B(n5139), .ZN(X1epw6) );
  AOI221_X1 U1830 ( .B1(n4424), .B2(n5299), .C1(n2730), .C2(n4888), .A(n4426), 
        .ZN(n5139) );
  XNOR2_X1 U1831 ( .A(n2545), .B(n5357), .ZN(Q1epw6) );
  AOI221_X1 U1832 ( .B1(n4424), .B2(n3083), .C1(n2730), .C2(n4878), .A(n4426), 
        .ZN(n5357) );
  XNOR2_X1 U1833 ( .A(n2545), .B(n4648), .ZN(J1epw6) );
  AOI221_X1 U1834 ( .B1(n4424), .B2(n5294), .C1(n2730), .C2(n4649), .A(n4426), 
        .ZN(n4648) );
  NAND4_X1 U1835 ( .A1(n5203), .A2(n5204), .A3(n5205), .A4(n5206), .ZN(n3059)
         );
  AOI22_X1 U1836 ( .A1(n5219), .A2(n5220), .B1(n417), .B2(n5221), .ZN(n5204)
         );
  NOR2_X1 U1837 ( .A1(n5207), .A2(n5208), .ZN(n5206) );
  AOI22_X1 U1838 ( .A1(n5222), .A2(n272), .B1(n1504), .B2(n4581), .ZN(n5203)
         );
  OAI222_X1 U1839 ( .A1(n4858), .A2(n3583), .B1(n4859), .B2(n5941), .C1(n623), 
        .C2(n2490), .ZN(n4901) );
  OAI222_X1 U1840 ( .A1(n4858), .A2(n3598), .B1(n4859), .B2(n5914), .C1(n4860), 
        .C2(n6241), .ZN(n4931) );
  OAI222_X1 U1841 ( .A1(n4858), .A2(n4278), .B1(n4859), .B2(n5960), .C1(n4860), 
        .C2(n6188), .ZN(n4945) );
  OAI222_X1 U1842 ( .A1(n627), .A2(n4181), .B1(n625), .B2(n5935), .C1(n4860), 
        .C2(n6264), .ZN(n5191) );
  OAI222_X1 U1843 ( .A1(n4858), .A2(n4178), .B1(n4859), .B2(n5915), .C1(n4860), 
        .C2(n6242), .ZN(n4857) );
  OAI222_X1 U1844 ( .A1(n627), .A2(n3591), .B1(n625), .B2(n5964), .C1(n4860), 
        .C2(n6212), .ZN(n5593) );
  OAI222_X1 U1845 ( .A1(n627), .A2(n4167), .B1(n625), .B2(n8251), .C1(n4860), 
        .C2(n6225), .ZN(n5143) );
  OAI222_X1 U1846 ( .A1(n627), .A2(n4007), .B1(n625), .B2(n5963), .C1(n4860), 
        .C2(n6210), .ZN(n5057) );
  OAI222_X1 U1847 ( .A1(n627), .A2(n3588), .B1(n625), .B2(n5956), .C1(n4860), 
        .C2(n6183), .ZN(n5361) );
  OAI222_X1 U1848 ( .A1(n627), .A2(n4086), .B1(n625), .B2(n5899), .C1(n4860), 
        .C2(n6229), .ZN(n5549) );
  OAI222_X1 U1849 ( .A1(n4858), .A2(n3611), .B1(n4859), .B2(n5938), .C1(n4860), 
        .C2(n6267), .ZN(n4969) );
  OAI222_X1 U1850 ( .A1(n3592), .A2(n627), .B1(n5990), .B2(n625), .C1(n2777), 
        .C2(n623), .ZN(n5768) );
  NOR2_X1 U1851 ( .A1(n678), .A2(n2633), .ZN(Tgfpw6[19]) );
  NOR2_X1 U1852 ( .A1(n4187), .A2(n3549), .ZN(n2376) );
  AOI21_X1 U1853 ( .B1(n4987), .B2(n4978), .A(n4669), .ZN(n4243) );
  NOR2_X1 U1854 ( .A1(n4187), .A2(n476), .ZN(n3527) );
  NOR2_X1 U1855 ( .A1(n679), .A2(n2631), .ZN(Tgfpw6[20]) );
  BUF_X1 U1856 ( .A(n4572), .Z(n464) );
  NAND2_X1 U1857 ( .A1(n435), .A2(n493), .ZN(n5214) );
  NOR2_X1 U1858 ( .A1(n678), .A2(n2630), .ZN(Tgfpw6[21]) );
  NOR3_X1 U1859 ( .A1(n3408), .A2(n3409), .A3(n3410), .ZN(n3407) );
  OR3_X1 U1860 ( .A1(n3411), .A2(n3412), .A3(n3413), .ZN(n3408) );
  NOR3_X1 U1861 ( .A1(n3392), .A2(n3393), .A3(n3394), .ZN(n3391) );
  NAND3_X1 U1862 ( .A1(n3395), .A2(n3396), .A3(n1552), .ZN(n3392) );
  INV_X1 U1863 ( .A(n3398), .ZN(n1552) );
  BUF_X1 U1864 ( .A(n5998), .Z(n567) );
  OAI22_X1 U1865 ( .A1(n4870), .A2(n6886), .B1(n4871), .B2(n6386), .ZN(n4935)
         );
  OAI22_X1 U1866 ( .A1(n4875), .A2(n7772), .B1(n4876), .B2(n5521), .ZN(n4953)
         );
  OAI22_X1 U1867 ( .A1(n4870), .A2(n3607), .B1(n577), .B2(n6355), .ZN(n5707)
         );
  OAI22_X1 U1868 ( .A1(n4870), .A2(n7603), .B1(n577), .B2(n6341), .ZN(n5379)
         );
  OAI22_X1 U1869 ( .A1(n4870), .A2(n6899), .B1(n4871), .B2(n6387), .ZN(n4869)
         );
  OAI22_X1 U1870 ( .A1(n4875), .A2(n7769), .B1(n4876), .B2(n5579), .ZN(n4927)
         );
  OAI22_X1 U1871 ( .A1(n4870), .A2(n7579), .B1(n577), .B2(n6328), .ZN(n5596)
         );
  OAI22_X1 U1872 ( .A1(n4870), .A2(n7342), .B1(n577), .B2(n6290), .ZN(n5170)
         );
  OAI22_X1 U1873 ( .A1(n4870), .A2(n7377), .B1(n4871), .B2(n6306), .ZN(n4964)
         );
  OAI22_X1 U1874 ( .A1(n4870), .A2(n4170), .B1(n577), .B2(n6372), .ZN(n5146)
         );
  OAI22_X1 U1875 ( .A1(n578), .A2(n7577), .B1(n577), .B2(n6329), .ZN(n5060) );
  OAI22_X1 U1876 ( .A1(n4870), .A2(n7573), .B1(n577), .B2(n6317), .ZN(n5364)
         );
  OAI22_X1 U1877 ( .A1(n4870), .A2(n7372), .B1(n4871), .B2(n6292), .ZN(n4904)
         );
  OAI22_X1 U1878 ( .A1(n4870), .A2(n7307), .B1(n4871), .B2(n6281), .ZN(n4972)
         );
  OAI22_X1 U1879 ( .A1(n4875), .A2(n7775), .B1(n4876), .B2(n5540), .ZN(n4886)
         );
  OAI22_X1 U1880 ( .A1(n4875), .A2(n7811), .B1(n4876), .B2(n5580), .ZN(n4897)
         );
  OAI22_X1 U1881 ( .A1(n4870), .A2(n8270), .B1(n577), .B2(n8267), .ZN(n5123)
         );
  OAI22_X1 U1882 ( .A1(n4870), .A2(n6918), .B1(n577), .B2(n6324), .ZN(n5440)
         );
  OAI22_X1 U1883 ( .A1(n572), .A2(n7815), .B1(n569), .B2(n5467), .ZN(n6440) );
  OAI22_X1 U1884 ( .A1(n572), .A2(n7754), .B1(n569), .B2(n5624), .ZN(n6429) );
  OAI22_X1 U1885 ( .A1(n572), .A2(n7781), .B1(n569), .B2(n5555), .ZN(n6436) );
  OAI22_X1 U1886 ( .A1(n572), .A2(n7751), .B1(n569), .B2(n5520), .ZN(n6444) );
  XNOR2_X1 U1887 ( .A(n4795), .B(n1977), .ZN(n1981) );
  NOR2_X1 U1888 ( .A1(n680), .A2(n2628), .ZN(Tgfpw6[23]) );
  INV_X1 U1889 ( .A(n5101), .ZN(n4078) );
  OAI22_X1 U1890 ( .A1(n564), .A2(n5718), .B1(n563), .B2(n6810), .ZN(n6463) );
  OAI22_X1 U1891 ( .A1(n6001), .A2(n5662), .B1(n6002), .B2(n6663), .ZN(n6099)
         );
  OAI22_X1 U1892 ( .A1(n6001), .A2(n5752), .B1(n6002), .B2(n6603), .ZN(n6095)
         );
  OAI22_X1 U1893 ( .A1(n564), .A2(n5799), .B1(n563), .B2(n6626), .ZN(n6471) );
  OAI22_X1 U1894 ( .A1(n564), .A2(n5682), .B1(n563), .B2(n6674), .ZN(n6467) );
  OAI22_X1 U1895 ( .A1(n6001), .A2(n5729), .B1(n6002), .B2(n6835), .ZN(n6087)
         );
  OAI22_X1 U1896 ( .A1(n6001), .A2(n5802), .B1(n6002), .B2(n6607), .ZN(n6459)
         );
  OAI22_X1 U1897 ( .A1(n6001), .A2(n5683), .B1(n6002), .B2(n6678), .ZN(n6091)
         );
  OAI22_X1 U1898 ( .A1(n5793), .A2(n564), .B1(n6863), .B2(n563), .ZN(n6501) );
  OAI22_X1 U1899 ( .A1(n5711), .A2(n564), .B1(n6668), .B2(n563), .ZN(n6496) );
  OAI22_X1 U1900 ( .A1(n5710), .A2(n564), .B1(n6657), .B2(n563), .ZN(n6010) );
  OAI22_X1 U1901 ( .A1(n5726), .A2(n564), .B1(n6600), .B2(n563), .ZN(n6507) );
  OAI22_X1 U1902 ( .A1(n5663), .A2(n564), .B1(n6638), .B2(n563), .ZN(n6522) );
  INV_X1 U1903 ( .A(n5984), .ZN(n2413) );
  INV_X1 U1904 ( .A(n2585), .ZN(n4669) );
  INV_X1 U1905 ( .A(n5323), .ZN(n2406) );
  NOR2_X1 U1906 ( .A1(n1907), .A2(n3527), .ZN(n1464) );
  NAND4_X1 U1907 ( .A1(n1799), .A2(n3420), .A3(n3421), .A4(n3422), .ZN(n3385)
         );
  INV_X1 U1908 ( .A(n3432), .ZN(n1799) );
  NOR3_X1 U1909 ( .A1(n3423), .A2(n3424), .A3(n3425), .ZN(n3422) );
  NOR3_X1 U1910 ( .A1(n3429), .A2(n3430), .A3(n3431), .ZN(n3421) );
  INV_X1 U1911 ( .A(n5943), .ZN(n2384) );
  INV_X1 U1912 ( .A(n5945), .ZN(n2403) );
  AOI22_X1 U1913 ( .A1(n878), .A2(n5212), .B1(n5213), .B2(n5225), .ZN(n5205)
         );
  OAI221_X1 U1914 ( .B1(n3800), .B2(n5214), .C1(n5215), .C2(n1528), .A(n4271), 
        .ZN(n5213) );
  AOI211_X1 U1915 ( .C1(n3077), .C2(n1538), .A(n5217), .B(n5218), .ZN(n5215)
         );
  NAND4_X1 U1916 ( .A1(n2873), .A2(n4194), .A3(n5223), .A4(n5224), .ZN(n5222)
         );
  AOI222_X1 U1917 ( .A1(n80), .A2(n266), .B1(n1478), .B2(n433), .C1(n474), 
        .C2(n4512), .ZN(n5224) );
  AOI22_X1 U1918 ( .A1(n3631), .A2(n5225), .B1(n429), .B2(n1663), .ZN(n5223)
         );
  INV_X1 U1919 ( .A(n3722), .ZN(n3631) );
  NAND2_X1 U1920 ( .A1(n1566), .A2(n435), .ZN(n3515) );
  INV_X1 U1921 ( .A(n4447), .ZN(n2326) );
  INV_X1 U1922 ( .A(n5536), .ZN(n2367) );
  INV_X1 U1923 ( .A(n5343), .ZN(n2347) );
  NOR2_X1 U1924 ( .A1(n680), .A2(n2626), .ZN(Tgfpw6[25]) );
  OAI22_X1 U1925 ( .A1(n3294), .A2(n2778), .B1(n3295), .B2(n2609), .ZN(Ksrhu6)
         );
  AOI222_X1 U1926 ( .A1(n101), .A2(n3297), .B1(n97), .B2(n1543), .C1(n99), 
        .C2(n224), .ZN(n3295) );
  INV_X1 U1927 ( .A(n4390), .ZN(n2459) );
  INV_X1 U1928 ( .A(n5538), .ZN(n2360) );
  INV_X1 U1929 ( .A(n5537), .ZN(n2370) );
  INV_X1 U1930 ( .A(n5342), .ZN(n2365) );
  INV_X1 U1931 ( .A(n5491), .ZN(n2460) );
  INV_X1 U1932 ( .A(n5283), .ZN(n2355) );
  INV_X1 U1933 ( .A(n4504), .ZN(n2474) );
  NOR2_X1 U1934 ( .A1(n679), .A2(n2625), .ZN(Tgfpw6[26]) );
  INV_X1 U1935 ( .A(n4747), .ZN(n3608) );
  BUF_X1 U1936 ( .A(n486), .Z(n485) );
  INV_X1 U1937 ( .A(n1977), .ZN(n2510) );
  INV_X1 U1938 ( .A(n5340), .ZN(n2387) );
  NOR2_X1 U1939 ( .A1(n679), .A2(n2624), .ZN(Tgfpw6[27]) );
  NOR2_X1 U1940 ( .A1(n679), .A2(n2636), .ZN(Tgfpw6[16]) );
  NOR2_X1 U1941 ( .A1(n2611), .A2(n2642), .ZN(Tgfpw6[10]) );
  NOR2_X1 U1942 ( .A1(n680), .A2(n2627), .ZN(Tgfpw6[24]) );
  NOR2_X1 U1943 ( .A1(n679), .A2(n2629), .ZN(Tgfpw6[22]) );
  AOI211_X1 U1944 ( .C1(n270), .C2(n5063), .A(n2932), .B(n2933), .ZN(n2931) );
  NAND3_X1 U1945 ( .A1(n5002), .A2(n4725), .A3(n2939), .ZN(n2930) );
  AOI22_X1 U1946 ( .A1(n2934), .A2(n2508), .B1(n98), .B2(n8260), .ZN(n2932) );
  NAND2_X1 U1947 ( .A1(n3515), .A2(n5265), .ZN(n5251) );
  NAND3_X1 U1948 ( .A1(n266), .A2(n516), .A3(n1566), .ZN(n5265) );
  INV_X1 U1949 ( .A(n4646), .ZN(n2411) );
  OAI21_X1 U1950 ( .B1(n25), .B2(n961), .A(n27), .ZN(n7726) );
  OAI21_X1 U1951 ( .B1(n28), .B2(n961), .A(n529), .ZN(n27) );
  NOR2_X1 U1952 ( .A1(n30), .A2(n31), .ZN(n25) );
  NAND4_X1 U1953 ( .A1(n66), .A2(n67), .A3(n68), .A4(n69), .ZN(n30) );
  INV_X1 U1954 ( .A(n3298), .ZN(n1543) );
  OAI21_X1 U1955 ( .B1(n3299), .B2(n5257), .A(n3301), .ZN(n3298) );
  OAI21_X1 U1956 ( .B1(n3302), .B2(n3303), .A(n5257), .ZN(n3301) );
  NOR4_X1 U1957 ( .A1(n3384), .A2(n3385), .A3(n3386), .A4(n3387), .ZN(n3299)
         );
  NOR2_X1 U1958 ( .A1(n679), .A2(n2623), .ZN(Tgfpw6[28]) );
  OAI221_X1 U1959 ( .B1(n1517), .B2(n33), .C1(n3766), .C2(n4738), .A(n36), 
        .ZN(n31) );
  AOI222_X1 U1960 ( .A1(n37), .A2(n38), .B1(n3550), .B2(n40), .C1(n41), .C2(
        n42), .ZN(n36) );
  INV_X1 U1961 ( .A(n65), .ZN(n1517) );
  OAI22_X1 U1962 ( .A1(n2528), .A2(n3749), .B1(n266), .B2(n2516), .ZN(n40) );
  INV_X1 U1963 ( .A(n4563), .ZN(n5273) );
  INV_X1 U1964 ( .A(n4562), .ZN(n5278) );
  INV_X1 U1965 ( .A(n5771), .ZN(n5282) );
  INV_X1 U1966 ( .A(n5550), .ZN(n5277) );
  NOR2_X1 U1967 ( .A1(n679), .A2(n2622), .ZN(Tgfpw6[29]) );
  NOR2_X1 U1968 ( .A1(n679), .A2(n2618), .ZN(Tgfpw6[3]) );
  NOR2_X1 U1969 ( .A1(n678), .A2(n2621), .ZN(Tgfpw6[2]) );
  NOR2_X1 U1970 ( .A1(n2611), .A2(n2613), .ZN(Tgfpw6[8]) );
  NOR2_X1 U1971 ( .A1(n679), .A2(n2620), .ZN(Tgfpw6[30]) );
  OAI221_X1 U1972 ( .B1(n3812), .B2(n3900), .C1(n1650), .C2(n3901), .A(n4279), 
        .ZN(\eq_3147/A[17] ) );
  NAND2_X1 U1973 ( .A1(N5fpw6[18]), .A2(n667), .ZN(n4279) );
  INV_X1 U1974 ( .A(Nxkbx6[20]), .ZN(n1650) );
  OAI221_X1 U1975 ( .B1(n3813), .B2(n3900), .C1(n1655), .C2(n3901), .A(n3916), 
        .ZN(\eq_3147/A[16] ) );
  NAND2_X1 U1976 ( .A1(N5fpw6[17]), .A2(n667), .ZN(n3916) );
  INV_X1 U1977 ( .A(Nxkbx6[19]), .ZN(n1655) );
  OAI221_X1 U1978 ( .B1(n3815), .B2(n664), .C1(n1677), .C2(n661), .A(n4045), 
        .ZN(\eq_3147/A[14] ) );
  NAND2_X1 U1979 ( .A1(N5fpw6[15]), .A2(n667), .ZN(n4045) );
  INV_X1 U1980 ( .A(Nxkbx6[17]), .ZN(n1677) );
  NOR2_X1 U1981 ( .A1(n679), .A2(n2619), .ZN(Tgfpw6[31]) );
  NAND4_X1 U1982 ( .A1(\add_3107/B[1] ), .A2(n952), .A3(n3895), .A4(Tnhpw6[0]), 
        .ZN(n3921) );
  OR3_X1 U1983 ( .A1(n3424), .A2(Affpw6[2]), .A3(n3442), .ZN(n4613) );
  NOR3_X1 U1984 ( .A1(n5065), .A2(n3576), .A3(n3571), .ZN(n2806) );
  OAI221_X1 U1985 ( .B1(n3817), .B2(n3900), .C1(n1696), .C2(n661), .A(n4201), 
        .ZN(\eq_3147/A[12] ) );
  NAND2_X1 U1986 ( .A1(N5fpw6[13]), .A2(n667), .ZN(n4201) );
  OAI221_X1 U1987 ( .B1(n3818), .B2(n664), .C1(n1717), .C2(n3901), .A(n3970), 
        .ZN(\eq_3147/A[11] ) );
  NAND2_X1 U1988 ( .A1(N5fpw6[12]), .A2(n667), .ZN(n3970) );
  NOR2_X2 U1989 ( .A1(n211), .A2(n3409), .ZN(n2217) );
  NOR2_X2 U1990 ( .A1(n224), .A2(n3398), .ZN(n2404) );
  AND2_X1 U1991 ( .A1(n3892), .A2(n3893), .ZN(HSIZE[1]) );
  OAI211_X1 U1992 ( .C1(n2693), .C2(n669), .A(n946), .B(n2154), .ZN(n3893) );
  OAI221_X1 U1993 ( .B1(n3819), .B2(n664), .C1(n1719), .C2(n3901), .A(n3918), 
        .ZN(\eq_3147/A[10] ) );
  NAND2_X1 U1994 ( .A1(N5fpw6[11]), .A2(n667), .ZN(n3918) );
  OAI221_X1 U1995 ( .B1(n3820), .B2(n664), .C1(n1764), .C2(n3901), .A(n4031), 
        .ZN(\eq_3147/A[9] ) );
  NAND2_X1 U1996 ( .A1(N5fpw6[10]), .A2(n667), .ZN(n4031) );
  OAI221_X1 U1997 ( .B1(n3821), .B2(n664), .C1(n1767), .C2(n661), .A(n3919), 
        .ZN(\eq_3147/A[8] ) );
  NAND2_X1 U1998 ( .A1(N5fpw6[9]), .A2(n667), .ZN(n3919) );
  OAI221_X1 U1999 ( .B1(n3791), .B2(n664), .C1(n1775), .C2(n661), .A(n3950), 
        .ZN(\eq_3147/A[6] ) );
  NAND2_X1 U2000 ( .A1(N5fpw6[7]), .A2(n667), .ZN(n3950) );
  OAI221_X1 U2001 ( .B1(n3792), .B2(n664), .C1(n1783), .C2(n3901), .A(n3902), 
        .ZN(\eq_3147/A[5] ) );
  NAND2_X1 U2002 ( .A1(N5fpw6[6]), .A2(n669), .ZN(n3902) );
  OAI221_X1 U2003 ( .B1(n3793), .B2(n664), .C1(n1786), .C2(n3901), .A(n4404), 
        .ZN(\eq_3147/A[4] ) );
  NAND2_X1 U2004 ( .A1(N5fpw6[5]), .A2(n667), .ZN(n4404) );
  OAI222_X1 U2005 ( .A1(n3315), .A2(n5387), .B1(n2713), .B2(n8307), .C1(n742), 
        .C2(n2712), .ZN(n4350) );
  OAI221_X1 U2006 ( .B1(n4332), .B2(n3458), .C1(n2813), .C2(n4334), .A(n2544), 
        .ZN(D5epw6) );
  INV_X1 U2007 ( .A(n3458), .ZN(n2813) );
  AOI221_X1 U2008 ( .B1(n4424), .B2(n3571), .C1(n2730), .C2(n4988), .A(n4426), 
        .ZN(n5609) );
  AOI221_X1 U2009 ( .B1(n4424), .B2(n3576), .C1(n2730), .C2(n4603), .A(n4426), 
        .ZN(n4601) );
  AOI221_X1 U2010 ( .B1(n4424), .B2(n5065), .C1(n2730), .C2(n4666), .A(n4426), 
        .ZN(n4686) );
  OAI21_X1 U2011 ( .B1(n6318), .B2(n6319), .A(n6320), .ZN(n6118) );
  NAND3_X1 U2012 ( .A1(n6321), .A2(n6322), .A3(n3925), .ZN(n6320) );
  AOI22_X1 U2013 ( .A1(n6323), .A2(n3061), .B1(n6305), .B2(n6307), .ZN(n6319)
         );
  AOI21_X1 U2014 ( .B1(n3925), .B2(n4420), .A(n6314), .ZN(n6323) );
  OAI221_X1 U2015 ( .B1(n2326), .B2(n3900), .C1(n1770), .C2(n3901), .A(n5413), 
        .ZN(\eq_3147/A[7] ) );
  NAND2_X1 U2016 ( .A1(N5fpw6[8]), .A2(n667), .ZN(n5413) );
  OAI221_X1 U2017 ( .B1(n3794), .B2(n3900), .C1(n1790), .C2(n661), .A(n3903), 
        .ZN(\eq_3147/A[3] ) );
  NAND2_X1 U2018 ( .A1(N5fpw6[4]), .A2(n669), .ZN(n3903) );
  OAI221_X1 U2019 ( .B1(n1795), .B2(n661), .C1(n3795), .C2(n3900), .A(n5104), 
        .ZN(\eq_3147/A[2] ) );
  NAND2_X1 U2020 ( .A1(N5fpw6[3]), .A2(n667), .ZN(n5104) );
  OAI221_X1 U2021 ( .B1(n2138), .B2(n4343), .C1(n4344), .C2(n2724), .A(n4345), 
        .ZN(n211) );
  AOI221_X1 U2022 ( .B1(n2339), .B2(n4346), .C1(n4347), .C2(n2363), .A(n4349), 
        .ZN(n4345) );
  OAI221_X1 U2023 ( .B1(n4522), .B2(n2716), .C1(n4343), .C2(n4523), .A(n5442), 
        .ZN(n224) );
  AOI221_X1 U2024 ( .B1(n4346), .B2(n4525), .C1(n4653), .C2(n4527), .A(n4349), 
        .ZN(n5442) );
  OAI221_X1 U2025 ( .B1(n2716), .B2(n4593), .C1(n4343), .C2(n4594), .A(n4817), 
        .ZN(n232) );
  AOI221_X1 U2026 ( .B1(n4653), .B2(n2207), .C1(n4590), .C2(n4346), .A(n4349), 
        .ZN(n4817) );
  OAI221_X1 U2027 ( .B1(n2415), .B2(n4343), .C1(n4638), .C2(n2724), .A(n5125), 
        .ZN(n100) );
  AOI221_X1 U2028 ( .B1(n4346), .B2(n2443), .C1(n4347), .C2(n2345), .A(n4349), 
        .ZN(n5125) );
  OAI221_X1 U2029 ( .B1(n4332), .B2(n3297), .C1(n2759), .C2(n4334), .A(n2544), 
        .ZN(Qbfpw6[30]) );
  INV_X1 U2030 ( .A(n3297), .ZN(n2759) );
  NOR2_X1 U2031 ( .A1(n3968), .A2(n5112), .ZN(n5255) );
  OAI222_X1 U2032 ( .A1(n2702), .A2(n8260), .B1(n4376), .B2(n442), .C1(n439), 
        .C2(n1581), .ZN(n3416) );
  OAI221_X1 U2033 ( .B1(n4332), .B2(n4939), .C1(n3602), .C2(n4334), .A(n2544), 
        .ZN(Qbfpw6[27]) );
  OAI221_X1 U2034 ( .B1(n4332), .B2(n4496), .C1(n3329), .C2(n4334), .A(n2544), 
        .ZN(Qbfpw6[25]) );
  OAI221_X1 U2035 ( .B1(n4332), .B2(n4678), .C1(n4063), .C2(n4334), .A(n2544), 
        .ZN(Qbfpw6[26]) );
  NOR2_X1 U2036 ( .A1(n6287), .A2(n6288), .ZN(n5303) );
  AOI21_X1 U2037 ( .B1(n3669), .B2(n8148), .A(n3668), .ZN(n6288) );
  AOI211_X1 U2038 ( .C1(n3666), .C2(n6262), .A(n3661), .B(n6261), .ZN(n6287)
         );
  INV_X1 U2039 ( .A(n6293), .ZN(n3661) );
  OAI221_X1 U2040 ( .B1(n4332), .B2(n102), .C1(n4376), .C2(n4334), .A(n2544), 
        .ZN(Qbfpw6[28]) );
  NOR2_X1 U2041 ( .A1(n5074), .A2(n3566), .ZN(n2807) );
  OAI221_X1 U2042 ( .B1(n4332), .B2(n4956), .C1(n3483), .C2(n4334), .A(n2544), 
        .ZN(Qbfpw6[24]) );
  OAI21_X1 U2043 ( .B1(n6213), .B2(n6214), .A(n6215), .ZN(n6143) );
  AND2_X1 U2044 ( .A1(n6141), .A2(n6211), .ZN(n6213) );
  OR3_X1 U2045 ( .A1(n6216), .A2(n6217), .A3(n3117), .ZN(n6215) );
  AOI22_X1 U2046 ( .A1(n2793), .A2(n6200), .B1(n6206), .B2(n2794), .ZN(n6214)
         );
  NAND2_X1 U2047 ( .A1(n474), .A2(n56), .ZN(n1572) );
  OAI22_X1 U2048 ( .A1(n6262), .A2(n5303), .B1(n6263), .B2(n3659), .ZN(n6209)
         );
  AND4_X1 U2049 ( .A1(n2851), .A2(n1972), .A3(n2850), .A4(n4060), .ZN(n4056)
         );
  NOR4_X1 U2050 ( .A1(n1527), .A2(n1526), .A3(n717), .A4(n1834), .ZN(n4060) );
  INV_X1 U2051 ( .A(n1961), .ZN(n1834) );
  OAI22_X1 U2052 ( .A1(n1814), .A2(n661), .B1(n3822), .B2(n3900), .ZN(n466) );
  OAI22_X1 U2053 ( .A1(n3120), .A2(n8246), .B1(n8233), .B2(n6233), .ZN(n6226)
         );
  INV_X1 U2054 ( .A(LOCKUP), .ZN(n2548) );
  NAND4_X1 U2055 ( .A1(n5780), .A2(n2444), .A3(n5781), .A4(n5782), .ZN(n5560)
         );
  NAND4_X1 U2056 ( .A1(n2185), .A2(n522), .A3(n4263), .A4(n265), .ZN(n5780) );
  OR3_X1 U2057 ( .A1(n503), .A2(n5787), .A3(n3730), .ZN(n5781) );
  AOI221_X1 U2058 ( .B1(n5783), .B2(n2363), .C1(n5220), .C2(n5784), .A(n5785), 
        .ZN(n5782) );
  AOI22_X1 U2059 ( .A1(n6132), .A2(n4282), .B1(n3640), .B2(n3638), .ZN(n6316)
         );
  AOI22_X1 U2060 ( .A1(n5321), .A2(n6327), .B1(n3063), .B2(n3062), .ZN(n6305)
         );
  OAI221_X1 U2061 ( .B1(n4332), .B2(n4531), .C1(n3032), .C2(n4334), .A(n2544), 
        .ZN(Qbfpw6[29]) );
  OAI22_X1 U2062 ( .A1(n2274), .A2(n2231), .B1(n755), .B2(n6387), .ZN(C4qhu6)
         );
  OAI22_X1 U2063 ( .A1(n2327), .A2(n2231), .B1(n755), .B2(n6377), .ZN(Gbshu6)
         );
  OAI22_X1 U2064 ( .A1(n2323), .A2(n2231), .B1(n755), .B2(n6372), .ZN(Gdqhu6)
         );
  OAI22_X1 U2065 ( .A1(n2284), .A2(n2231), .B1(n755), .B2(n6355), .ZN(Gxrhu6)
         );
  OAI22_X1 U2066 ( .A1(n2311), .A2(n2231), .B1(n755), .B2(n6329), .ZN(Nlphu6)
         );
  OAI22_X1 U2067 ( .A1(n2340), .A2(n2231), .B1(n755), .B2(n6328), .ZN(Nzphu6)
         );
  OAI22_X1 U2068 ( .A1(n2331), .A2(n2231), .B1(n755), .B2(n6317), .ZN(R8qhu6)
         );
  OAI22_X1 U2069 ( .A1(n2278), .A2(n2231), .B1(n755), .B2(n6306), .ZN(V1shu6)
         );
  OAI22_X1 U2070 ( .A1(n2205), .A2(n2231), .B1(n755), .B2(n6281), .ZN(Yuphu6)
         );
  OAI221_X1 U2071 ( .B1(n4632), .B2(n2715), .C1(n2415), .C2(n2718), .A(n4634), 
        .ZN(n337) );
  AOI221_X1 U2072 ( .B1(n4440), .B2(n2345), .C1(n4636), .C2(n2175), .A(n2158), 
        .ZN(n4634) );
  INV_X1 U2073 ( .A(n4638), .ZN(n2175) );
  OAI221_X1 U2074 ( .B1(n2429), .B2(n2715), .C1(n2718), .C2(n2389), .A(n4689), 
        .ZN(n347) );
  AOI221_X1 U2075 ( .B1(n4440), .B2(n2350), .C1(n4636), .C2(n2383), .A(n2158), 
        .ZN(n4689) );
  OAI221_X1 U2076 ( .B1(n4593), .B2(n2720), .C1(n2718), .C2(n4594), .A(n5267), 
        .ZN(n331) );
  AOI221_X1 U2077 ( .B1(n4636), .B2(n2207), .C1(n4439), .C2(n4590), .A(n2158), 
        .ZN(n5267) );
  OAI221_X1 U2078 ( .B1(n3780), .B2(n442), .C1(n439), .C2(n1614), .A(n4155), 
        .ZN(n3440) );
  AOI221_X1 U2079 ( .B1(n4156), .B2(n2745), .C1(n2279), .C2(n4159), .A(
        Affpw6[23]), .ZN(n4155) );
  OAI22_X1 U2080 ( .A1(n2549), .A2(Qbfpw6[23]), .B1(n2550), .B2(n4162), .ZN(
        n4159) );
  OAI21_X1 U2081 ( .B1(n2279), .B2(n4162), .A(n243), .ZN(n4156) );
  OAI221_X1 U2082 ( .B1(n4412), .B2(n2703), .C1(n4411), .C2(n2719), .A(n4630), 
        .ZN(n402) );
  AOI221_X1 U2083 ( .B1(n4267), .B2(n4416), .C1(n4269), .C2(n4414), .A(n2148), 
        .ZN(n4630) );
  OAI221_X1 U2084 ( .B1(n4344), .B2(n2719), .C1(n4143), .C2(n2703), .A(n5176), 
        .ZN(n368) );
  AOI221_X1 U2085 ( .B1(n4269), .B2(n2339), .C1(n4267), .C2(n4350), .A(n2148), 
        .ZN(n5176) );
  OAI221_X1 U2086 ( .B1(n4522), .B2(n2720), .C1(n2718), .C2(n4523), .A(n5130), 
        .ZN(n325) );
  AOI221_X1 U2087 ( .B1(n4439), .B2(n4525), .C1(n4636), .C2(n4527), .A(n2158), 
        .ZN(n5130) );
  OAI221_X1 U2088 ( .B1(n5553), .B2(n4343), .C1(n4837), .C2(n2724), .A(n5655), 
        .ZN(n246) );
  AOI221_X1 U2089 ( .B1(n4346), .B2(n4840), .C1(n4347), .C2(n2341), .A(n4349), 
        .ZN(n5655) );
  OAI221_X1 U2090 ( .B1(n2435), .B2(n2715), .C1(n5553), .C2(n2718), .A(n5554), 
        .ZN(n341) );
  AOI221_X1 U2091 ( .B1(n4440), .B2(n2341), .C1(n4636), .C2(n2385), .A(n2158), 
        .ZN(n5554) );
  OAI221_X1 U2092 ( .B1(n2718), .B2(n2204), .C1(n4264), .C2(n2708), .A(n4438), 
        .ZN(n358) );
  AOI221_X1 U2093 ( .B1(n4439), .B2(n4270), .C1(n4440), .C2(n2351), .A(n2158), 
        .ZN(n4438) );
  OAI221_X1 U2094 ( .B1(n4343), .B2(n2204), .C1(n4264), .C2(n2724), .A(n4492), 
        .ZN(n263) );
  AOI221_X1 U2095 ( .B1(n4270), .B2(n4346), .C1(n2351), .C2(n4347), .A(n4349), 
        .ZN(n4492) );
  OAI221_X1 U2096 ( .B1(n5127), .B2(n2703), .C1(n4638), .C2(n2719), .A(n5777), 
        .ZN(n386) );
  AOI221_X1 U2097 ( .B1(n4267), .B2(n4654), .C1(n4269), .C2(n2443), .A(n2148), 
        .ZN(n5777) );
  OAI221_X1 U2098 ( .B1(n4393), .B2(n2708), .C1(n2718), .C2(n2203), .A(n5043), 
        .ZN(n362) );
  AOI221_X1 U2099 ( .B1(n4440), .B2(n4398), .C1(n4439), .C2(n4399), .A(n2158), 
        .ZN(n5043) );
  AOI22_X1 U2100 ( .A1(n4435), .A2(n6145), .B1(n6226), .B2(n3117), .ZN(n6206)
         );
  NOR3_X1 U2101 ( .A1(n4205), .A2(n272), .A3(n4826), .ZN(n4235) );
  OAI221_X1 U2102 ( .B1(n6200), .B2(n6143), .C1(n6201), .C2(n2789), .A(n6203), 
        .ZN(n6190) );
  OR3_X1 U2103 ( .A1(n2792), .A2(n6204), .A3(n6141), .ZN(n6203) );
  INV_X1 U2104 ( .A(n5310), .ZN(n2789) );
  AOI221_X1 U2105 ( .B1(n7381), .B2(n4187), .C1(n476), .C2(n3549), .A(n4635), 
        .ZN(n5264) );
  NOR2_X1 U2106 ( .A1(n3797), .A2(n3789), .ZN(Idfpw6[31]) );
  NOR2_X1 U2107 ( .A1(n6333), .A2(n6334), .ZN(n6311) );
  AOI21_X1 U2108 ( .B1(n8153), .B2(n3930), .A(n3928), .ZN(n6333) );
  AOI221_X1 U2109 ( .B1(n6335), .B2(n3926), .C1(n6322), .C2(n6321), .A(n6336), 
        .ZN(n6334) );
  AOI22_X1 U2110 ( .A1(n4420), .A2(n6312), .B1(n6337), .B2(n4431), .ZN(n6336)
         );
  INV_X1 U2111 ( .A(n56), .ZN(n3550) );
  OAI222_X1 U2112 ( .A1(n4858), .A2(n3586), .B1(n4859), .B2(n5948), .C1(n623), 
        .C2(n6177), .ZN(n4923) );
  OAI222_X1 U2113 ( .A1(n4858), .A2(n8184), .B1(n4859), .B2(n8189), .C1(n623), 
        .C2(n8181), .ZN(n4914) );
  OAI222_X1 U2114 ( .A1(n4858), .A2(n3781), .B1(n4859), .B2(n5959), .C1(n4860), 
        .C2(n6207), .ZN(n4949) );
  OAI222_X1 U2115 ( .A1(n627), .A2(n3596), .B1(n625), .B2(n5901), .C1(n4860), 
        .C2(n6234), .ZN(n5376) );
  OAI222_X1 U2116 ( .A1(n627), .A2(n3581), .B1(n625), .B2(n5940), .C1(n4860), 
        .C2(n6271), .ZN(n5167) );
  OAI222_X1 U2117 ( .A1(n4858), .A2(n4066), .B1(n4859), .B2(n5961), .C1(n4860), 
        .C2(n6202), .ZN(n4961) );
  OAI222_X1 U2118 ( .A1(n627), .A2(n3864), .B1(n625), .B2(n5905), .C1(n4860), 
        .C2(n6239), .ZN(n5617) );
  OAI222_X1 U2119 ( .A1(n627), .A2(n3650), .B1(n625), .B2(n3653), .C1(n4860), 
        .C2(n6220), .ZN(n5006) );
  OAI222_X1 U2120 ( .A1(n627), .A2(n8211), .B1(n625), .B2(n8216), .C1(n4860), 
        .C2(n8208), .ZN(n4997) );
  OAI222_X1 U2121 ( .A1(n627), .A2(n3279), .B1(n625), .B2(n5924), .C1(n4860), 
        .C2(n6257), .ZN(n4982) );
  OAI222_X1 U2122 ( .A1(n627), .A2(n4003), .B1(n625), .B2(n5989), .C1(n4860), 
        .C2(n6218), .ZN(n5082) );
  OAI221_X1 U2123 ( .B1(n4063), .B2(n448), .C1(n439), .C2(n1597), .A(n4675), 
        .ZN(n3431) );
  AOI211_X1 U2124 ( .C1(n4676), .C2(Qbfpw6[26]), .A(Affpw6[26]), .B(n4677), 
        .ZN(n4675) );
  OAI22_X1 U2125 ( .A1(n2550), .A2(n2328), .B1(n4446), .B2(n4679), .ZN(n4676)
         );
  NOR3_X1 U2126 ( .A1(n2328), .A2(Qbfpw6[26]), .A3(n2549), .ZN(n4677) );
  NAND2_X1 U2127 ( .A1(n5867), .A2(n5868), .ZN(n2472) );
  NAND2_X1 U2128 ( .A1(n5863), .A2(n5243), .ZN(n3449) );
  NAND2_X1 U2129 ( .A1(n5867), .A2(n5861), .ZN(n3862) );
  NAND3_X1 U2130 ( .A1(n5255), .A2(n5111), .A3(n5862), .ZN(n1636) );
  OAI22_X1 U2131 ( .A1(n659), .A2(n3335), .B1(n650), .B2(n4498), .ZN(n4497) );
  NOR3_X1 U2132 ( .A1(n4499), .A2(n4500), .A3(n4501), .ZN(n4498) );
  OAI22_X1 U2133 ( .A1(n4288), .A2(n8097), .B1(n4291), .B2(n8066), .ZN(n4501)
         );
  OAI222_X1 U2134 ( .A1(n4502), .A2(n5834), .B1(n4503), .B2(n3324), .C1(n646), 
        .C2(n8119), .ZN(n4500) );
  NAND3_X1 U2135 ( .A1(n2307), .A2(n4069), .A3(N439), .ZN(n111) );
  OAI21_X1 U2136 ( .B1(n2616), .B2(n4064), .A(n4071), .ZN(n4069) );
  NAND4_X1 U2137 ( .A1(n736), .A2(n477), .A3(n4667), .A4(n5284), .ZN(n4071) );
  NAND3_X1 U2138 ( .A1(n2333), .A2(n4062), .A3(N438), .ZN(n124) );
  OAI21_X1 U2139 ( .B1(n2615), .B2(n4064), .A(n4065), .ZN(n4062) );
  NAND4_X1 U2140 ( .A1(n697), .A2(n477), .A3(n4667), .A4(n5284), .ZN(n4065) );
  OAI22_X1 U2141 ( .A1(n5900), .A2(n2219), .B1(n5457), .B2(n2220), .ZN(n5803)
         );
  INV_X1 U2142 ( .A(n5902), .ZN(n2220) );
  NAND2_X1 U2143 ( .A1(n5861), .A2(n5243), .ZN(n4843) );
  AOI22_X1 U2144 ( .A1(n4436), .A2(n6145), .B1(n3118), .B2(n3117), .ZN(n6200)
         );
  INV_X1 U2145 ( .A(n6222), .ZN(n4436) );
  NAND2_X1 U2146 ( .A1(n5864), .A2(n5243), .ZN(n3778) );
  AOI22_X1 U2147 ( .A1(n6141), .A2(n2799), .B1(n3033), .B2(n2797), .ZN(n6205)
         );
  NAND2_X1 U2148 ( .A1(n5867), .A2(n5878), .ZN(n3199) );
  NAND2_X1 U2149 ( .A1(n5867), .A2(n5869), .ZN(n3742) );
  AOI22_X1 U2150 ( .A1(n8244), .A2(n6125), .B1(n8230), .B2(n3064), .ZN(n6350)
         );
  NAND2_X1 U2151 ( .A1(n5863), .A2(n5867), .ZN(n3558) );
  NAND2_X1 U2152 ( .A1(n5889), .A2(n5867), .ZN(n4276) );
  NAND4_X1 U2153 ( .A1(n5824), .A2(n3936), .A3(n5826), .A4(n5827), .ZN(n5262)
         );
  AOI221_X1 U2154 ( .B1(n3934), .B2(n8199), .C1(n3987), .C2(n8256), .A(n5850), 
        .ZN(n5824) );
  NOR4_X1 U2155 ( .A1(n5841), .A2(n5842), .A3(n5843), .A4(n5844), .ZN(n5826)
         );
  INV_X1 U2156 ( .A(n5845), .ZN(n3936) );
  INV_X1 U2157 ( .A(n4426), .ZN(n2597) );
  NAND2_X1 U2158 ( .A1(n5889), .A2(n5243), .ZN(n3639) );
  NAND2_X1 U2159 ( .A1(n131), .A2(n132), .ZN(n128) );
  OAI211_X1 U2160 ( .C1(n133), .C2(n134), .A(n135), .B(HSIZE[1]), .ZN(n132) );
  NOR4_X1 U2161 ( .A1(n170), .A2(n1726), .A3(n1772), .A4(n328), .ZN(n133) );
  AOI21_X1 U2162 ( .B1(n154), .B2(n155), .A(HADDR[5]), .ZN(n134) );
  NAND2_X1 U2163 ( .A1(n5870), .A2(n5798), .ZN(n2526) );
  OAI22_X1 U2164 ( .A1(n761), .A2(n8119), .B1(n2252), .B2(n757), .ZN(Pkrhu6)
         );
  OAI22_X1 U2165 ( .A1(n761), .A2(n8101), .B1(n2228), .B2(n2229), .ZN(Zrphu6)
         );
  OAI22_X1 U2166 ( .A1(n683), .A2(n8097), .B1(n2252), .B2(n2362), .ZN(Fmrhu6)
         );
  OAI22_X1 U2167 ( .A1(n683), .A2(n8086), .B1(n2228), .B2(n2362), .ZN(Ptphu6)
         );
  OAI22_X1 U2168 ( .A1(n768), .A2(n8066), .B1(n2252), .B2(n764), .ZN(Ikrhu6)
         );
  OAI22_X1 U2169 ( .A1(n767), .A2(n8056), .B1(n2228), .B2(n2218), .ZN(Srphu6)
         );
  OAI22_X1 U2170 ( .A1(n714), .A2(n7769), .B1(n2252), .B2(n2285), .ZN(Rlrhu6)
         );
  OAI22_X1 U2171 ( .A1(n688), .A2(n7571), .B1(n2252), .B2(n2344), .ZN(Njrhu6)
         );
  OAI22_X1 U2172 ( .A1(n690), .A2(n6886), .B1(n2228), .B2(n2344), .ZN(Xqphu6)
         );
  OAI22_X1 U2173 ( .A1(n738), .A2(n6674), .B1(n2228), .B2(n2253), .ZN(Jqphu6)
         );
  OAI22_X1 U2174 ( .A1(n739), .A2(n6599), .B1(n2252), .B2(n737), .ZN(Zirhu6)
         );
  OAI22_X1 U2175 ( .A1(n780), .A2(n6588), .B1(n2252), .B2(n776), .ZN(Dlrhu6)
         );
  OAI22_X1 U2176 ( .A1(n779), .A2(n6524), .B1(n2228), .B2(n776), .ZN(Nsphu6)
         );
  OAI22_X1 U2177 ( .A1(n755), .A2(n6386), .B1(n2228), .B2(n2231), .ZN(Cqphu6)
         );
  OAI22_X1 U2178 ( .A1(n753), .A2(n6313), .B1(n2252), .B2(n751), .ZN(Sirhu6)
         );
  OAI22_X1 U2179 ( .A1(n706), .A2(n6241), .B1(n2228), .B2(n2289), .ZN(Itphu6)
         );
  OAI22_X1 U2180 ( .A1(n709), .A2(n6177), .B1(n2252), .B2(n2289), .ZN(Ylrhu6)
         );
  OAI22_X1 U2181 ( .A1(n685), .A2(n6142), .B1(n2228), .B2(n684), .ZN(Lrphu6)
         );
  OAI22_X1 U2182 ( .A1(n403), .A2(n5948), .B1(n2252), .B2(n729), .ZN(Mmrhu6)
         );
  OAI22_X1 U2183 ( .A1(n403), .A2(n5914), .B1(n2228), .B2(n722), .ZN(Wtphu6)
         );
  OAI22_X1 U2184 ( .A1(n775), .A2(n5891), .B1(n2228), .B2(n771), .ZN(Erphu6)
         );
  OAI22_X1 U2185 ( .A1(n775), .A2(n5834), .B1(n2252), .B2(n2214), .ZN(Ujrhu6)
         );
  OAI22_X1 U2186 ( .A1(n749), .A2(n5736), .B1(n2252), .B2(n2237), .ZN(Klrhu6)
         );
  OAI22_X1 U2187 ( .A1(n748), .A2(n5682), .B1(n2228), .B2(n2237), .ZN(Usphu6)
         );
  OAI22_X1 U2188 ( .A1(n695), .A2(n5579), .B1(n2252), .B2(n691), .ZN(Gjrhu6)
         );
  OAI22_X1 U2189 ( .A1(n695), .A2(n5523), .B1(n2228), .B2(n691), .ZN(Qqphu6)
         );
  OAI22_X1 U2190 ( .A1(n743), .A2(n5428), .B1(n2228), .B2(n2249), .ZN(Gsphu6)
         );
  OAI22_X1 U2191 ( .A1(n744), .A2(n5326), .B1(n2252), .B2(n2249), .ZN(Wkrhu6)
         );
  OAI22_X1 U2192 ( .A1(n787), .A2(n3598), .B1(n2228), .B2(n784), .ZN(Duphu6)
         );
  OAI22_X1 U2193 ( .A1(n399), .A2(n3586), .B1(n2252), .B2(n783), .ZN(Tmrhu6)
         );
  OAI22_X1 U2194 ( .A1(n714), .A2(n3341), .B1(n2228), .B2(n2285), .ZN(Btphu6)
         );
  OAI22_X1 U2195 ( .A1(n686), .A2(n3324), .B1(n2252), .B2(n684), .ZN(Bkrhu6)
         );
  NAND2_X1 U2196 ( .A1(n5864), .A2(n5255), .ZN(n4121) );
  OAI22_X1 U2197 ( .A1(n683), .A2(n8282), .B1(n2278), .B2(n2362), .ZN(B5shu6)
         );
  OAI22_X1 U2198 ( .A1(n403), .A2(n8251), .B1(n2323), .B2(n729), .ZN(Ahqhu6)
         );
  OAI22_X1 U2199 ( .A1(n761), .A2(n8132), .B1(n2323), .B2(n757), .ZN(Dfqhu6)
         );
  OAI22_X1 U2200 ( .A1(n760), .A2(n8126), .B1(n2340), .B2(n757), .ZN(K1qhu6)
         );
  OAI22_X1 U2201 ( .A1(n760), .A2(n8125), .B1(n2311), .B2(n757), .ZN(Knphu6)
         );
  OAI22_X1 U2202 ( .A1(n761), .A2(n8123), .B1(n2278), .B2(n757), .ZN(L3shu6)
         );
  OAI22_X1 U2203 ( .A1(n760), .A2(n8121), .B1(n2331), .B2(n757), .ZN(Oaqhu6)
         );
  OAI22_X1 U2204 ( .A1(n761), .A2(n8113), .B1(n2205), .B2(n2229), .ZN(Vwphu6)
         );
  OAI22_X1 U2205 ( .A1(n761), .A2(n8112), .B1(n2327), .B2(n2229), .ZN(Wcshu6)
         );
  OAI22_X1 U2206 ( .A1(n760), .A2(n8107), .B1(n2284), .B2(n2229), .ZN(Wyrhu6)
         );
  OAI22_X1 U2207 ( .A1(n761), .A2(n8102), .B1(n2274), .B2(n2229), .ZN(Z5qhu6)
         );
  OAI22_X1 U2208 ( .A1(n683), .A2(n8092), .B1(n2284), .B2(n2362), .ZN(M0shu6)
         );
  OAI22_X1 U2209 ( .A1(n768), .A2(n8071), .B1(n2278), .B2(n764), .ZN(E3shu6)
         );
  OAI22_X1 U2210 ( .A1(n768), .A2(n8058), .B1(n2284), .B2(n2218), .ZN(Pyrhu6)
         );
  OAI22_X1 U2211 ( .A1(n714), .A2(n7806), .B1(n2323), .B2(n2285), .ZN(Fgqhu6)
         );
  OAI22_X1 U2212 ( .A1(n713), .A2(n7790), .B1(n2340), .B2(n2285), .ZN(M2qhu6)
         );
  OAI22_X1 U2213 ( .A1(n713), .A2(n7787), .B1(n2311), .B2(n2285), .ZN(Mophu6)
         );
  OAI22_X1 U2214 ( .A1(n714), .A2(n7784), .B1(n2278), .B2(n2285), .ZN(N4shu6)
         );
  OAI22_X1 U2215 ( .A1(n713), .A2(n7778), .B1(n2331), .B2(n2285), .ZN(Qbqhu6)
         );
  OAI22_X1 U2216 ( .A1(n713), .A2(n7757), .B1(n2205), .B2(n2285), .ZN(Xxphu6)
         );
  OAI22_X1 U2217 ( .A1(n714), .A2(n7751), .B1(n2327), .B2(n2285), .ZN(Ydshu6)
         );
  OAI22_X1 U2218 ( .A1(n713), .A2(n7704), .B1(n2284), .B2(n2285), .ZN(Yzrhu6)
         );
  OAI22_X1 U2219 ( .A1(n688), .A2(n7695), .B1(n2327), .B2(n2344), .ZN(Bcshu6)
         );
  OAI22_X1 U2220 ( .A1(n688), .A2(n7579), .B1(n2340), .B2(n2344), .ZN(I0qhu6)
         );
  OAI22_X1 U2221 ( .A1(n690), .A2(n7577), .B1(n2311), .B2(n2344), .ZN(Imphu6)
         );
  OAI22_X1 U2222 ( .A1(n688), .A2(n7573), .B1(n2331), .B2(n2344), .ZN(M9qhu6)
         );
  OAI22_X1 U2223 ( .A1(n688), .A2(n7377), .B1(n2278), .B2(n2344), .ZN(Q2shu6)
         );
  OAI22_X1 U2224 ( .A1(n688), .A2(n7307), .B1(n2205), .B2(n2344), .ZN(Tvphu6)
         );
  OAI22_X1 U2225 ( .A1(n690), .A2(n6899), .B1(n2274), .B2(n2344), .ZN(X4qhu6)
         );
  OAI22_X1 U2226 ( .A1(n739), .A2(n6810), .B1(n2205), .B2(n737), .ZN(Fvphu6)
         );
  OAI22_X1 U2227 ( .A1(n738), .A2(n6678), .B1(n2274), .B2(n2253), .ZN(J4qhu6)
         );
  OAI22_X1 U2228 ( .A1(n739), .A2(n6668), .B1(n2327), .B2(n2253), .ZN(Nbshu6)
         );
  OAI22_X1 U2229 ( .A1(n738), .A2(n6663), .B1(n2323), .B2(n2253), .ZN(Ndqhu6)
         );
  OAI22_X1 U2230 ( .A1(n739), .A2(n6650), .B1(n2284), .B2(n2253), .ZN(Nxrhu6)
         );
  OAI22_X1 U2231 ( .A1(n739), .A2(n6626), .B1(n2311), .B2(n737), .ZN(Ulphu6)
         );
  OAI22_X1 U2232 ( .A1(n739), .A2(n6607), .B1(n2340), .B2(n737), .ZN(Uzphu6)
         );
  OAI22_X1 U2233 ( .A1(n739), .A2(n6603), .B1(n2331), .B2(n737), .ZN(Y8qhu6)
         );
  OAI22_X1 U2234 ( .A1(n779), .A2(n6595), .B1(n2331), .B2(n2210), .ZN(Cbqhu6)
         );
  OAI22_X1 U2235 ( .A1(n780), .A2(n6574), .B1(n2205), .B2(n776), .ZN(Jxphu6)
         );
  OAI22_X1 U2236 ( .A1(n779), .A2(n6571), .B1(n2327), .B2(n776), .ZN(Kdshu6)
         );
  OAI22_X1 U2237 ( .A1(n779), .A2(n6560), .B1(n2284), .B2(n776), .ZN(Kzrhu6)
         );
  OAI22_X1 U2238 ( .A1(n779), .A2(n6526), .B1(n2274), .B2(n776), .ZN(N6qhu6)
         );
  OAI22_X1 U2239 ( .A1(n780), .A2(n6484), .B1(n2323), .B2(n2210), .ZN(Rfqhu6)
         );
  OAI22_X1 U2240 ( .A1(n780), .A2(n6425), .B1(n2340), .B2(n2210), .ZN(Y1qhu6)
         );
  OAI22_X1 U2241 ( .A1(n779), .A2(n6399), .B1(n2311), .B2(n2210), .ZN(Ynphu6)
         );
  OAI22_X1 U2242 ( .A1(n779), .A2(n6395), .B1(n2278), .B2(n2210), .ZN(Z3shu6)
         );
  OAI22_X1 U2243 ( .A1(n709), .A2(n6267), .B1(n2205), .B2(n2289), .ZN(Eyphu6)
         );
  OAI22_X1 U2244 ( .A1(n706), .A2(n6266), .B1(n2284), .B2(n2289), .ZN(F0shu6)
         );
  OAI22_X1 U2245 ( .A1(n709), .A2(n6264), .B1(n2327), .B2(n704), .ZN(Feshu6)
         );
  OAI22_X1 U2246 ( .A1(n706), .A2(n6242), .B1(n2274), .B2(n2289), .ZN(I7qhu6)
         );
  OAI22_X1 U2247 ( .A1(n706), .A2(n6225), .B1(n2323), .B2(n2289), .ZN(Mgqhu6)
         );
  OAI22_X1 U2248 ( .A1(n706), .A2(n6212), .B1(n2340), .B2(n2289), .ZN(T2qhu6)
         );
  OAI22_X1 U2249 ( .A1(n709), .A2(n6210), .B1(n2311), .B2(n2289), .ZN(Tophu6)
         );
  OAI22_X1 U2250 ( .A1(n706), .A2(n6202), .B1(n2278), .B2(n2289), .ZN(U4shu6)
         );
  OAI22_X1 U2251 ( .A1(n709), .A2(n6183), .B1(n2331), .B2(n2289), .ZN(Xbqhu6)
         );
  OAI22_X1 U2252 ( .A1(n685), .A2(n6148), .B1(n2284), .B2(n684), .ZN(Iyrhu6)
         );
  OAI22_X1 U2253 ( .A1(n686), .A2(n6080), .B1(n2278), .B2(n2348), .ZN(X2shu6)
         );
  OAI22_X1 U2254 ( .A1(n731), .A2(n5964), .B1(n2340), .B2(n722), .ZN(H3qhu6)
         );
  OAI22_X1 U2255 ( .A1(n403), .A2(n5963), .B1(n2311), .B2(n729), .ZN(Hpphu6)
         );
  OAI22_X1 U2256 ( .A1(n403), .A2(n5961), .B1(n2278), .B2(n729), .ZN(I5shu6)
         );
  OAI22_X1 U2257 ( .A1(n403), .A2(n5956), .B1(n2331), .B2(n729), .ZN(Lcqhu6)
         );
  OAI22_X1 U2258 ( .A1(n403), .A2(n5938), .B1(n2205), .B2(n722), .ZN(Syphu6)
         );
  OAI22_X1 U2259 ( .A1(n403), .A2(n5937), .B1(n2284), .B2(n722), .ZN(T0shu6)
         );
  OAI22_X1 U2260 ( .A1(n403), .A2(n5935), .B1(n2327), .B2(n722), .ZN(Teshu6)
         );
  OAI22_X1 U2261 ( .A1(n403), .A2(n5915), .B1(n2274), .B2(n722), .ZN(W7qhu6)
         );
  OAI22_X1 U2262 ( .A1(n775), .A2(n5895), .B1(n2278), .B2(n2214), .ZN(D6shu6)
         );
  OAI22_X1 U2263 ( .A1(n775), .A2(n5873), .B1(n2284), .B2(n2214), .ZN(O1shu6)
         );
  OAI22_X1 U2264 ( .A1(n749), .A2(n5802), .B1(n2340), .B2(n2237), .ZN(F2qhu6)
         );
  OAI22_X1 U2265 ( .A1(n749), .A2(n5799), .B1(n2311), .B2(n747), .ZN(Fophu6)
         );
  OAI22_X1 U2266 ( .A1(n749), .A2(n5794), .B1(n2278), .B2(n2237), .ZN(G4shu6)
         );
  OAI22_X1 U2267 ( .A1(n749), .A2(n5752), .B1(n2331), .B2(n2237), .ZN(Jbqhu6)
         );
  OAI22_X1 U2268 ( .A1(n749), .A2(n5718), .B1(n2205), .B2(n2237), .ZN(Qxphu6)
         );
  OAI22_X1 U2269 ( .A1(n749), .A2(n5711), .B1(n2327), .B2(n2237), .ZN(Rdshu6)
         );
  OAI22_X1 U2270 ( .A1(n748), .A2(n5689), .B1(n2284), .B2(n2237), .ZN(Rzrhu6)
         );
  OAI22_X1 U2271 ( .A1(n748), .A2(n5683), .B1(n2274), .B2(n2237), .ZN(U6qhu6)
         );
  OAI22_X1 U2272 ( .A1(n749), .A2(n5662), .B1(n2323), .B2(n2237), .ZN(Yfqhu6)
         );
  OAI22_X1 U2273 ( .A1(n694), .A2(n5606), .B1(n2340), .B2(n691), .ZN(B0qhu6)
         );
  OAI22_X1 U2274 ( .A1(n694), .A2(n5598), .B1(n2311), .B2(n2315), .ZN(Bmphu6)
         );
  OAI22_X1 U2275 ( .A1(n694), .A2(n5584), .B1(n2331), .B2(n691), .ZN(F9qhu6)
         );
  OAI22_X1 U2276 ( .A1(n695), .A2(n5556), .B1(n2278), .B2(n691), .ZN(J2shu6)
         );
  OAI22_X1 U2277 ( .A1(n694), .A2(n5534), .B1(n2205), .B2(n691), .ZN(Mvphu6)
         );
  OAI22_X1 U2278 ( .A1(n695), .A2(n5526), .B1(n2274), .B2(n691), .ZN(Q4qhu6)
         );
  OAI22_X1 U2279 ( .A1(n694), .A2(n5520), .B1(n2327), .B2(n2315), .ZN(Ubshu6)
         );
  OAI22_X1 U2280 ( .A1(n695), .A2(n5507), .B1(n2323), .B2(n2315), .ZN(Udqhu6)
         );
  OAI22_X1 U2281 ( .A1(n694), .A2(n5493), .B1(n2284), .B2(n2315), .ZN(Uxrhu6)
         );
  OAI22_X1 U2282 ( .A1(n744), .A2(n5463), .B1(n2205), .B2(n2249), .ZN(Cxphu6)
         );
  OAI22_X1 U2283 ( .A1(n744), .A2(n5462), .B1(n2327), .B2(n2249), .ZN(Ddshu6)
         );
  OAI22_X1 U2284 ( .A1(n744), .A2(n5451), .B1(n2284), .B2(n740), .ZN(Dzrhu6)
         );
  OAI22_X1 U2285 ( .A1(n744), .A2(n5449), .B1(n2274), .B2(n2249), .ZN(G6qhu6)
         );
  OAI22_X1 U2286 ( .A1(n744), .A2(n5410), .B1(n2323), .B2(n2249), .ZN(Kfqhu6)
         );
  OAI22_X1 U2287 ( .A1(n744), .A2(n5372), .B1(n2340), .B2(n2249), .ZN(R1qhu6)
         );
  OAI22_X1 U2288 ( .A1(n744), .A2(n5370), .B1(n2311), .B2(n2249), .ZN(Rnphu6)
         );
  OAI22_X1 U2289 ( .A1(n744), .A2(n5369), .B1(n2278), .B2(n2249), .ZN(S3shu6)
         );
  OAI22_X1 U2290 ( .A1(n744), .A2(n5334), .B1(n2331), .B2(n2249), .ZN(Vaqhu6)
         );
  OAI22_X1 U2291 ( .A1(n399), .A2(n4181), .B1(n2327), .B2(n784), .ZN(Afshu6)
         );
  OAI22_X1 U2292 ( .A1(n714), .A2(n4179), .B1(n2274), .B2(n2285), .ZN(B7qhu6)
         );
  OAI22_X1 U2293 ( .A1(n787), .A2(n4178), .B1(n2274), .B2(n783), .ZN(D8qhu6)
         );
  OAI22_X1 U2294 ( .A1(n690), .A2(n4170), .B1(n2323), .B2(n2344), .ZN(Beqhu6)
         );
  OAI22_X1 U2295 ( .A1(n399), .A2(n4167), .B1(n2323), .B2(n784), .ZN(Hhqhu6)
         );
  OAI22_X1 U2296 ( .A1(n739), .A2(n4070), .B1(n2278), .B2(n2253), .ZN(C2shu6)
         );
  OAI22_X1 U2297 ( .A1(n787), .A2(n4066), .B1(n2278), .B2(n783), .ZN(P5shu6)
         );
  OAI22_X1 U2298 ( .A1(n399), .A2(n4007), .B1(n2311), .B2(n784), .ZN(Opphu6)
         );
  OAI22_X1 U2299 ( .A1(n787), .A2(n3611), .B1(n2205), .B2(n783), .ZN(Zyphu6)
         );
  OAI22_X1 U2300 ( .A1(n690), .A2(n3607), .B1(n2284), .B2(n2344), .ZN(Byrhu6)
         );
  OAI22_X1 U2301 ( .A1(n787), .A2(n3604), .B1(n2284), .B2(n783), .ZN(A1shu6)
         );
  OAI22_X1 U2302 ( .A1(n399), .A2(n3591), .B1(n2340), .B2(n784), .ZN(O3qhu6)
         );
  OAI22_X1 U2303 ( .A1(n787), .A2(n3588), .B1(n2331), .B2(n783), .ZN(Scqhu6)
         );
  NAND2_X1 U2304 ( .A1(n5864), .A2(n5798), .ZN(n2426) );
  NAND2_X1 U2305 ( .A1(n5869), .A2(n5243), .ZN(n3958) );
  NAND2_X1 U2306 ( .A1(n5863), .A2(n5798), .ZN(n2685) );
  NAND2_X1 U2307 ( .A1(n5870), .A2(n5243), .ZN(n3677) );
  NAND2_X1 U2308 ( .A1(n5868), .A2(n5243), .ZN(n3644) );
  NAND2_X1 U2309 ( .A1(n5863), .A2(n5255), .ZN(n2800) );
  NAND2_X1 U2310 ( .A1(n5870), .A2(n5255), .ZN(n2824) );
  NAND2_X1 U2311 ( .A1(n5870), .A2(n5867), .ZN(n3612) );
  NAND2_X1 U2312 ( .A1(n2562), .A2(n1454), .ZN(n3723) );
  NOR2_X1 U2313 ( .A1(n4426), .A2(n4166), .ZN(n5694) );
  NAND2_X1 U2314 ( .A1(n5798), .A2(n5244), .ZN(n455) );
  NAND2_X1 U2315 ( .A1(n5798), .A2(n5861), .ZN(n3597) );
  NAND2_X1 U2316 ( .A1(n5798), .A2(n5869), .ZN(n2536) );
  OAI22_X1 U2317 ( .A1(n4875), .A2(n8186), .B1(n4876), .B2(n8192), .ZN(n4918)
         );
  OAI22_X1 U2318 ( .A1(n4870), .A2(n6871), .B1(n577), .B2(n6380), .ZN(n5620)
         );
  OAI22_X1 U2319 ( .A1(n4870), .A2(n7644), .B1(n577), .B2(n6352), .ZN(n5009)
         );
  OAI22_X1 U2320 ( .A1(n4870), .A2(n8215), .B1(n4871), .B2(n8212), .ZN(n5000)
         );
  OAI22_X1 U2321 ( .A1(n4870), .A2(n7261), .B1(n4871), .B2(n6280), .ZN(n4985)
         );
  OAI22_X1 U2322 ( .A1(n4870), .A2(n7580), .B1(n577), .B2(n6330), .ZN(n5085)
         );
  OAI22_X1 U2323 ( .A1(n2321), .A2(n2231), .B1(n755), .B2(n8267), .ZN(Rgphu6)
         );
  OAI22_X1 U2324 ( .A1(n2239), .A2(n2231), .B1(n755), .B2(n6349), .ZN(Igvhu6)
         );
  OAI22_X1 U2325 ( .A1(n2399), .A2(n751), .B1(n755), .B2(n4273), .ZN(B9vhu6)
         );
  NAND2_X1 U2326 ( .A1(n5798), .A2(n5878), .ZN(n4013) );
  NAND3_X1 U2327 ( .A1(n4417), .A2(n4418), .A3(n4419), .ZN(n3410) );
  NAND3_X1 U2328 ( .A1(n3813), .A2(n2745), .A3(N3epw6), .ZN(n4418) );
  AOI22_X1 U2329 ( .A1(n2551), .A2(n4425), .B1(Nxkbx6[19]), .B2(n438), .ZN(
        n4417) );
  AOI211_X1 U2330 ( .C1(n2282), .C2(n4421), .A(Affpw6[18]), .B(n632), .ZN(
        n4419) );
  OAI22_X1 U2331 ( .A1(n6001), .A2(n5725), .B1(n6002), .B2(n6826), .ZN(n6058)
         );
  OAI22_X1 U2333 ( .A1(n6001), .A2(n5789), .B1(n6002), .B2(n3783), .ZN(n6046)
         );
  OAI22_X1 U2334 ( .A1(n6001), .A2(n8217), .B1(n6002), .B2(n8207), .ZN(n6050)
         );
  OAI22_X1 U2335 ( .A1(n6001), .A2(n5654), .B1(n6002), .B2(n6646), .ZN(n6054)
         );
  OAI22_X1 U2336 ( .A1(n6222), .A2(n3118), .B1(n6231), .B2(n6226), .ZN(n6230)
         );
  OAI22_X1 U2337 ( .A1(n6001), .A2(n5794), .B1(n6002), .B2(n4070), .ZN(n6067)
         );
  OAI22_X1 U2338 ( .A1(n6001), .A2(n5689), .B1(n6002), .B2(n6650), .ZN(n6063)
         );
  OAI22_X1 U2339 ( .A1(n6001), .A2(n5709), .B1(n6002), .B2(n6771), .ZN(n6417)
         );
  OAI22_X1 U2340 ( .A1(n6001), .A2(n8190), .B1(n6002), .B2(n8180), .ZN(n6421)
         );
  OAI22_X1 U2341 ( .A1(n6001), .A2(n5676), .B1(n6002), .B2(n6669), .ZN(n6409)
         );
  OAI22_X1 U2342 ( .A1(n6001), .A2(n5736), .B1(n6002), .B2(n6599), .ZN(n6071)
         );
  OAI22_X1 U2343 ( .A1(n6001), .A2(n5810), .B1(n6002), .B2(n6636), .ZN(n6413)
         );
  OAI22_X1 U2344 ( .A1(n6001), .A2(n5669), .B1(n6002), .B2(n6639), .ZN(n6075)
         );
  NAND2_X1 U2345 ( .A1(n5867), .A2(n5864), .ZN(n5838) );
  NOR2_X1 U2346 ( .A1(n5070), .A2(n1706), .ZN(n5648) );
  OAI22_X1 U2347 ( .A1(n6285), .A2(n3664), .B1(n6262), .B2(n3666), .ZN(n6293)
         );
  INV_X1 U2348 ( .A(n6286), .ZN(n3664) );
  NAND2_X1 U2349 ( .A1(n5878), .A2(n5243), .ZN(n4039) );
  INV_X1 U2350 ( .A(n5986), .ZN(n2437) );
  INV_X1 U2351 ( .A(n5983), .ZN(n2390) );
  NAND2_X1 U2352 ( .A1(n5861), .A2(n5255), .ZN(n3624) );
  NAND2_X1 U2353 ( .A1(n5868), .A2(n5798), .ZN(n3649) );
  NAND2_X1 U2354 ( .A1(n5869), .A2(n5255), .ZN(n4472) );
  AND3_X1 U2355 ( .A1(n5105), .A2(n5126), .A3(n5880), .ZN(n5244) );
  INV_X1 U2356 ( .A(n6216), .ZN(n4437) );
  NAND2_X1 U2357 ( .A1(n5889), .A2(n5798), .ZN(n3542) );
  INV_X1 U2358 ( .A(n5445), .ZN(n2438) );
  AOI22_X1 U2359 ( .A1(n3986), .A2(n8244), .B1(n3934), .B2(n4467), .ZN(n5893)
         );
  NAND2_X1 U2360 ( .A1(n5255), .A2(n5878), .ZN(n3579) );
  OAI21_X1 U2361 ( .B1(n6301), .B2(n6360), .A(n6361), .ZN(n6115) );
  NAND3_X1 U2362 ( .A1(n6362), .A2(n6363), .A3(n3019), .ZN(n6361) );
  AOI22_X1 U2363 ( .A1(n6364), .A2(n6181), .B1(n3018), .B2(n3635), .ZN(n6360)
         );
  AOI21_X1 U2364 ( .B1(n6316), .B2(n6366), .A(n6187), .ZN(n6364) );
  AND2_X1 U2365 ( .A1(Ntkbx6[27]), .A2(n2962), .ZN(Ovihu6) );
  OAI22_X1 U2366 ( .A1(n701), .A2(n1582), .B1(n696), .B2(n3871), .ZN(n2962) );
  INV_X1 U2367 ( .A(n1430), .ZN(n2511) );
  OAI22_X1 U2368 ( .A1(n1525), .A2(n3008), .B1(n4056), .B2(n4057), .ZN(E5xhu6)
         );
  INV_X1 U2369 ( .A(n4057), .ZN(n1525) );
  NAND2_X1 U2370 ( .A1(N701), .A2(n4058), .ZN(n4057) );
  NAND4_X1 U2371 ( .A1(n4056), .A2(n4059), .A3(n2446), .A4(n1436), .ZN(n4058)
         );
  AND2_X1 U2372 ( .A1(Ntkbx6[28]), .A2(n2405), .ZN(Wwihu6) );
  OAI22_X1 U2373 ( .A1(n697), .A2(n1580), .B1(n4110), .B2(n2297), .ZN(n2405)
         );
  AND2_X1 U2374 ( .A1(n5879), .A2(n5880), .ZN(n5868) );
  NAND3_X1 U2375 ( .A1(n4595), .A2(n4596), .A3(n4597), .ZN(n3401) );
  NAND3_X1 U2376 ( .A1(n3809), .A2(n2745), .A3(I4epw6), .ZN(n4596) );
  AOI22_X1 U2377 ( .A1(n2551), .A2(n4603), .B1(Nxkbx6[22]), .B2(n438), .ZN(
        n4595) );
  AOI211_X1 U2378 ( .C1(n2286), .C2(n4599), .A(Affpw6[21]), .B(n632), .ZN(
        n4597) );
  NAND3_X1 U2379 ( .A1(n5603), .A2(n5604), .A3(n5605), .ZN(n3393) );
  NAND3_X1 U2380 ( .A1(n3812), .A2(n2745), .A3(U3epw6), .ZN(n5604) );
  AOI22_X1 U2381 ( .A1(n2551), .A2(n4988), .B1(Nxkbx6[20]), .B2(n438), .ZN(
        n5603) );
  AOI211_X1 U2382 ( .C1(n2317), .C2(n5607), .A(Affpw6[19]), .B(n632), .ZN(
        n5605) );
  AND2_X1 U2383 ( .A1(Nvkbx6[28]), .A2(n3962), .ZN(Gglhu6) );
  OAI22_X1 U2384 ( .A1(n4110), .A2(n733), .B1(n736), .B2(n1580), .ZN(n3962) );
  AND2_X1 U2385 ( .A1(Nvkbx6[27]), .A2(n2263), .ZN(Zelhu6) );
  OAI22_X1 U2386 ( .A1(n733), .A2(n3871), .B1(n736), .B2(n1582), .ZN(n2263) );
  AND2_X1 U2387 ( .A1(Ntkbx6[29]), .A2(n4025), .ZN(Eyihu6) );
  OAI22_X1 U2388 ( .A1(n4761), .A2(n2297), .B1(n697), .B2(n1573), .ZN(n4025)
         );
  INV_X1 U2389 ( .A(n6338), .ZN(n3928) );
  NAND3_X1 U2390 ( .A1(n4655), .A2(n4656), .A3(n4657), .ZN(n3399) );
  NAND3_X1 U2391 ( .A1(n3810), .A2(n2745), .A3(B4epw6), .ZN(n4656) );
  AOI22_X1 U2392 ( .A1(n2551), .A2(n4666), .B1(Nxkbx6[21]), .B2(n438), .ZN(
        n4655) );
  AOI211_X1 U2393 ( .C1(n2290), .C2(n4659), .A(Affpw6[20]), .B(n632), .ZN(
        n4657) );
  AND2_X1 U2394 ( .A1(n5888), .A2(n5880), .ZN(n5889) );
  INV_X1 U2395 ( .A(n6132), .ZN(n3638) );
  AOI21_X1 U2396 ( .B1(n6350), .B2(n6327), .A(n6332), .ZN(n6348) );
  OAI22_X1 U2397 ( .A1(n779), .A2(n8276), .B1(n2321), .B2(n2210), .ZN(Cjphu6)
         );
  OAI22_X1 U2398 ( .A1(n695), .A2(n8274), .B1(n2321), .B2(n2315), .ZN(Fhphu6)
         );
  OAI22_X1 U2399 ( .A1(n761), .A2(n8131), .B1(n2271), .B2(n2229), .ZN(Dyshu6)
         );
  OAI22_X1 U2400 ( .A1(n768), .A2(n8074), .B1(n2399), .B2(n2218), .ZN(Bxshu6)
         );
  OAI22_X1 U2401 ( .A1(n714), .A2(n7818), .B1(n2335), .B2(n2285), .ZN(C9shu6)
         );
  OAI22_X1 U2402 ( .A1(n714), .A2(n7811), .B1(n2217), .B2(n2285), .ZN(D5thu6)
         );
  OAI22_X1 U2403 ( .A1(n714), .A2(n7809), .B1(n2399), .B2(n2285), .ZN(F6thu6)
         );
  OAI22_X1 U2404 ( .A1(n690), .A2(n7643), .B1(n2271), .B2(n687), .ZN(Dcthu6)
         );
  OAI22_X1 U2405 ( .A1(n688), .A2(n7603), .B1(n2335), .B2(n2344), .ZN(F7shu6)
         );
  OAI22_X1 U2406 ( .A1(n739), .A2(n6819), .B1(n2213), .B2(n2253), .ZN(Ftrhu6)
         );
  OAI22_X1 U2407 ( .A1(n780), .A2(n6590), .B1(n2213), .B2(n2210), .ZN(Cvrhu6)
         );
  OAI22_X1 U2408 ( .A1(n779), .A2(n6586), .B1(n2239), .B2(n2210), .ZN(E9thu6)
         );
  OAI22_X1 U2409 ( .A1(n753), .A2(n6291), .B1(n2271), .B2(n2231), .ZN(W9vhu6)
         );
  OAI22_X1 U2410 ( .A1(n748), .A2(n5789), .B1(n2271), .B2(n2237), .ZN(H7thu6)
         );
  OAI22_X1 U2411 ( .A1(n694), .A2(n5624), .B1(n2239), .B2(n2315), .ZN(Aethu6)
         );
  OAI22_X1 U2412 ( .A1(n694), .A2(n5580), .B1(n2217), .B2(n2315), .ZN(Fdthu6)
         );
  OAI22_X1 U2413 ( .A1(n743), .A2(n5464), .B1(n2399), .B2(n2249), .ZN(Bbthu6)
         );
  OAI22_X1 U2414 ( .A1(n738), .A2(n3783), .B1(n2271), .B2(n737), .ZN(Davhu6)
         );
  OAI22_X1 U2415 ( .A1(n761), .A2(n3482), .B1(n2335), .B2(n2229), .ZN(A8shu6)
         );
  OAI22_X1 U2416 ( .A1(n755), .A2(n2815), .B1(n2217), .B2(n751), .ZN(Cdvhu6)
         );
  OAI22_X1 U2417 ( .A1(n709), .A2(n2777), .B1(n2239), .B2(n2289), .ZN(A0thu6)
         );
  OAI22_X1 U2418 ( .A1(n749), .A2(n2758), .B1(n2404), .B2(n2237), .ZN(A7thu6)
         );
  INV_X1 U2419 ( .A(n5336), .ZN(n2432) );
  INV_X1 U2420 ( .A(n6145), .ZN(n3117) );
  OAI22_X1 U2421 ( .A1(n714), .A2(n7772), .B1(n2271), .B2(n2285), .ZN(R5thu6)
         );
  OAI22_X1 U2422 ( .A1(n779), .A2(n6452), .B1(n2271), .B2(n2210), .ZN(X8thu6)
         );
  OAI22_X1 U2423 ( .A1(n706), .A2(n6207), .B1(n2271), .B2(n2289), .ZN(Tzshu6)
         );
  OAI22_X1 U2424 ( .A1(n403), .A2(n5959), .B1(n2271), .B2(n729), .ZN(L2thu6)
         );
  OAI22_X1 U2425 ( .A1(n694), .A2(n5521), .B1(n2271), .B2(n2315), .ZN(Tdthu6)
         );
  OAI22_X1 U2426 ( .A1(n744), .A2(n5394), .B1(n2271), .B2(n2249), .ZN(Nathu6)
         );
  OAI22_X1 U2427 ( .A1(n399), .A2(n3781), .B1(n2271), .B2(n783), .ZN(U3thu6)
         );
  OAI22_X1 U2428 ( .A1(n749), .A2(n8272), .B1(n2321), .B2(n2237), .ZN(Jjphu6)
         );
  OAI22_X1 U2429 ( .A1(n403), .A2(n8271), .B1(n2321), .B2(n729), .ZN(Lkphu6)
         );
  OAI22_X1 U2430 ( .A1(n690), .A2(n8270), .B1(n2321), .B2(n687), .ZN(Mhphu6)
         );
  OAI22_X1 U2431 ( .A1(n760), .A2(n8269), .B1(n2321), .B2(n757), .ZN(Oiphu6)
         );
  OAI22_X1 U2432 ( .A1(n714), .A2(n8268), .B1(n2321), .B2(n712), .ZN(Qjphu6)
         );
  OAI22_X1 U2433 ( .A1(n787), .A2(n8266), .B1(n2321), .B2(n783), .ZN(Skphu6)
         );
  OAI22_X1 U2434 ( .A1(n744), .A2(n8264), .B1(n2321), .B2(n2249), .ZN(Viphu6)
         );
  OAI22_X1 U2435 ( .A1(n706), .A2(n8263), .B1(n2321), .B2(n2289), .ZN(Xjphu6)
         );
  OAI22_X1 U2436 ( .A1(n739), .A2(n8262), .B1(n2321), .B2(n737), .ZN(Ygphu6)
         );
  OAI22_X1 U2437 ( .A1(n760), .A2(n8124), .B1(n2239), .B2(n757), .ZN(Kyshu6)
         );
  OAI22_X1 U2438 ( .A1(n713), .A2(n7754), .B1(n2239), .B2(n2285), .ZN(Y5thu6)
         );
  OAI22_X1 U2439 ( .A1(n690), .A2(n7575), .B1(n2239), .B2(n687), .ZN(Kcthu6)
         );
  OAI22_X1 U2440 ( .A1(n739), .A2(n6600), .B1(n2239), .B2(n737), .ZN(Zevhu6)
         );
  OAI22_X1 U2441 ( .A1(n403), .A2(n5990), .B1(n2239), .B2(n729), .ZN(E2thu6)
         );
  OAI22_X1 U2442 ( .A1(n749), .A2(n5726), .B1(n2239), .B2(n2237), .ZN(O7thu6)
         );
  OAI22_X1 U2443 ( .A1(n743), .A2(n5348), .B1(n2239), .B2(n2249), .ZN(Uathu6)
         );
  OAI22_X1 U2444 ( .A1(n399), .A2(n3592), .B1(n2239), .B2(n784), .ZN(N3thu6)
         );
  INV_X1 U2445 ( .A(n4679), .ZN(n2328) );
  OAI22_X1 U2446 ( .A1(n761), .A2(n8117), .B1(n2399), .B2(n2229), .ZN(Ryshu6)
         );
  OAI22_X1 U2447 ( .A1(n683), .A2(n8076), .B1(n2399), .B2(n2362), .ZN(X1thu6)
         );
  OAI22_X1 U2448 ( .A1(n690), .A2(n7370), .B1(n2399), .B2(n2344), .ZN(Rcthu6)
         );
  OAI22_X1 U2449 ( .A1(n738), .A2(n6686), .B1(n2399), .B2(n2253), .ZN(I9vhu6)
         );
  OAI22_X1 U2450 ( .A1(n779), .A2(n6537), .B1(n2399), .B2(n776), .ZN(L9thu6)
         );
  OAI22_X1 U2451 ( .A1(n709), .A2(n6249), .B1(n2399), .B2(n2289), .ZN(H0thu6)
         );
  OAI22_X1 U2452 ( .A1(n686), .A2(n6138), .B1(n2399), .B2(n684), .ZN(Lvshu6)
         );
  OAI22_X1 U2453 ( .A1(n403), .A2(n5976), .B1(n2399), .B2(n722), .ZN(G3thu6)
         );
  OAI22_X1 U2454 ( .A1(n775), .A2(n5832), .B1(n2399), .B2(n2214), .ZN(Vtshu6)
         );
  OAI22_X1 U2455 ( .A1(n748), .A2(n5673), .B1(n2399), .B2(n2237), .ZN(V7thu6)
         );
  OAI22_X1 U2456 ( .A1(n694), .A2(n5562), .B1(n2399), .B2(n691), .ZN(Hethu6)
         );
  OAI22_X1 U2457 ( .A1(n399), .A2(n4272), .B1(n2399), .B2(n784), .ZN(P4thu6)
         );
  OAI22_X1 U2458 ( .A1(n760), .A2(n8118), .B1(n2217), .B2(n2229), .ZN(Pxshu6)
         );
  OAI22_X1 U2459 ( .A1(n688), .A2(n7512), .B1(n2217), .B2(n687), .ZN(Pbthu6)
         );
  OAI22_X1 U2460 ( .A1(n738), .A2(n6677), .B1(n2217), .B2(n2253), .ZN(Jdvhu6)
         );
  OAI22_X1 U2461 ( .A1(n780), .A2(n6577), .B1(n2217), .B2(n776), .ZN(J8thu6)
         );
  OAI22_X1 U2462 ( .A1(n709), .A2(n6253), .B1(n2217), .B2(n2289), .ZN(Fzshu6)
         );
  OAI22_X1 U2463 ( .A1(n403), .A2(n5898), .B1(n2217), .B2(n722), .ZN(Z2thu6)
         );
  OAI22_X1 U2465 ( .A1(n748), .A2(n5684), .B1(n2217), .B2(n2237), .ZN(T6thu6)
         );
  OAI22_X1 U2466 ( .A1(n744), .A2(n5319), .B1(n2217), .B2(n2249), .ZN(Z9thu6)
         );
  OAI22_X1 U2468 ( .A1(n787), .A2(n3593), .B1(n2217), .B2(n784), .ZN(I4thu6)
         );
  OAI22_X1 U2469 ( .A1(n761), .A2(n8108), .B1(n2404), .B2(n2229), .ZN(Wxshu6)
         );
  OAI22_X1 U2470 ( .A1(n714), .A2(n7793), .B1(n2404), .B2(n712), .ZN(K5thu6)
         );
  OAI22_X1 U2471 ( .A1(n690), .A2(n6918), .B1(n2404), .B2(n2344), .ZN(Wbthu6)
         );
  OAI22_X1 U2472 ( .A1(n739), .A2(n6605), .B1(n2404), .B2(n737), .ZN(Vcvhu6)
         );
  OAI22_X1 U2473 ( .A1(n779), .A2(n6486), .B1(n2404), .B2(n2210), .ZN(Q8thu6)
         );
  OAI22_X1 U2474 ( .A1(n709), .A2(n6221), .B1(n2404), .B2(n2289), .ZN(Mzshu6)
         );
  OAI22_X1 U2475 ( .A1(n403), .A2(n5939), .B1(n2404), .B2(n722), .ZN(S2thu6)
         );
  OAI22_X1 U2476 ( .A1(n695), .A2(n5541), .B1(n2404), .B2(n691), .ZN(Mdthu6)
         );
  OAI22_X1 U2477 ( .A1(n743), .A2(n5433), .B1(n2404), .B2(n740), .ZN(Gathu6)
         );
  OAI22_X1 U2478 ( .A1(n399), .A2(n3601), .B1(n2404), .B2(n783), .ZN(B4thu6)
         );
  OAI22_X1 U2479 ( .A1(n761), .A2(n8120), .B1(n2213), .B2(n757), .ZN(Ourhu6)
         );
  OAI22_X1 U2480 ( .A1(n714), .A2(n7775), .B1(n2213), .B2(n712), .ZN(Qvrhu6)
         );
  OAI22_X1 U2481 ( .A1(n690), .A2(n7341), .B1(n2213), .B2(n2344), .ZN(Ttrhu6)
         );
  OAI22_X1 U2483 ( .A1(n709), .A2(n6178), .B1(n2213), .B2(n2289), .ZN(Xvrhu6)
         );
  OAI22_X1 U2484 ( .A1(n403), .A2(n5955), .B1(n2213), .B2(n729), .ZN(Lwrhu6)
         );
  OAI22_X1 U2485 ( .A1(n749), .A2(n5739), .B1(n2213), .B2(n747), .ZN(Jvrhu6)
         );
  OAI22_X1 U2486 ( .A1(n694), .A2(n5540), .B1(n2213), .B2(n691), .ZN(Mtrhu6)
         );
  OAI22_X1 U2487 ( .A1(n744), .A2(n5333), .B1(n2213), .B2(n2249), .ZN(Vurhu6)
         );
  OAI22_X1 U2488 ( .A1(n787), .A2(n3587), .B1(n2213), .B2(n783), .ZN(Swrhu6)
         );
  OAI22_X1 U2489 ( .A1(n738), .A2(n6639), .B1(n2335), .B2(n2253), .ZN(R6shu6)
         );
  OAI22_X1 U2490 ( .A1(n780), .A2(n6504), .B1(n2335), .B2(n776), .ZN(O8shu6)
         );
  OAI22_X1 U2491 ( .A1(n709), .A2(n6234), .B1(n2335), .B2(n704), .ZN(J9shu6)
         );
  OAI22_X1 U2492 ( .A1(n731), .A2(n5901), .B1(n2335), .B2(n722), .ZN(X9shu6)
         );
  OAI22_X1 U2493 ( .A1(n748), .A2(n5669), .B1(n2335), .B2(n2237), .ZN(V8shu6)
         );
  OAI22_X1 U2494 ( .A1(n694), .A2(n5470), .B1(n2335), .B2(n2315), .ZN(Y6shu6)
         );
  OAI22_X1 U2495 ( .A1(n743), .A2(n5419), .B1(n2335), .B2(n740), .ZN(H8shu6)
         );
  OAI22_X1 U2496 ( .A1(n787), .A2(n3596), .B1(n2335), .B2(n784), .ZN(Eashu6)
         );
  INV_X1 U2497 ( .A(n5329), .ZN(n2442) );
  INV_X1 U2498 ( .A(n5290), .ZN(n2400) );
  INV_X1 U2499 ( .A(n5456), .ZN(n2224) );
  INV_X1 U2500 ( .A(n5695), .ZN(n2324) );
  INV_X1 U2501 ( .A(n6321), .ZN(n4432) );
  INV_X1 U2502 ( .A(n5501), .ZN(n2427) );
  INV_X1 U2503 ( .A(n5337), .ZN(n2436) );
  INV_X1 U2504 ( .A(n5472), .ZN(n2392) );
  OAI22_X1 U2505 ( .A1(n2335), .A2(n2231), .B1(n755), .B2(n6341), .ZN(K6shu6)
         );
  OAI22_X1 U2506 ( .A1(n2404), .A2(n2231), .B1(n753), .B2(n6324), .ZN(Ocvhu6)
         );
  OAI22_X1 U2507 ( .A1(n2213), .A2(n2231), .B1(n755), .B2(n6289), .ZN(Ysrhu6)
         );
  INV_X1 U2508 ( .A(n2154), .ZN(n2107) );
  OAI22_X1 U2509 ( .A1(n94), .A2(n961), .B1(n95), .B2(n8260), .ZN(n7727) );
  AOI21_X1 U2510 ( .B1(n97), .B2(n98), .A(n961), .ZN(n95) );
  AOI221_X1 U2511 ( .B1(n99), .B2(n100), .C1(n101), .C2(n102), .A(n103), .ZN(
        n94) );
  AND3_X1 U2512 ( .A1(n104), .A2(n2508), .A3(n97), .ZN(n103) );
  NAND2_X1 U2513 ( .A1(N5fpw6[2]), .A2(n667), .ZN(n4114) );
  INV_X1 U2514 ( .A(n1599), .ZN(n3113) );
  INV_X1 U2515 ( .A(n4496), .ZN(n3329) );
  OR4_X1 U2516 ( .A1(Affpw6[24]), .A2(n635), .A3(n5367), .A4(n5368), .ZN(n3412) );
  NOR3_X1 U2517 ( .A1(n3806), .A2(Qbfpw6[24]), .A3(n2549), .ZN(n5367) );
  OAI222_X1 U2518 ( .A1(n3483), .A2(n448), .B1(n2541), .B2(n5371), .C1(n4154), 
        .C2(n1608), .ZN(n5368) );
  AOI22_X1 U2519 ( .A1(n2313), .A2(n4254), .B1(n4253), .B2(n3806), .ZN(n5371)
         );
  INV_X1 U2520 ( .A(n6139), .ZN(n2809) );
  INV_X1 U2521 ( .A(n6141), .ZN(n2797) );
  INV_X1 U2522 ( .A(n6126), .ZN(n4465) );
  INV_X1 U2523 ( .A(n6135), .ZN(n3668) );
  INV_X1 U2524 ( .A(n5321), .ZN(n3062) );
  NAND2_X1 U2526 ( .A1(n8165), .A2(n8166), .ZN(n6322) );
  NAND4_X1 U2527 ( .A1(n1395), .A2(n1393), .A3(n1388), .A4(n1386), .ZN(n390)
         );
  NAND4_X1 U2528 ( .A1(n1117), .A2(n1115), .A3(n1114), .A4(n1113), .ZN(n391)
         );
  INV_X1 U2529 ( .A(n6245), .ZN(n3036) );
  INV_X1 U2530 ( .A(n6125), .ZN(n3064) );
  INV_X1 U2531 ( .A(n6233), .ZN(n3120) );
  INV_X1 U2532 ( .A(n5328), .ZN(n2419) );
  NAND3_X1 U2533 ( .A1(n2226), .A2(n4459), .A3(n5457), .ZN(n5823) );
  INV_X1 U2534 ( .A(n5324), .ZN(n2397) );
  AND3_X1 U2535 ( .A1(n2173), .A2(n2113), .A3(n5800), .ZN(n2171) );
  INV_X1 U2536 ( .A(n5297), .ZN(n2173) );
  OAI221_X1 U2538 ( .B1(n5801), .B2(n2215), .C1(n3784), .C2(n5803), .A(n5260), 
        .ZN(n5800) );
  OAI211_X1 U2539 ( .C1(n2216), .C2(n5261), .A(n5823), .B(n5262), .ZN(n5801)
         );
  INV_X1 U2540 ( .A(\eq_3147/A[0] ), .ZN(n1802) );
  INV_X1 U2541 ( .A(n6131), .ZN(n3643) );
  NAND3_X1 U2542 ( .A1(n4276), .A2(n1781), .A3(n1796), .ZN(n5809) );
  INV_X1 U2543 ( .A(n4678), .ZN(n4063) );
  INV_X1 U2544 ( .A(n4956), .ZN(n3483) );
  INV_X1 U2545 ( .A(n443), .ZN(n1808) );
  AND3_X1 U2546 ( .A1(n5151), .A2(n5152), .A3(n5153), .ZN(n3395) );
  NAND3_X1 U2547 ( .A1(n3808), .A2(n2745), .A3(n2535), .ZN(n5152) );
  AOI22_X1 U2548 ( .A1(n2551), .A2(n4941), .B1(Nxkbx6[23]), .B2(n438), .ZN(
        n5151) );
  AOI211_X1 U2549 ( .C1(n2309), .C2(n5155), .A(Affpw6[22]), .B(n632), .ZN(
        n5153) );
  NAND3_X1 U2550 ( .A1(n5649), .A2(n511), .A3(n5650), .ZN(n5637) );
  NAND4_X1 U2551 ( .A1(n5220), .A2(n1567), .A3(n493), .A4(n7375), .ZN(n5649)
         );
  NAND3_X1 U2552 ( .A1(n2562), .A2(n1626), .A3(n2563), .ZN(n5650) );
  NAND2_X1 U2553 ( .A1(n3062), .A2(n6326), .ZN(n6315) );
  AND3_X1 U2554 ( .A1(n5226), .A2(n5227), .A3(n5228), .ZN(n5199) );
  AOI221_X1 U2555 ( .B1(n492), .B2(n5232), .C1(n2562), .C2(n5233), .A(n5234), 
        .ZN(n5227) );
  NOR4_X1 U2556 ( .A1(n5229), .A2(n5230), .A3(n2575), .A4(n1661), .ZN(n5228)
         );
  AOI222_X1 U2557 ( .A1(n3189), .A2(n1663), .B1(n878), .B2(n5235), .C1(n2496), 
        .C2(n2517), .ZN(n5226) );
  OAI21_X1 U2558 ( .B1(n1537), .B2(n2104), .A(n3842), .ZN(Hyuhu6) );
  INV_X1 U2559 ( .A(HWRITE), .ZN(n2104) );
  NAND3_X1 U2560 ( .A1(n2964), .A2(n3634), .A3(n1537), .ZN(n3842) );
  OAI21_X1 U2561 ( .B1(n114), .B2(n115), .A(n3013), .ZN(n7729) );
  INV_X1 U2562 ( .A(n117), .ZN(n3013) );
  AOI21_X1 U2563 ( .B1(n119), .B2(n118), .A(N701), .ZN(n114) );
  NOR2_X1 U2564 ( .A1(n1526), .A2(n1527), .ZN(n115) );
  INV_X1 U2565 ( .A(n4800), .ZN(n3278) );
  INV_X1 U2566 ( .A(n4664), .ZN(n2440) );
  AND4_X1 U2567 ( .A1(n2974), .A2(n5790), .A3(n5791), .A4(n5792), .ZN(n742) );
  AOI221_X1 U2568 ( .B1(n2985), .B2(n8157), .C1(n2884), .C2(n4467), .A(n5925), 
        .ZN(n5791) );
  AOI221_X1 U2569 ( .B1(n2866), .B2(n8294), .C1(n2852), .C2(n8292), .A(n5926), 
        .ZN(n5790) );
  INV_X1 U2570 ( .A(n5927), .ZN(n2974) );
  OR3_X1 U2571 ( .A1(n5250), .A2(n5251), .A3(n5252), .ZN(n3721) );
  NOR4_X1 U2572 ( .A1(n492), .A2(n5263), .A3(n4688), .A4(n3723), .ZN(n5250) );
  NOR3_X1 U2573 ( .A1(n5264), .A2(n2376), .A3(n1907), .ZN(n5263) );
  INV_X1 U2574 ( .A(n6248), .ZN(n2799) );
  INV_X1 U2575 ( .A(n6231), .ZN(n4435) );
  OAI22_X1 U2576 ( .A1(n4528), .A2(n961), .B1(n4529), .B2(n2729), .ZN(Bgvhu6)
         );
  AOI21_X1 U2577 ( .B1(n97), .B2(n2507), .A(n963), .ZN(n4529) );
  AOI221_X1 U2578 ( .B1(n99), .B2(n232), .C1(n101), .C2(n4531), .A(n4532), 
        .ZN(n4528) );
  AND3_X1 U2579 ( .A1(n97), .A2(n4530), .A3(n2946), .ZN(n4532) );
  INV_X1 U2580 ( .A(n6309), .ZN(n4420) );
  INV_X1 U2581 ( .A(n6263), .ZN(n3666) );
  INV_X1 U2582 ( .A(n6335), .ZN(n4431) );
  INV_X1 U2583 ( .A(n5261), .ZN(n3784) );
  INV_X1 U2584 ( .A(n6392), .ZN(n3640) );
  INV_X1 U2585 ( .A(n6247), .ZN(n3033) );
  INV_X1 U2586 ( .A(n6337), .ZN(n3926) );
  AOI21_X1 U2587 ( .B1(n6309), .B2(n5318), .A(n6310), .ZN(n6186) );
  AND3_X1 U2588 ( .A1(n6311), .A2(n6312), .A3(n3056), .ZN(n6310) );
  NOR2_X1 U2589 ( .A1(n2611), .A2(n2643), .ZN(Tgfpw6[0]) );
  INV_X1 U2590 ( .A(n6325), .ZN(n3061) );
  OAI221_X1 U2591 ( .B1(n3925), .B2(n6312), .C1(n6307), .C2(n6305), .A(n6315), 
        .ZN(n6325) );
  INV_X1 U2592 ( .A(n2946), .ZN(n1523) );
  AND2_X1 U2593 ( .A1(Nvkbx6[29]), .A2(n3043), .ZN(Nhlhu6) );
  OAI22_X1 U2594 ( .A1(n4761), .A2(n733), .B1(n736), .B2(n1573), .ZN(n3043) );
  INV_X1 U2595 ( .A(n6223), .ZN(n2793) );
  OAI21_X1 U2596 ( .B1(n2794), .B2(n6206), .A(n6224), .ZN(n6223) );
  OAI22_X1 U2597 ( .A1(n6141), .A2(n6204), .B1(n2797), .B2(n6201), .ZN(n6224)
         );
  INV_X1 U2598 ( .A(n5819), .ZN(n2215) );
  AOI22_X1 U2599 ( .A1(n2219), .A2(n5821), .B1(n8200), .B2(n5453), .ZN(n5819)
         );
  AOI22_X1 U2600 ( .A1(n6154), .A2(n3775), .B1(n6108), .B2(n6155), .ZN(n5457)
         );
  OAI22_X1 U2601 ( .A1(n2222), .A2(n5821), .B1(n5902), .B2(n5900), .ZN(n6155)
         );
  INV_X1 U2602 ( .A(n6158), .ZN(n2222) );
  AOI21_X1 U2603 ( .B1(n5900), .B2(n5902), .A(n6159), .ZN(n6158) );
  NAND4_X1 U2604 ( .A1(n1514), .A2(n1510), .A3(n1509), .A4(n1508), .ZN(n394)
         );
  NAND4_X1 U2605 ( .A1(n1254), .A2(n1252), .A3(n1250), .A4(n1243), .ZN(n396)
         );
  AOI21_X1 U2606 ( .B1(n2149), .B2(n1351), .A(n1366), .ZN(n856) );
  NOR2_X1 U2607 ( .A1(n2262), .A2(n524), .ZN(n473) );
  NOR2_X1 U2608 ( .A1(n3549), .A2(n2124), .ZN(n1672) );
  NOR2_X1 U2609 ( .A1(n3878), .A2(n2693), .ZN(n4851) );
  NOR2_X2 U2610 ( .A1(n393), .A2(n3432), .ZN(n2299) );
  INV_X1 U2611 ( .A(n1407), .ZN(n1832) );
  OR2_X1 U2612 ( .A1(n3878), .A2(n2439), .ZN(n3874) );
  INV_X1 U2613 ( .A(n1371), .ZN(n4123) );
  NAND2_X1 U2614 ( .A1(n1144), .A2(SLEEPHOLDACKn), .ZN(n449) );
  NOR3_X1 U2615 ( .A1(n4673), .A2(n5297), .A3(n2500), .ZN(n4791) );
  NOR2_X1 U2616 ( .A1(n741), .A2(n1020), .ZN(n839) );
  NOR2_X1 U2617 ( .A1(n4635), .A2(n524), .ZN(n1685) );
  NOR2_X1 U2618 ( .A1(n5042), .A2(n270), .ZN(n1752) );
  OAI221_X1 U2619 ( .B1(n4393), .B2(n2724), .C1(n4343), .C2(n2203), .A(n5385), 
        .ZN(n269) );
  AOI221_X1 U2620 ( .B1(n4398), .B2(n4347), .C1(n4399), .C2(n4346), .A(n4349), 
        .ZN(n5385) );
  AOI221_X1 U2621 ( .B1(n4148), .B2(n4527), .C1(n4525), .C2(n4150), .A(n5150), 
        .ZN(n282) );
  OAI22_X1 U2622 ( .A1(n2724), .A2(n4522), .B1(n2710), .B2(n4523), .ZN(n5150)
         );
  NOR2_X1 U2623 ( .A1(n2233), .A2(n806), .ZN(n792) );
  NOR3_X1 U2624 ( .A1(HADDR[11]), .A2(HADDR[10]), .A3(HADDR[2]), .ZN(n163) );
  NAND3_X1 U2625 ( .A1(n2098), .A2(n3899), .A3(n911), .ZN(n741) );
  INV_X1 U2626 ( .A(n1351), .ZN(n3899) );
  OAI221_X1 U2627 ( .B1(n4522), .B2(n2703), .C1(n4523), .C2(n2723), .A(n4524), 
        .ZN(n375) );
  AOI221_X1 U2628 ( .B1(n4269), .B2(n4525), .C1(n4526), .C2(n4527), .A(n2148), 
        .ZN(n4524) );
  OAI221_X1 U2629 ( .B1(n2708), .B2(n4344), .C1(n2715), .C2(n4488), .A(n4489), 
        .ZN(n319) );
  AOI221_X1 U2630 ( .B1(n4490), .B2(n4350), .C1(n4440), .C2(n2363), .A(n2158), 
        .ZN(n4489) );
  NOR2_X1 U2631 ( .A1(n3911), .A2(n1324), .ZN(n2395) );
  OAI221_X1 U2632 ( .B1(n4143), .B2(n2724), .C1(n2138), .C2(n2710), .A(n4147), 
        .ZN(n276) );
  AOI22_X1 U2633 ( .A1(n4148), .A2(n2185), .B1(n4150), .B2(n2339), .ZN(n4147)
         );
  INV_X1 U2634 ( .A(n793), .ZN(n2164) );
  INV_X1 U2635 ( .A(n1684), .ZN(n2256) );
  OAI22_X1 U2636 ( .A1(n6285), .A2(n5303), .B1(n6286), .B2(n3659), .ZN(n6189)
         );
  OAI22_X1 U2637 ( .A1(n3300), .A2(n8245), .B1(n8231), .B2(n6275), .ZN(n6265)
         );
  OAI22_X1 U2638 ( .A1(n3292), .A2(n3867), .B1(n3293), .B2(n5306), .ZN(n6192)
         );
  INV_X1 U2640 ( .A(n6268), .ZN(n3867) );
  NAND4_X1 U2641 ( .A1(HADDR[15]), .A2(\eq_3147/A[11] ), .A3(\eq_3147/A[12] ), 
        .A4(n941), .ZN(n141) );
  NOR2_X1 U2642 ( .A1(n354), .A2(n2065), .ZN(n806) );
  AND3_X1 U2643 ( .A1(n2145), .A2(n3396), .A3(n5089), .ZN(n2318) );
  NOR3_X1 U2644 ( .A1(n635), .A2(Affpw6[5]), .A3(n2298), .ZN(n5089) );
  AOI22_X1 U2645 ( .A1(n6132), .A2(n6367), .B1(n6368), .B2(n3638), .ZN(n6181)
         );
  OAI21_X1 U2646 ( .B1(n5453), .B2(n5454), .A(n4791), .ZN(n750) );
  AOI21_X1 U2647 ( .B1(n5455), .B2(n5456), .A(n5457), .ZN(n5454) );
  NOR2_X1 U2648 ( .A1(n5309), .A2(n2792), .ZN(n5458) );
  OAI221_X1 U2649 ( .B1(n2717), .B2(n4393), .C1(n2203), .C2(n2710), .A(n5066), 
        .ZN(n312) );
  AOI22_X1 U2650 ( .A1(n4150), .A2(n4399), .B1(n4653), .B2(n4398), .ZN(n5066)
         );
  OAI221_X1 U2651 ( .B1(n2204), .B2(n2710), .C1(n2717), .C2(n4264), .A(n4754), 
        .ZN(n307) );
  AOI22_X1 U2652 ( .A1(n4653), .A2(n2351), .B1(n4150), .B2(n4270), .ZN(n4754)
         );
  OAI221_X1 U2653 ( .B1(n2717), .B2(n4638), .C1(n4632), .C2(n2721), .A(n4652), 
        .ZN(n292) );
  AOI22_X1 U2654 ( .A1(n4653), .A2(n2345), .B1(n4415), .B2(n4654), .ZN(n4652)
         );
  INV_X1 U2656 ( .A(n1482), .ZN(n3123) );
  NOR3_X1 U2657 ( .A1(n4910), .A2(n3686), .A3(n4932), .ZN(n2952) );
  OAI22_X1 U2658 ( .A1(n2276), .A2(n2231), .B1(n755), .B2(n8212), .ZN(S4rhu6)
         );
  OAI22_X1 U2659 ( .A1(n2343), .A2(n751), .B1(n755), .B2(n6380), .ZN(D0rhu6)
         );
  OAI22_X1 U2660 ( .A1(n2314), .A2(n2231), .B1(n755), .B2(n6330), .ZN(Kmqhu6)
         );
  OAI22_X1 U2661 ( .A1(n2230), .A2(n2231), .B1(n755), .B2(n6280), .ZN(Zqqhu6)
         );
  OAI221_X1 U2662 ( .B1(n3608), .B2(n4153), .C1(n4154), .C2(n1767), .A(n4737), 
        .ZN(n3429) );
  AOI221_X1 U2663 ( .B1(n2291), .B2(n4739), .C1(n4740), .C2(Qbfpw6_10), .A(
        Affpw6[10]), .ZN(n4737) );
  OAI22_X1 U2664 ( .A1(n2549), .A2(Qbfpw6_10), .B1(n2550), .B2(n4741), .ZN(
        n4739) );
  NOR2_X1 U2665 ( .A1(n4446), .A2(n2291), .ZN(n4740) );
  OAI221_X1 U2666 ( .B1(n4393), .B2(n2719), .C1(n2203), .C2(n2723), .A(n4396), 
        .ZN(n3051) );
  AOI221_X1 U2667 ( .B1(n4397), .B2(n4398), .C1(n4269), .C2(n4399), .A(n2148), 
        .ZN(n4396) );
  OAI221_X1 U2668 ( .B1(n4262), .B2(n2703), .C1(n4264), .C2(n2719), .A(n4266), 
        .ZN(n453) );
  AOI221_X1 U2669 ( .B1(n4267), .B2(n4268), .C1(n4269), .C2(n4270), .A(n2148), 
        .ZN(n4266) );
  OAI221_X1 U2670 ( .B1(n4593), .B2(n2703), .C1(n4594), .C2(n2723), .A(n5102), 
        .ZN(n379) );
  AOI221_X1 U2671 ( .B1(n4526), .B2(n2207), .C1(n4269), .C2(n4590), .A(n2148), 
        .ZN(n5102) );
  OAI221_X1 U2672 ( .B1(n4836), .B2(n2703), .C1(n4837), .C2(n2719), .A(n4838), 
        .ZN(n393) );
  AOI221_X1 U2673 ( .B1(n4267), .B2(n2398), .C1(n4269), .C2(n4840), .A(n2148), 
        .ZN(n4838) );
  OAI221_X1 U2674 ( .B1(n1786), .B2(n2513), .C1(n458), .C2(n4816), .A(n374), 
        .ZN(n7812) );
  AOI221_X1 U2675 ( .B1(n934), .B2(n375), .C1(Zsfpw6[5]), .C2(n931), .A(n213), 
        .ZN(n374) );
  OAI221_X1 U2676 ( .B1(n1783), .B2(n2513), .C1(n458), .C2(n4811), .A(n367), 
        .ZN(n7807) );
  AOI221_X1 U2677 ( .B1(n934), .B2(n368), .C1(Zsfpw6[6]), .C2(n931), .A(n213), 
        .ZN(n367) );
  OAI221_X1 U2678 ( .B1(n1775), .B2(n2513), .C1(n458), .C2(n4810), .A(n361), 
        .ZN(n7804) );
  AOI221_X1 U2679 ( .B1(n210), .B2(n362), .C1(Zsfpw6[7]), .C2(n931), .A(n213), 
        .ZN(n361) );
  OAI221_X1 U2680 ( .B1(n1767), .B2(n2513), .C1(n458), .C2(n4807), .A(n346), 
        .ZN(n7798) );
  AOI221_X1 U2681 ( .B1(n934), .B2(n347), .C1(Zsfpw6[9]), .C2(n931), .A(n213), 
        .ZN(n346) );
  OAI221_X1 U2682 ( .B1(n1764), .B2(n2513), .C1(n458), .C2(n4806), .A(n340), 
        .ZN(n7795) );
  AOI221_X1 U2683 ( .B1(n934), .B2(n341), .C1(Zsfpw6[10]), .C2(n212), .A(n213), 
        .ZN(n340) );
  OAI221_X1 U2684 ( .B1(n1719), .B2(n2513), .C1(n458), .C2(n4805), .A(n336), 
        .ZN(n7794) );
  AOI221_X1 U2685 ( .B1(n934), .B2(n337), .C1(Zsfpw6[11]), .C2(n212), .A(n213), 
        .ZN(n336) );
  OAI221_X1 U2686 ( .B1(n1717), .B2(n2513), .C1(n458), .C2(n4802), .A(n330), 
        .ZN(n7791) );
  AOI221_X1 U2687 ( .B1(n210), .B2(n331), .C1(Zsfpw6[12]), .C2(n931), .A(n213), 
        .ZN(n330) );
  OAI221_X1 U2688 ( .B1(n1696), .B2(n2513), .C1(n458), .C2(n4801), .A(n324), 
        .ZN(n7788) );
  AOI221_X1 U2689 ( .B1(n210), .B2(n325), .C1(Zsfpw6[13]), .C2(n931), .A(n213), 
        .ZN(n324) );
  OAI221_X1 U2690 ( .B1(n1604), .B2(n2513), .C1(n458), .C2(n4799), .A(n262), 
        .ZN(n7755) );
  AOI221_X1 U2691 ( .B1(n210), .B2(n263), .C1(Zsfpw6[24]), .C2(n931), .A(n213), 
        .ZN(n262) );
  OAI221_X1 U2692 ( .B1(n1597), .B2(n2513), .C1(n458), .C2(n4797), .A(n251), 
        .ZN(n7752) );
  AOI221_X1 U2693 ( .B1(n210), .B2(n252), .C1(Zsfpw6[25]), .C2(n931), .A(n213), 
        .ZN(n251) );
  OAI221_X1 U2694 ( .B1(n1804), .B2(n2513), .C1(n458), .C2(n4795), .A(n401), 
        .ZN(n7822) );
  AOI221_X1 U2695 ( .B1(n934), .B2(n402), .C1(Zsfpw6[1]), .C2(n931), .A(n213), 
        .ZN(n401) );
  OAI221_X1 U2696 ( .B1(n1801), .B2(n2513), .C1(n2569), .C2(n4787), .A(n392), 
        .ZN(n7819) );
  AOI221_X1 U2697 ( .B1(n934), .B2(n393), .C1(Zsfpw6[2]), .C2(n931), .A(n213), 
        .ZN(n392) );
  OAI221_X1 U2698 ( .B1(n1795), .B2(n2513), .C1(n2569), .C2(n4783), .A(n385), 
        .ZN(n7816) );
  AOI221_X1 U2699 ( .B1(n934), .B2(n386), .C1(Zsfpw6[3]), .C2(n931), .A(n213), 
        .ZN(n385) );
  OAI221_X1 U2700 ( .B1(n1790), .B2(n2513), .C1(n2569), .C2(n4782), .A(n378), 
        .ZN(n7813) );
  AOI221_X1 U2701 ( .B1(n934), .B2(n379), .C1(Zsfpw6[4]), .C2(n931), .A(n213), 
        .ZN(n378) );
  OAI221_X1 U2702 ( .B1(n1770), .B2(n2513), .C1(n458), .C2(n4777), .A(n357), 
        .ZN(n7803) );
  AOI221_X1 U2703 ( .B1(n934), .B2(n358), .C1(Zsfpw6[8]), .C2(n931), .A(n213), 
        .ZN(n357) );
  OAI221_X1 U2705 ( .B1(n1692), .B2(n2513), .C1(n458), .C2(n4776), .A(n318), 
        .ZN(n7785) );
  AOI221_X1 U2707 ( .B1(n210), .B2(n319), .C1(Zsfpw6[14]), .C2(n931), .A(n213), 
        .ZN(n318) );
  OAI221_X1 U2708 ( .B1(n1608), .B2(n2513), .C1(n458), .C2(n4764), .A(n268), 
        .ZN(n7758) );
  AOI221_X1 U2709 ( .B1(n210), .B2(n269), .C1(Zsfpw6[23]), .C2(n931), .A(n213), 
        .ZN(n268) );
  OAI221_X1 U2710 ( .B1(n1575), .B2(n2513), .C1(n458), .C2(n4761), .A(n231), 
        .ZN(n7743) );
  AOI221_X1 U2712 ( .B1(n210), .B2(n232), .C1(Zsfpw6[28]), .C2(n212), .A(n213), 
        .ZN(n231) );
  OAI221_X1 U2713 ( .B1(n1581), .B2(n2513), .C1(n458), .C2(n4110), .A(n238), 
        .ZN(n7746) );
  AOI221_X1 U2714 ( .B1(n210), .B2(n100), .C1(Zsfpw6[27]), .C2(n212), .A(n213), 
        .ZN(n238) );
  OAI221_X1 U2715 ( .B1(n1590), .B2(n2513), .C1(n458), .C2(n3871), .A(n245), 
        .ZN(n7749) );
  AOI221_X1 U2716 ( .B1(n210), .B2(n246), .C1(Zsfpw6[26]), .C2(n212), .A(n213), 
        .ZN(n245) );
  OAI221_X1 U2717 ( .B1(n1551), .B2(n2513), .C1(n458), .C2(n3124), .A(n223), 
        .ZN(n7741) );
  AOI221_X1 U2718 ( .B1(n210), .B2(n224), .C1(Zsfpw6[29]), .C2(n212), .A(n213), 
        .ZN(n223) );
  NAND3_X1 U2719 ( .A1(n5011), .A2(n2754), .A3(n5012), .ZN(n4047) );
  AOI22_X1 U2720 ( .A1(n2562), .A2(n2742), .B1(n228), .B2(n225), .ZN(n5012) );
  NAND3_X1 U2721 ( .A1(n266), .A2(n538), .A3(n5013), .ZN(n5011) );
  AOI22_X1 U2722 ( .A1(n3019), .A2(n6369), .B1(n6370), .B2(n6127), .ZN(n6187)
         );
  OAI221_X1 U2723 ( .B1(n4172), .B2(n442), .C1(n439), .C2(n1719), .A(n4639), 
        .ZN(n3430) );
  AOI211_X1 U2724 ( .C1(J1epw6), .C2(n4640), .A(Affpw6[12]), .B(n4641), .ZN(
        n4639) );
  NOR3_X1 U2725 ( .A1(n3819), .A2(n2549), .A3(J1epw6), .ZN(n4641) );
  OAI22_X1 U2726 ( .A1(n4446), .A2(n2287), .B1(n2550), .B2(n3819), .ZN(n4640)
         );
  OAI221_X1 U2727 ( .B1(n3337), .B2(n448), .C1(n439), .C2(n1770), .A(n4443), 
        .ZN(n3427) );
  AOI211_X1 U2728 ( .C1(Q5phu6), .C2(n4444), .A(Affpw6[9]), .B(n4445), .ZN(
        n4443) );
  OAI22_X1 U2729 ( .A1(n2550), .A2(n2326), .B1(n4446), .B2(n4447), .ZN(n4444)
         );
  NOR3_X1 U2730 ( .A1(Q5phu6), .A2(n2549), .A3(n2326), .ZN(n4445) );
  AOI22_X1 U2731 ( .A1(n5306), .A2(n3868), .B1(n6265), .B2(n3292), .ZN(n6208)
         );
  OAI221_X1 U2732 ( .B1(n2817), .B2(n448), .C1(n4154), .C2(n1764), .A(n5581), 
        .ZN(n3411) );
  AOI211_X1 U2733 ( .C1(C1epw6), .C2(n5582), .A(Affpw6[11]), .B(n5583), .ZN(
        n5581) );
  NOR3_X1 U2734 ( .A1(n3820), .A2(n2549), .A3(C1epw6), .ZN(n5583) );
  OAI22_X1 U2735 ( .A1(n4446), .A2(n2316), .B1(n2550), .B2(n3820), .ZN(n5582)
         );
  NOR2_X1 U2736 ( .A1(n6373), .A2(n6374), .ZN(n6127) );
  AOI21_X1 U2737 ( .B1(n3276), .B2(n8134), .A(n3274), .ZN(n6373) );
  AOI221_X1 U2738 ( .B1(n6375), .B2(n6371), .C1(n6363), .C2(n6362), .A(n6376), 
        .ZN(n6374) );
  AOI22_X1 U2739 ( .A1(n3020), .A2(n6370), .B1(n3021), .B2(n3272), .ZN(n6376)
         );
  OAI222_X1 U2740 ( .A1(n4858), .A2(n3587), .B1(n4859), .B2(n5955), .C1(n623), 
        .C2(n6178), .ZN(n4882) );
  OAI222_X1 U2741 ( .A1(n4858), .A2(n3593), .B1(n4859), .B2(n5898), .C1(n623), 
        .C2(n6253), .ZN(n4893) );
  OAI222_X1 U2742 ( .A1(n627), .A2(n3604), .B1(n625), .B2(n5937), .C1(n4860), 
        .C2(n6266), .ZN(n5704) );
  OAI222_X1 U2743 ( .A1(n627), .A2(n8266), .B1(n625), .B2(n8271), .C1(n4860), 
        .C2(n8263), .ZN(n5120) );
  OAI222_X1 U2744 ( .A1(n627), .A2(n3601), .B1(n625), .B2(n5939), .C1(n4860), 
        .C2(n6221), .ZN(n5437) );
  OAI221_X1 U2745 ( .B1(n4164), .B2(n448), .C1(n439), .C2(n1696), .A(n5131), 
        .ZN(n3414) );
  AOI211_X1 U2746 ( .C1(X1epw6), .C2(n5132), .A(Affpw6[14]), .B(n5133), .ZN(
        n5131) );
  NOR3_X1 U2747 ( .A1(n3817), .A2(n2549), .A3(X1epw6), .ZN(n5133) );
  OAI221_X1 U2748 ( .B1(n3040), .B2(n442), .C1(n439), .C2(n1717), .A(n5349), 
        .ZN(n3418) );
  AOI211_X1 U2749 ( .C1(Q1epw6), .C2(n5350), .A(Affpw6[13]), .B(n5351), .ZN(
        n5349) );
  NOR3_X1 U2750 ( .A1(n3818), .A2(n2549), .A3(Q1epw6), .ZN(n5351) );
  OAI22_X1 U2751 ( .A1(n4446), .A2(n2312), .B1(n2550), .B2(n3818), .ZN(n5350)
         );
  OAI21_X1 U2752 ( .B1(n3923), .B2(n4152), .A(N701), .ZN(n1364) );
  AOI211_X1 U2753 ( .C1(n3682), .C2(n475), .A(n1752), .B(n472), .ZN(n4372) );
  AND2_X1 U2754 ( .A1(n2139), .A2(n3434), .ZN(n2236) );
  AOI21_X1 U2755 ( .B1(n8150), .B2(n5192), .A(n2809), .ZN(n6211) );
  OAI22_X1 U2756 ( .A1(n6371), .A2(n6127), .B1(n3272), .B2(n3019), .ZN(n6366)
         );
  NAND2_X1 U2757 ( .A1(n792), .A2(n3289), .ZN(n798) );
  NAND4_X1 U2758 ( .A1(n450), .A2(n1977), .A3(n1430), .A4(n524), .ZN(n3289) );
  INV_X1 U2759 ( .A(n1612), .ZN(n5063) );
  OR2_X1 U2760 ( .A1(n796), .A2(n797), .ZN(n745) );
  OAI22_X1 U2761 ( .A1(n3274), .A2(n8248), .B1(n8236), .B2(n6379), .ZN(n6375)
         );
  NOR2_X1 U2762 ( .A1(n4241), .A2(n1612), .ZN(n489) );
  AOI22_X1 U2763 ( .A1(n254), .A2(n1539), .B1(n1455), .B2(n435), .ZN(n4081) );
  INV_X1 U2764 ( .A(n2375), .ZN(n2277) );
  NAND4_X1 U2765 ( .A1(n5951), .A2(n5952), .A3(n5953), .A4(n5954), .ZN(n1110)
         );
  AOI221_X1 U2766 ( .B1(n2882), .B2(n8161), .C1(n2978), .C2(n4453), .A(n5957), 
        .ZN(n5954) );
  AOI222_X1 U2767 ( .A1(n2886), .A2(n4482), .B1(n2858), .B2(n4473), .C1(n2866), 
        .C2(n5192), .ZN(n5953) );
  AOI221_X1 U2768 ( .B1(n2985), .B2(n8158), .C1(n2884), .C2(n4466), .A(n5965), 
        .ZN(n5951) );
  NAND2_X1 U2770 ( .A1(n3510), .A2(n2568), .ZN(n1571) );
  OAI22_X1 U2771 ( .A1(n760), .A2(n8130), .B1(n2269), .B2(n2229), .ZN(Ebrhu6)
         );
  OAI22_X1 U2772 ( .A1(n714), .A2(n7802), .B1(n2269), .B2(n2285), .ZN(Gcrhu6)
         );
  OAI22_X1 U2773 ( .A1(n688), .A2(n7644), .B1(n2269), .B2(n2344), .ZN(Carhu6)
         );
  OAI22_X1 U2774 ( .A1(n738), .A2(n6646), .B1(n2269), .B2(n2253), .ZN(O9rhu6)
         );
  OAI22_X1 U2775 ( .A1(n780), .A2(n6480), .B1(n2269), .B2(n2210), .ZN(Sbrhu6)
         );
  OAI22_X1 U2776 ( .A1(n755), .A2(n6352), .B1(n2269), .B2(n2231), .ZN(H9rhu6)
         );
  OAI22_X1 U2777 ( .A1(n709), .A2(n6220), .B1(n2269), .B2(n704), .ZN(Ncrhu6)
         );
  OAI22_X1 U2778 ( .A1(n749), .A2(n5654), .B1(n2269), .B2(n2237), .ZN(Zbrhu6)
         );
  OAI22_X1 U2779 ( .A1(n694), .A2(n5485), .B1(n2269), .B2(n2315), .ZN(V9rhu6)
         );
  OAI22_X1 U2780 ( .A1(n743), .A2(n5409), .B1(n2269), .B2(n2249), .ZN(Lbrhu6)
         );
  OAI22_X1 U2781 ( .A1(n403), .A2(n3653), .B1(n2269), .B2(n729), .ZN(Bdrhu6)
         );
  OAI22_X1 U2782 ( .A1(n787), .A2(n3650), .B1(n2269), .B2(n784), .ZN(Idrhu6)
         );
  OAI22_X1 U2783 ( .A1(n779), .A2(n8221), .B1(n2276), .B2(n2210), .ZN(D7rhu6)
         );
  OAI22_X1 U2784 ( .A1(n694), .A2(n8219), .B1(n2276), .B2(n2315), .ZN(G5rhu6)
         );
  OAI22_X1 U2785 ( .A1(n749), .A2(n8217), .B1(n2276), .B2(n747), .ZN(K7rhu6)
         );
  OAI22_X1 U2786 ( .A1(n403), .A2(n8216), .B1(n2276), .B2(n729), .ZN(M8rhu6)
         );
  OAI22_X1 U2787 ( .A1(n690), .A2(n8215), .B1(n2276), .B2(n2344), .ZN(N5rhu6)
         );
  OAI22_X1 U2788 ( .A1(n761), .A2(n8214), .B1(n2276), .B2(n757), .ZN(P6rhu6)
         );
  OAI22_X1 U2789 ( .A1(n714), .A2(n8213), .B1(n2276), .B2(n2285), .ZN(R7rhu6)
         );
  OAI22_X1 U2790 ( .A1(n399), .A2(n8211), .B1(n2276), .B2(n783), .ZN(T8rhu6)
         );
  OAI22_X1 U2791 ( .A1(n744), .A2(n8209), .B1(n2276), .B2(n2249), .ZN(W6rhu6)
         );
  OAI22_X1 U2792 ( .A1(n709), .A2(n8208), .B1(n2276), .B2(n2289), .ZN(Y7rhu6)
         );
  OAI22_X1 U2793 ( .A1(n739), .A2(n8207), .B1(n2276), .B2(n737), .ZN(Z4rhu6)
         );
  OAI22_X1 U2794 ( .A1(n761), .A2(n8128), .B1(n2314), .B2(n2229), .ZN(Hoqhu6)
         );
  OAI22_X1 U2795 ( .A1(n760), .A2(n8109), .B1(n2230), .B2(n2229), .ZN(Wsqhu6)
         );
  OAI22_X1 U2796 ( .A1(n714), .A2(n7821), .B1(n2343), .B2(n712), .ZN(C3rhu6)
         );
  OAI22_X1 U2797 ( .A1(n714), .A2(n7797), .B1(n2314), .B2(n2285), .ZN(Jpqhu6)
         );
  OAI22_X1 U2798 ( .A1(n714), .A2(n7745), .B1(n2230), .B2(n2285), .ZN(Ytqhu6)
         );
  OAI22_X1 U2799 ( .A1(n690), .A2(n7580), .B1(n2314), .B2(n2344), .ZN(Fnqhu6)
         );
  OAI22_X1 U2800 ( .A1(n690), .A2(n7261), .B1(n2230), .B2(n2344), .ZN(Urqhu6)
         );
  OAI22_X1 U2801 ( .A1(n690), .A2(n6871), .B1(n2343), .B2(n2344), .ZN(Y0rhu6)
         );
  OAI22_X1 U2802 ( .A1(n739), .A2(n6771), .B1(n2230), .B2(n2253), .ZN(Grqhu6)
         );
  OAI22_X1 U2803 ( .A1(n739), .A2(n6669), .B1(n2343), .B2(n2253), .ZN(K0rhu6)
         );
  OAI22_X1 U2804 ( .A1(n738), .A2(n6636), .B1(n2314), .B2(n737), .ZN(Rmqhu6)
         );
  OAI22_X1 U2805 ( .A1(n779), .A2(n6564), .B1(n2230), .B2(n776), .ZN(Ktqhu6)
         );
  OAI22_X1 U2806 ( .A1(n779), .A2(n6518), .B1(n2343), .B2(n776), .ZN(O2rhu6)
         );
  OAI22_X1 U2807 ( .A1(n780), .A2(n6478), .B1(n2314), .B2(n2210), .ZN(Voqhu6)
         );
  OAI22_X1 U2808 ( .A1(n709), .A2(n6257), .B1(n2230), .B2(n704), .ZN(Fuqhu6)
         );
  OAI22_X1 U2809 ( .A1(n709), .A2(n6239), .B1(n2343), .B2(n704), .ZN(J3rhu6)
         );
  OAI22_X1 U2810 ( .A1(n709), .A2(n6218), .B1(n2314), .B2(n704), .ZN(Qpqhu6)
         );
  OAI22_X1 U2811 ( .A1(n403), .A2(n5989), .B1(n2314), .B2(n722), .ZN(Eqqhu6)
         );
  OAI22_X1 U2812 ( .A1(n403), .A2(n5924), .B1(n2230), .B2(n722), .ZN(Tuqhu6)
         );
  OAI22_X1 U2813 ( .A1(n731), .A2(n5905), .B1(n2343), .B2(n722), .ZN(X3rhu6)
         );
  OAI22_X1 U2814 ( .A1(n749), .A2(n5810), .B1(n2314), .B2(n747), .ZN(Cpqhu6)
         );
  OAI22_X1 U2815 ( .A1(n749), .A2(n5709), .B1(n2230), .B2(n2237), .ZN(Rtqhu6)
         );
  OAI22_X1 U2816 ( .A1(n749), .A2(n5676), .B1(n2343), .B2(n2237), .ZN(V2rhu6)
         );
  OAI22_X1 U2817 ( .A1(n694), .A2(n5532), .B1(n2230), .B2(n691), .ZN(Nrqhu6)
         );
  OAI22_X1 U2818 ( .A1(n695), .A2(n5522), .B1(n2343), .B2(n2315), .ZN(R0rhu6)
         );
  OAI22_X1 U2819 ( .A1(n695), .A2(n5465), .B1(n2314), .B2(n2315), .ZN(Ymqhu6)
         );
  OAI22_X1 U2820 ( .A1(n744), .A2(n5460), .B1(n2230), .B2(n2249), .ZN(Dtqhu6)
         );
  OAI22_X1 U2821 ( .A1(n744), .A2(n5427), .B1(n2343), .B2(n740), .ZN(H2rhu6)
         );
  OAI22_X1 U2822 ( .A1(n744), .A2(n5386), .B1(n2314), .B2(n740), .ZN(Ooqhu6)
         );
  OAI22_X1 U2823 ( .A1(n399), .A2(n4003), .B1(n2314), .B2(n784), .ZN(Lqqhu6)
         );
  OAI22_X1 U2824 ( .A1(n761), .A2(n3865), .B1(n2343), .B2(n2229), .ZN(A2rhu6)
         );
  OAI22_X1 U2825 ( .A1(n787), .A2(n3864), .B1(n2343), .B2(n784), .ZN(E4rhu6)
         );
  OAI22_X1 U2826 ( .A1(n399), .A2(n3279), .B1(n2230), .B2(n784), .ZN(Avqhu6)
         );
  AOI21_X1 U2827 ( .B1(SLEEPHOLDACKn), .B2(n4674), .A(n2124), .ZN(n3510) );
  INV_X1 U2828 ( .A(n1108), .ZN(n4119) );
  NAND3_X1 U2829 ( .A1(n3211), .A2(n449), .A3(n1613), .ZN(n4241) );
  NAND2_X1 U2830 ( .A1(n5243), .A2(n5244), .ZN(n4835) );
  OAI21_X1 U2831 ( .B1(n6161), .B2(n6162), .A(n5456), .ZN(n6108) );
  NAND3_X1 U2832 ( .A1(n4475), .A2(n4476), .A3(n4477), .ZN(n3400) );
  NAND3_X1 U2833 ( .A1(n3816), .A2(n2745), .A3(L2epw6), .ZN(n4476) );
  AOI22_X1 U2834 ( .A1(n2551), .A2(n4471), .B1(Nxkbx6[16]), .B2(n438), .ZN(
        n4475) );
  AOI211_X1 U2835 ( .C1(n2283), .C2(n4479), .A(Affpw6[15]), .B(n632), .ZN(
        n4477) );
  OAI22_X1 U2836 ( .A1(n6001), .A2(n5684), .B1(n6002), .B2(n6677), .ZN(n6036)
         );
  OAI22_X1 U2837 ( .A1(n6001), .A2(n2758), .B1(n6002), .B2(n6605), .ZN(n6031)
         );
  OAI22_X1 U2838 ( .A1(n6001), .A2(n5739), .B1(n6002), .B2(n6819), .ZN(n6027)
         );
  INV_X1 U2839 ( .A(n918), .ZN(n3886) );
  AOI21_X1 U2840 ( .B1(n8292), .B2(n8294), .A(n8156), .ZN(n6261) );
  OAI22_X1 U2841 ( .A1(n6268), .A2(n3293), .B1(n6273), .B2(n6265), .ZN(n6272)
         );
  INV_X1 U2842 ( .A(n5186), .ZN(n4180) );
  OAI22_X1 U2843 ( .A1(n564), .A2(n8272), .B1(n563), .B2(n8262), .ZN(n6023) );
  INV_X1 U2844 ( .A(n4519), .ZN(n4275) );
  AOI21_X1 U2845 ( .B1(n8237), .B2(n8239), .A(n4285), .ZN(n6388) );
  AOI21_X1 U2846 ( .B1(n8240), .B2(n8250), .A(n4465), .ZN(n6345) );
  INV_X1 U2847 ( .A(n922), .ZN(n3894) );
  INV_X1 U2848 ( .A(n4488), .ZN(n2339) );
  NOR2_X1 U2849 ( .A1(n4908), .A2(n3690), .ZN(n501) );
  INV_X1 U2850 ( .A(n5286), .ZN(n2447) );
  INV_X1 U2851 ( .A(n4344), .ZN(n2185) );
  INV_X1 U2852 ( .A(n6276), .ZN(n3869) );
  NAND3_X1 U2853 ( .A1(n270), .A2(n4318), .A3(n1612), .ZN(n4373) );
  NAND2_X1 U2854 ( .A1(n3898), .A2(n443), .ZN(n2959) );
  NOR2_X1 U2855 ( .A1(n2698), .A2(n2262), .ZN(n4375) );
  NAND3_X1 U2856 ( .A1(n4792), .A2(n4793), .A3(n4794), .ZN(n3402) );
  NAND3_X1 U2857 ( .A1(n3814), .A2(n2745), .A3(G3epw6), .ZN(n4793) );
  AOI22_X1 U2858 ( .A1(n2551), .A2(n4800), .B1(Nxkbx6[18]), .B2(n438), .ZN(
        n4792) );
  AOI211_X1 U2859 ( .C1(n2320), .C2(n4796), .A(Affpw6[17]), .B(n632), .ZN(
        n4794) );
  NAND3_X1 U2860 ( .A1(n5067), .A2(n5068), .A3(n5069), .ZN(n3403) );
  NAND3_X1 U2861 ( .A1(n3815), .A2(n2745), .A3(Z2epw6), .ZN(n5068) );
  AOI22_X1 U2862 ( .A1(n2551), .A2(n4909), .B1(Nxkbx6[17]), .B2(n438), .ZN(
        n5067) );
  AOI211_X1 U2863 ( .C1(n2296), .C2(n5071), .A(Affpw6[16]), .B(n632), .ZN(
        n5069) );
  INV_X1 U2864 ( .A(n6379), .ZN(n3274) );
  OAI22_X1 U2865 ( .A1(n695), .A2(n8192), .B1(n2209), .B2(n2315), .ZN(Cwqhu6)
         );
  OAI22_X1 U2866 ( .A1(n748), .A2(n8190), .B1(n2209), .B2(n2237), .ZN(Gyqhu6)
         );
  OAI22_X1 U2867 ( .A1(n755), .A2(n8185), .B1(n2209), .B2(n2231), .ZN(Ovqhu6)
         );
  OAI22_X1 U2868 ( .A1(n761), .A2(n8129), .B1(n2236), .B2(n2229), .ZN(Eprhu6)
         );
  OAI22_X1 U2869 ( .A1(n768), .A2(n8070), .B1(n2255), .B2(n2218), .ZN(Ehshu6)
         );
  OAI22_X1 U2870 ( .A1(n714), .A2(n7815), .B1(n2318), .B2(n712), .ZN(Cnshu6)
         );
  OAI22_X1 U2871 ( .A1(n690), .A2(n7668), .B1(n2299), .B2(n2344), .ZN(Bqshu6)
         );
  OAI22_X1 U2872 ( .A1(n739), .A2(n6863), .B1(n2255), .B2(n2253), .ZN(Cgshu6)
         );
  OAI22_X1 U2873 ( .A1(n738), .A2(n6835), .B1(n2248), .B2(n2253), .ZN(Ciqhu6)
         );
  OAI22_X1 U2874 ( .A1(n738), .A2(n6826), .B1(n2325), .B2(n2253), .ZN(Derhu6)
         );
  OAI22_X1 U2875 ( .A1(n779), .A2(n6585), .B1(n2248), .B2(n2210), .ZN(Gkqhu6)
         );
  OAI22_X1 U2876 ( .A1(n753), .A2(n6378), .B1(n2288), .B2(n751), .ZN(Eevhu6)
         );
  OAI22_X1 U2877 ( .A1(n755), .A2(n6294), .B1(n2255), .B2(n2231), .ZN(Vfshu6)
         );
  OAI22_X1 U2878 ( .A1(n755), .A2(n6292), .B1(n2248), .B2(n2231), .ZN(Vhqhu6)
         );
  OAI22_X1 U2879 ( .A1(n709), .A2(n6271), .B1(n2325), .B2(n704), .ZN(Chrhu6)
         );
  OAI22_X1 U2880 ( .A1(n706), .A2(n6260), .B1(n2299), .B2(n2289), .ZN(Fsshu6)
         );
  OAI22_X1 U2881 ( .A1(n772), .A2(n5894), .B1(n2255), .B2(n2214), .ZN(Dkshu6)
         );
  OAI22_X1 U2882 ( .A1(n749), .A2(n5793), .B1(n2255), .B2(n2237), .ZN(Gishu6)
         );
  OAI22_X1 U2883 ( .A1(n744), .A2(n5461), .B1(n2299), .B2(n2249), .ZN(Drshu6)
         );
  OAI22_X1 U2884 ( .A1(n688), .A2(n4352), .B1(n2236), .B2(n687), .ZN(Corhu6)
         );
  OAI22_X1 U2885 ( .A1(n683), .A2(n4280), .B1(n2255), .B2(n2362), .ZN(Bjshu6)
         );
  OAI22_X1 U2886 ( .A1(n760), .A2(n4109), .B1(n2318), .B2(n757), .ZN(Amshu6)
         );
  OAI22_X1 U2887 ( .A1(n779), .A2(n3343), .B1(n2288), .B2(n776), .ZN(C8thu6)
         );
  OAI22_X1 U2888 ( .A1(n744), .A2(n2727), .B1(n2325), .B2(n2249), .ZN(Agrhu6)
         );
  OAI22_X1 U2889 ( .A1(n706), .A2(n2490), .B1(n2248), .B2(n2289), .ZN(Blqhu6)
         );
  INV_X1 U2890 ( .A(n5499), .ZN(n2457) );
  INV_X1 U2891 ( .A(n5489), .ZN(n2451) );
  INV_X1 U2892 ( .A(n5287), .ZN(n2207) );
  AOI221_X1 U2893 ( .B1(n3364), .B2(n4690), .C1(n853), .C2(n4705), .A(n5288), 
        .ZN(n5287) );
  OAI22_X1 U2894 ( .A1(n3106), .A2(n2388), .B1(n8316), .B2(n2713), .ZN(n5288)
         );
  OAI211_X1 U2895 ( .C1(n458), .C2(n8193), .A(n273), .B(n296), .ZN(n7773) );
  AOI222_X1 U2896 ( .A1(n275), .A2(Nxkbx6[20]), .B1(Zsfpw6[18]), .B2(n931), 
        .C1(n934), .C2(n297), .ZN(n296) );
  OAI211_X1 U2897 ( .C1(n458), .C2(n8174), .A(n273), .B(n301), .ZN(n7776) );
  AOI222_X1 U2898 ( .A1(n275), .A2(Nxkbx6[19]), .B1(Zsfpw6[17]), .B2(n931), 
        .C1(n934), .C2(n302), .ZN(n301) );
  OAI211_X1 U2899 ( .C1(n458), .C2(n4774), .A(n273), .B(n311), .ZN(n7782) );
  AOI222_X1 U2900 ( .A1(n275), .A2(Nxkbx6[17]), .B1(Zsfpw6[15]), .B2(n931), 
        .C1(n934), .C2(n312), .ZN(n311) );
  OAI211_X1 U2901 ( .C1(n458), .C2(n4773), .A(n273), .B(n306), .ZN(n7779) );
  AOI222_X1 U2902 ( .A1(n275), .A2(Nxkbx6[18]), .B1(Zsfpw6[16]), .B2(n931), 
        .C1(n934), .C2(n307), .ZN(n306) );
  OAI211_X1 U2903 ( .C1(n458), .C2(n4772), .A(n273), .B(n286), .ZN(n7767) );
  AOI222_X1 U2904 ( .A1(n275), .A2(Nxkbx6[22]), .B1(Zsfpw6[20]), .B2(n931), 
        .C1(n934), .C2(n2206), .ZN(n286) );
  OAI211_X1 U2905 ( .C1(n458), .C2(n4766), .A(n273), .B(n280), .ZN(n7764) );
  AOI222_X1 U2906 ( .A1(n275), .A2(Nxkbx6[23]), .B1(Zsfpw6[21]), .B2(n931), 
        .C1(n934), .C2(n2190), .ZN(n280) );
  INV_X1 U2907 ( .A(n282), .ZN(n2190) );
  OAI211_X1 U2908 ( .C1(n458), .C2(n4765), .A(n273), .B(n274), .ZN(n7761) );
  AOI222_X1 U2909 ( .A1(n275), .A2(Nxkbx6[24]), .B1(Zsfpw6[22]), .B2(n931), 
        .C1(n934), .C2(n276), .ZN(n274) );
  OAI211_X1 U2910 ( .C1(n458), .C2(n4184), .A(n273), .B(n291), .ZN(n7770) );
  AOI222_X1 U2911 ( .A1(n275), .A2(Nxkbx6[21]), .B1(Zsfpw6[19]), .B2(n931), 
        .C1(n210), .C2(n292), .ZN(n291) );
  OAI22_X1 U2912 ( .A1(n403), .A2(n8189), .B1(n2209), .B2(n729), .ZN(Izqhu6)
         );
  OAI22_X1 U2913 ( .A1(n690), .A2(n8188), .B1(n2209), .B2(n687), .ZN(Jwqhu6)
         );
  OAI22_X1 U2914 ( .A1(n760), .A2(n8187), .B1(n2209), .B2(n757), .ZN(Lxqhu6)
         );
  OAI22_X1 U2915 ( .A1(n714), .A2(n8186), .B1(n2209), .B2(n2285), .ZN(Nyqhu6)
         );
  OAI22_X1 U2916 ( .A1(n399), .A2(n8184), .B1(n2209), .B2(n783), .ZN(Pzqhu6)
         );
  OAI22_X1 U2917 ( .A1(n744), .A2(n8182), .B1(n2209), .B2(n2249), .ZN(Sxqhu6)
         );
  OAI22_X1 U2918 ( .A1(n706), .A2(n8181), .B1(n2209), .B2(n2289), .ZN(Uyqhu6)
         );
  OAI22_X1 U2919 ( .A1(n738), .A2(n8180), .B1(n2209), .B2(n737), .ZN(Vvqhu6)
         );
  OAI22_X1 U2920 ( .A1(n780), .A2(n8178), .B1(n2209), .B2(n2210), .ZN(Zxqhu6)
         );
  OAI22_X1 U2921 ( .A1(n760), .A2(n8110), .B1(n2299), .B2(n2229), .ZN(Wqshu6)
         );
  OAI22_X1 U2922 ( .A1(n714), .A2(n7748), .B1(n2299), .B2(n2285), .ZN(Yrshu6)
         );
  OAI22_X1 U2923 ( .A1(n738), .A2(n6657), .B1(n2299), .B2(n2253), .ZN(Npshu6)
         );
  OAI22_X1 U2924 ( .A1(n780), .A2(n6570), .B1(n2299), .B2(n776), .ZN(Krshu6)
         );
  OAI22_X1 U2925 ( .A1(n403), .A2(n5928), .B1(n2299), .B2(n722), .ZN(Tsshu6)
         );
  OAI22_X1 U2926 ( .A1(n748), .A2(n5710), .B1(n2299), .B2(n747), .ZN(Rrshu6)
         );
  OAI22_X1 U2927 ( .A1(n694), .A2(n5506), .B1(n2299), .B2(n2315), .ZN(Upshu6)
         );
  OAI22_X1 U2928 ( .A1(n399), .A2(n3774), .B1(n2299), .B2(n784), .ZN(Atshu6)
         );
  OAI22_X1 U2929 ( .A1(n755), .A2(n6351), .B1(n2236), .B2(n2231), .ZN(Hnrhu6)
         );
  OAI22_X1 U2930 ( .A1(n760), .A2(n8122), .B1(n2255), .B2(n757), .ZN(Lhshu6)
         );
  OAI22_X1 U2931 ( .A1(n761), .A2(n8115), .B1(n2248), .B2(n2229), .ZN(Sjqhu6)
         );
  OAI22_X1 U2932 ( .A1(n714), .A2(n7781), .B1(n2255), .B2(n712), .ZN(Nishu6)
         );
  OAI22_X1 U2933 ( .A1(n714), .A2(n7766), .B1(n2248), .B2(n2285), .ZN(Ukqhu6)
         );
  OAI22_X1 U2934 ( .A1(n690), .A2(n7376), .B1(n2255), .B2(n2344), .ZN(Qgshu6)
         );
  OAI22_X1 U2935 ( .A1(n690), .A2(n7372), .B1(n2248), .B2(n2344), .ZN(Qiqhu6)
         );
  OAI22_X1 U2936 ( .A1(n780), .A2(n6394), .B1(n2255), .B2(n2210), .ZN(Zhshu6)
         );
  OAI22_X1 U2937 ( .A1(n709), .A2(n6188), .B1(n2255), .B2(n2289), .ZN(Uishu6)
         );
  OAI22_X1 U2938 ( .A1(n686), .A2(n6039), .B1(n2255), .B2(n2348), .ZN(Xgshu6)
         );
  OAI22_X1 U2939 ( .A1(n403), .A2(n5960), .B1(n2255), .B2(n729), .ZN(Ijshu6)
         );
  OAI22_X1 U2940 ( .A1(n731), .A2(n5941), .B1(n2248), .B2(n729), .ZN(Plqhu6)
         );
  OAI22_X1 U2941 ( .A1(n749), .A2(n5729), .B1(n2248), .B2(n747), .ZN(Nkqhu6)
         );
  OAI22_X1 U2942 ( .A1(n695), .A2(n5555), .B1(n2255), .B2(n691), .ZN(Jgshu6)
         );
  OAI22_X1 U2943 ( .A1(n694), .A2(n5552), .B1(n2248), .B2(n691), .ZN(Jiqhu6)
         );
  OAI22_X1 U2944 ( .A1(n744), .A2(n5352), .B1(n2255), .B2(n2249), .ZN(Shshu6)
         );
  OAI22_X1 U2945 ( .A1(n744), .A2(n5317), .B1(n2248), .B2(n2249), .ZN(Zjqhu6)
         );
  OAI22_X1 U2946 ( .A1(n787), .A2(n4278), .B1(n2255), .B2(n783), .ZN(Pjshu6)
         );
  OAI22_X1 U2947 ( .A1(n787), .A2(n3583), .B1(n2248), .B2(n783), .ZN(Wlqhu6)
         );
  OAI22_X1 U2948 ( .A1(n760), .A2(n8127), .B1(n2288), .B2(n757), .ZN(Ixshu6)
         );
  OAI22_X1 U2949 ( .A1(n760), .A2(n8114), .B1(n2325), .B2(n757), .ZN(Tfrhu6)
         );
  OAI22_X1 U2950 ( .A1(n683), .A2(n8088), .B1(n2288), .B2(n2362), .ZN(O0thu6)
         );
  OAI22_X1 U2951 ( .A1(n683), .A2(n8078), .B1(n2236), .B2(n681), .ZN(Uqrhu6)
         );
  OAI22_X1 U2953 ( .A1(n767), .A2(n8055), .B1(n2288), .B2(n2218), .ZN(Svshu6)
         );
  OAI22_X1 U2954 ( .A1(n767), .A2(n7922), .B1(n2236), .B2(n2218), .ZN(Xorhu6)
         );
  OAI22_X1 U2955 ( .A1(n714), .A2(n7800), .B1(n2236), .B2(n2285), .ZN(Gqrhu6)
         );
  OAI22_X1 U2956 ( .A1(n714), .A2(n7763), .B1(n2325), .B2(n712), .ZN(Vgrhu6)
         );
  OAI22_X1 U2957 ( .A1(n714), .A2(n7760), .B1(n2288), .B2(n2285), .ZN(W4thu6)
         );
  OAI22_X1 U2958 ( .A1(n690), .A2(n7600), .B1(n2318), .B2(n687), .ZN(Flshu6)
         );
  OAI22_X1 U2959 ( .A1(n688), .A2(n7578), .B1(n2288), .B2(n2344), .ZN(Ibthu6)
         );
  OAI22_X1 U2960 ( .A1(n690), .A2(n7342), .B1(n2325), .B2(n2344), .ZN(Rerhu6)
         );
  OAI22_X1 U2961 ( .A1(n738), .A2(n6642), .B1(n2236), .B2(n2253), .ZN(Onrhu6)
         );
  OAI22_X1 U2962 ( .A1(n738), .A2(n6638), .B1(n2318), .B2(n737), .ZN(Rkshu6)
         );
  OAI22_X1 U2963 ( .A1(n739), .A2(n6628), .B1(n2288), .B2(n737), .ZN(Sevhu6)
         );
  OAI22_X1 U2964 ( .A1(n779), .A2(n6583), .B1(n2325), .B2(n776), .ZN(Hgrhu6)
         );
  OAI22_X1 U2965 ( .A1(n779), .A2(n6487), .B1(n2318), .B2(n776), .ZN(Omshu6)
         );
  OAI22_X1 U2966 ( .A1(n780), .A2(n6479), .B1(n2236), .B2(n776), .ZN(Sprhu6)
         );
  OAI22_X1 U2967 ( .A1(n706), .A2(n6229), .B1(n2318), .B2(n2289), .ZN(Jnshu6)
         );
  OAI22_X1 U2968 ( .A1(n709), .A2(n6219), .B1(n2236), .B2(n2289), .ZN(Nqrhu6)
         );
  OAI22_X1 U2969 ( .A1(n709), .A2(n6176), .B1(n2288), .B2(n2289), .ZN(Yyshu6)
         );
  OAI22_X1 U2970 ( .A1(n748), .A2(n5730), .B1(n2288), .B2(n2237), .ZN(M6thu6)
         );
  OAI22_X1 U2971 ( .A1(n749), .A2(n5725), .B1(n2325), .B2(n2237), .ZN(Ogrhu6)
         );
  OAI22_X1 U2972 ( .A1(n748), .A2(n5663), .B1(n2318), .B2(n747), .ZN(Vmshu6)
         );
  OAI22_X1 U2973 ( .A1(n749), .A2(n5642), .B1(n2236), .B2(n2237), .ZN(Zprhu6)
         );
  OAI22_X1 U2974 ( .A1(n695), .A2(n5551), .B1(n2325), .B2(n691), .ZN(Kerhu6)
         );
  OAI22_X1 U2975 ( .A1(n695), .A2(n5484), .B1(n2236), .B2(n691), .ZN(Vnrhu6)
         );
  OAI22_X1 U2976 ( .A1(n694), .A2(n5468), .B1(n2288), .B2(n2315), .ZN(Ycthu6)
         );
  OAI22_X1 U2977 ( .A1(n694), .A2(n5467), .B1(n2318), .B2(n691), .ZN(Ykshu6)
         );
  OAI22_X1 U2978 ( .A1(n744), .A2(n5411), .B1(n2318), .B2(n740), .ZN(Hmshu6)
         );
  OAI22_X1 U2979 ( .A1(n744), .A2(n5403), .B1(n2236), .B2(n2249), .ZN(Lprhu6)
         );
  OAI22_X1 U2980 ( .A1(n744), .A2(n5366), .B1(n2288), .B2(n740), .ZN(S9thu6)
         );
  OAI22_X1 U2981 ( .A1(n403), .A2(n5940), .B1(n2325), .B2(n729), .ZN(Qhrhu6)
         );
  OAI22_X1 U2982 ( .A1(n731), .A2(n5899), .B1(n2318), .B2(n722), .ZN(Xnshu6)
         );
  OAI22_X1 U2983 ( .A1(n787), .A2(n4086), .B1(n2318), .B2(n784), .ZN(Eoshu6)
         );
  OAI22_X1 U2984 ( .A1(n787), .A2(n3581), .B1(n2325), .B2(n783), .ZN(Xhrhu6)
         );
  OAI22_X1 U2985 ( .A1(n802), .A2(n5236), .B1(n2163), .B2(n804), .ZN(n7871) );
  AOI21_X1 U2986 ( .B1(n3712), .B2(n805), .A(n961), .ZN(n802) );
  NAND2_X1 U2987 ( .A1(N701), .A2(n805), .ZN(n804) );
  OAI21_X1 U2988 ( .B1(n808), .B2(n3762), .A(n810), .ZN(n805) );
  OAI22_X1 U2989 ( .A1(n798), .A2(n3620), .B1(n3532), .B2(n796), .ZN(n7870) );
  INV_X1 U2990 ( .A(n801), .ZN(n3532) );
  OAI22_X1 U2991 ( .A1(n3486), .A2(n3044), .B1(n2514), .B2(n3046), .ZN(Nfvhu6)
         );
  INV_X1 U2992 ( .A(n3044), .ZN(n2514) );
  NAND2_X1 U2993 ( .A1(n3052), .A2(n3053), .ZN(n3044) );
  AOI22_X1 U2994 ( .A1(n1815), .A2(n3066), .B1(n3049), .B2(n3484), .ZN(n3046)
         );
  NAND4_X1 U2995 ( .A1(n845), .A2(n846), .A3(n2026), .A4(n2033), .ZN(n7875) );
  AOI221_X1 U2996 ( .B1(n239), .B2(n4145), .C1(n856), .C2(n3042), .A(n858), 
        .ZN(n845) );
  INV_X1 U2997 ( .A(n852), .ZN(n2026) );
  INV_X1 U2998 ( .A(n849), .ZN(n2033) );
  INV_X1 U2999 ( .A(n5400), .ZN(n2203) );
  OAI222_X1 U3000 ( .A1(n3314), .A2(n5387), .B1(n2713), .B2(n8314), .C1(n874), 
        .C2(n2712), .ZN(n5400) );
  INV_X1 U3001 ( .A(n5498), .ZN(n2456) );
  OAI22_X1 U3002 ( .A1(n2299), .A2(n751), .B1(n755), .B2(n6365), .ZN(Gpshu6)
         );
  OAI22_X1 U3003 ( .A1(n2318), .A2(n2231), .B1(n753), .B2(n6331), .ZN(Kkshu6)
         );
  OAI22_X1 U3004 ( .A1(n2325), .A2(n2231), .B1(n753), .B2(n6290), .ZN(Wdrhu6)
         );
  INV_X1 U3005 ( .A(n6362), .ZN(n3024) );
  INV_X1 U3006 ( .A(n5306), .ZN(n3292) );
  OAI21_X1 U3007 ( .B1(n158), .B2(n159), .A(n316), .ZN(n154) );
  AND4_X1 U3008 ( .A1(n1772), .A2(HADDR[9]), .A3(n163), .A4(n164), .ZN(n158)
         );
  AOI21_X1 U3009 ( .B1(n161), .B2(n162), .A(HADDR[9]), .ZN(n159) );
  NAND3_X1 U3010 ( .A1(n163), .A2(HADDR[8]), .A3(n164), .ZN(n162) );
  NAND2_X1 U3011 ( .A1(n2585), .A2(n4987), .ZN(n4318) );
  INV_X1 U3012 ( .A(n6130), .ZN(n4285) );
  INV_X1 U3013 ( .A(n6137), .ZN(n8156) );
  NAND4_X1 U3015 ( .A1(n1999), .A2(n1116), .A3(n2020), .A4(n1118), .ZN(n7899)
         );
  INV_X1 U3016 ( .A(n1129), .ZN(n1999) );
  AOI221_X1 U3017 ( .B1(n876), .B2(LOCKUP), .C1(n884), .C2(Gqgpw6[19]), .A(
        n1120), .ZN(n1118) );
  INV_X1 U3018 ( .A(n1121), .ZN(n2020) );
  INV_X1 U3019 ( .A(n6275), .ZN(n3300) );
  NAND2_X1 U3020 ( .A1(n5210), .A2(n8144), .ZN(n6363) );
  NAND2_X1 U3021 ( .A1(n165), .A2(n1779), .ZN(n161) );
  INV_X1 U3022 ( .A(HADDR[7]), .ZN(n1779) );
  OAI21_X1 U3023 ( .B1(HADDR[2]), .B2(n365), .A(HADDR[11]), .ZN(n167) );
  INV_X1 U3024 ( .A(n1613), .ZN(n2251) );
  INV_X1 U3025 ( .A(n4268), .ZN(n2204) );
  INV_X1 U3026 ( .A(n102), .ZN(n4376) );
  INV_X1 U3027 ( .A(n4531), .ZN(n3032) );
  INV_X1 U3028 ( .A(n171), .ZN(n1726) );
  OAI21_X1 U3029 ( .B1(HADDR[2]), .B2(HADDR[3]), .A(HADDR[7]), .ZN(n173) );
  NAND3_X1 U3030 ( .A1(HADDR[11]), .A2(HADDR[4]), .A3(n952), .ZN(n172) );
  INV_X1 U3031 ( .A(n1566), .ZN(n4521) );
  INV_X1 U3032 ( .A(n1135), .ZN(n4118) );
  INV_X1 U3033 ( .A(n4878), .ZN(n3040) );
  INV_X1 U3034 ( .A(n4938), .ZN(n2817) );
  INV_X1 U3035 ( .A(n4888), .ZN(n4164) );
  INV_X1 U3036 ( .A(n4649), .ZN(n4172) );
  INV_X1 U3038 ( .A(n4449), .ZN(n3337) );
  INV_X1 U3039 ( .A(n4955), .ZN(n4006) );
  INV_X1 U3040 ( .A(n4939), .ZN(n3602) );
  OR4_X1 U3041 ( .A1(n1726), .A2(n328), .A3(HADDR[11]), .A4(HADDR[8]), .ZN(
        n155) );
  INV_X1 U3042 ( .A(n4168), .ZN(n3780) );
  INV_X1 U3043 ( .A(n1136), .ZN(n3911) );
  NAND2_X1 U3044 ( .A1(n8143), .A2(n3870), .ZN(n6277) );
  AND2_X1 U3045 ( .A1(n6388), .A2(n6132), .ZN(n6301) );
  AND2_X1 U3046 ( .A1(n6332), .A2(n5321), .ZN(n6314) );
  INV_X1 U3047 ( .A(n795), .ZN(n2181) );
  AND2_X1 U3048 ( .A1(n6345), .A2(n5321), .ZN(n6318) );
  INV_X1 U3049 ( .A(n4589), .ZN(n2206) );
  AOI221_X1 U3050 ( .B1(n4590), .B2(n4150), .C1(n4148), .C2(n2207), .A(n4592), 
        .ZN(n4589) );
  OAI22_X1 U3051 ( .A1(n2724), .A2(n4593), .B1(n2710), .B2(n4594), .ZN(n4592)
         );
  INV_X1 U3052 ( .A(n6393), .ZN(n4282) );
  INV_X1 U3053 ( .A(n6273), .ZN(n3868) );
  OR3_X1 U3054 ( .A1(n3511), .A2(n5231), .A3(n1660), .ZN(n5229) );
  INV_X1 U3055 ( .A(n3269), .ZN(n4587) );
  INV_X1 U3056 ( .A(n6371), .ZN(n3021) );
  INV_X1 U3057 ( .A(n4080), .ZN(n3767) );
  NAND2_X1 U3058 ( .A1(n796), .A2(n3281), .ZN(L0vhu6) );
  NAND4_X1 U3059 ( .A1(n2167), .A2(n2118), .A3(n1430), .A4(n2234), .ZN(n3281)
         );
  INV_X1 U3060 ( .A(n6369), .ZN(n3020) );
  NAND2_X1 U3061 ( .A1(n793), .A2(n3991), .ZN(Fivhu6) );
  OAI21_X1 U3062 ( .B1(n3992), .B2(n806), .A(n2233), .ZN(n3991) );
  AOI21_X1 U3063 ( .B1(n3565), .B2(N701), .A(n354), .ZN(n3992) );
  OAI21_X1 U3064 ( .B1(n6483), .B2(n3109), .A(n254), .ZN(n6482) );
  AOI21_X1 U3065 ( .B1(n6485), .B2(n3351), .A(n3112), .ZN(n6483) );
  INV_X1 U3066 ( .A(n6447), .ZN(n3109) );
  INV_X1 U3067 ( .A(n180), .ZN(n1851) );
  OAI22_X1 U3068 ( .A1(n3106), .A2(n2368), .B1(n8324), .B2(n2713), .ZN(n5338)
         );
  OAI21_X1 U3069 ( .B1(n3213), .B2(n3214), .A(N701), .ZN(n1694) );
  OAI211_X1 U3070 ( .C1(n4205), .C2(n426), .A(n1888), .B(n2122), .ZN(n3214) );
  OAI221_X1 U3071 ( .B1(n3218), .B2(n4608), .C1(n2262), .C2(n1923), .A(n3220), 
        .ZN(n3213) );
  INV_X1 U3072 ( .A(n3217), .ZN(n1888) );
  NAND2_X1 U3073 ( .A1(n3488), .A2(n450), .ZN(n1997) );
  AOI221_X1 U3074 ( .B1(n900), .B2(n4705), .C1(n3313), .C2(n4690), .A(n5496), 
        .ZN(n4523) );
  OAI22_X1 U3075 ( .A1(n3106), .A2(n2428), .B1(n8308), .B2(n2713), .ZN(n5496)
         );
  AOI221_X1 U3076 ( .B1(n1213), .B2(n4705), .C1(n3364), .C2(n4717), .A(n4775), 
        .ZN(n4264) );
  OAI22_X1 U3077 ( .A1(n3104), .A2(n2368), .B1(n8320), .B2(n2713), .ZN(n4775)
         );
  OAI22_X1 U3078 ( .A1(n254), .A2(n6445), .B1(n7355), .B2(n6446), .ZN(n4556)
         );
  AOI21_X1 U3079 ( .B1(n6445), .B2(n6447), .A(n4559), .ZN(n6446) );
  NAND3_X1 U3080 ( .A1(n955), .A2(N701), .A3(n3850), .ZN(n909) );
  INV_X1 U3081 ( .A(HWDATA[22]), .ZN(n2671) );
  INV_X1 U3082 ( .A(HWDATA[23]), .ZN(n2676) );
  OAI21_X1 U3083 ( .B1(n4299), .B2(n4300), .A(N701), .ZN(n1916) );
  NAND4_X1 U3084 ( .A1(n2122), .A2(n1970), .A3(n1910), .A4(n4302), .ZN(n4300)
         );
  NAND4_X1 U3085 ( .A1(n3187), .A2(n447), .A3(n4311), .A4(n4312), .ZN(n4299)
         );
  AOI222_X1 U3086 ( .A1(n496), .A2(n4303), .B1(n1588), .B2(n1674), .C1(n1488), 
        .C2(n1594), .ZN(n4302) );
  OAI222_X1 U3087 ( .A1(n2416), .A2(n5387), .B1(n1180), .B2(n2712), .C1(n2713), 
        .C2(n8306), .ZN(n4399) );
  INV_X1 U3088 ( .A(n3334), .ZN(n2416) );
  OAI222_X1 U3089 ( .A1(n2820), .A2(n2712), .B1(n3373), .B2(n5387), .C1(n2713), 
        .C2(n8329), .ZN(n4398) );
  INV_X1 U3090 ( .A(n997), .ZN(n2820) );
  AOI221_X1 U3091 ( .B1(n3326), .B2(n4717), .C1(n3323), .C2(n4690), .A(n5685), 
        .ZN(n5553) );
  OAI22_X1 U3092 ( .A1(n2712), .A2(n2827), .B1(n8311), .B2(n2713), .ZN(n5685)
         );
  AOI221_X1 U3093 ( .B1(n1343), .B2(n4705), .C1(n3379), .C2(n4690), .A(n4706), 
        .ZN(n4412) );
  OAI22_X1 U3094 ( .A1(n3106), .A2(n2358), .B1(n8327), .B2(n2713), .ZN(n4706)
         );
  INV_X1 U3095 ( .A(n119), .ZN(n3012) );
  AOI221_X1 U3096 ( .B1(n3361), .B2(n4717), .C1(n3368), .C2(n4690), .A(n5678), 
        .ZN(n4837) );
  OAI22_X1 U3097 ( .A1(n2712), .A2(n2835), .B1(n8318), .B2(n2713), .ZN(n5678)
         );
  NAND4_X1 U3098 ( .A1(n677), .A2(n689), .A3(n897), .A4(n2233), .ZN(n676) );
  NAND2_X1 U3099 ( .A1(n692), .A2(n3766), .ZN(n689) );
  AOI211_X1 U3100 ( .C1(n5313), .C2(n6534), .A(n6536), .B(n2596), .ZN(n5622)
         );
  INV_X1 U3101 ( .A(n6538), .ZN(n2596) );
  AOI22_X1 U3102 ( .A1(n6529), .A2(n3571), .B1(n6530), .B2(n5304), .ZN(n6538)
         );
  INV_X1 U3103 ( .A(n705), .ZN(n2119) );
  INV_X1 U3104 ( .A(n710), .ZN(n3259) );
  OAI221_X1 U3105 ( .B1(n2400), .B2(n3347), .C1(n2390), .C2(n3358), .A(n5444), 
        .ZN(n3322) );
  AOI22_X1 U3106 ( .A1(n629), .A2(n4664), .B1(n568), .B2(n5445), .ZN(n5444) );
  OAI222_X1 U3107 ( .A1(n439), .A2(n1795), .B1(n2700), .B2(n5105), .C1(n3956), 
        .C2(n4153), .ZN(n3394) );
  OAI221_X1 U3108 ( .B1(n2457), .B2(n387), .C1(n2427), .C2(n3358), .A(n5335), 
        .ZN(n3318) );
  AOI22_X1 U3109 ( .A1(n4734), .A2(n5336), .B1(n4763), .B2(n5337), .ZN(n5335)
         );
  OAI221_X1 U3110 ( .B1(n2406), .B2(n387), .C1(n2384), .C2(n3358), .A(n5539), 
        .ZN(n3365) );
  AOI22_X1 U3111 ( .A1(n4734), .A2(n5340), .B1(n4763), .B2(n4646), .ZN(n5539)
         );
  AOI221_X1 U3112 ( .B1(n3381), .B2(n4690), .C1(n1267), .C2(n4705), .A(n6455), 
        .ZN(n5127) );
  OAI22_X1 U3113 ( .A1(n8325), .A2(n2713), .B1(n3106), .B2(n2366), .ZN(n6455)
         );
  NOR3_X1 U3114 ( .A1(n2430), .A2(n5786), .A3(n5564), .ZN(n5558) );
  OAI221_X1 U3115 ( .B1(n2413), .B2(n3358), .C1(n2397), .C2(n459), .A(n5982), 
        .ZN(n3361) );
  AOI22_X1 U3116 ( .A1(n568), .A2(n5983), .B1(n629), .B2(n5472), .ZN(n5982) );
  OAI221_X1 U3117 ( .B1(n2419), .B2(n3358), .C1(n2427), .C2(n3347), .A(n6060), 
        .ZN(n3328) );
  AOI22_X1 U3118 ( .A1(n629), .A2(n5336), .B1(n568), .B2(n5337), .ZN(n6060) );
  INV_X1 U3119 ( .A(n711), .ZN(n2111) );
  OAI221_X1 U3120 ( .B1(n2437), .B2(n631), .C1(n2438), .C2(n459), .A(n6043), 
        .ZN(n3325) );
  AOI22_X1 U3121 ( .A1(n5280), .A2(n4664), .B1(n568), .B2(n5329), .ZN(n6043)
         );
  OAI221_X1 U3122 ( .B1(n2406), .B2(n631), .C1(n2387), .C2(n3358), .A(n5944), 
        .ZN(n3368) );
  AOI22_X1 U3123 ( .A1(n4734), .A2(n4646), .B1(n568), .B2(n5945), .ZN(n5944)
         );
  OAI221_X1 U3125 ( .B1(n2347), .B2(n631), .C1(n2355), .C2(n459), .A(n5950), 
        .ZN(n3380) );
  AOI22_X1 U3127 ( .A1(n5280), .A2(n5491), .B1(n568), .B2(n5538), .ZN(n5950)
         );
  OAI221_X1 U3128 ( .B1(n2347), .B2(n3347), .C1(n2355), .C2(n3358), .A(n6493), 
        .ZN(n3381) );
  AOI22_X1 U3129 ( .A1(n629), .A2(n5538), .B1(n568), .B2(n5342), .ZN(n6493) );
  OAI221_X1 U3130 ( .B1(n2384), .B2(n387), .C1(n2365), .C2(n3358), .A(n5942), 
        .ZN(n3382) );
  AOI22_X1 U3131 ( .A1(n4734), .A2(n5536), .B1(n4763), .B2(n5537), .ZN(n5942)
         );
  OAI221_X1 U3132 ( .B1(n2451), .B2(n3347), .C1(n2456), .C2(n3358), .A(n5285), 
        .ZN(n3339) );
  AOI22_X1 U3133 ( .A1(n568), .A2(n4390), .B1(n629), .B2(n5286), .ZN(n5285) );
  OAI221_X1 U3134 ( .B1(n2457), .B2(n3347), .C1(n2436), .C2(n3358), .A(n5929), 
        .ZN(n3340) );
  AOI22_X1 U3135 ( .A1(n568), .A2(n5489), .B1(n4763), .B2(n5498), .ZN(n5929)
         );
  NOR2_X1 U3136 ( .A1(HADDR[3]), .A2(HADDR[4]), .ZN(n164) );
  OAI221_X1 U3137 ( .B1(n2432), .B2(n387), .C1(n2442), .C2(n3358), .A(n5930), 
        .ZN(n3326) );
  AOI22_X1 U3138 ( .A1(n4734), .A2(n5328), .B1(n4763), .B2(n5501), .ZN(n5930)
         );
  OAI221_X1 U3139 ( .B1(n1021), .B2(n2712), .C1(n2713), .C2(n8312), .A(n4716), 
        .ZN(n4416) );
  AOI22_X1 U3140 ( .A1(n4717), .A2(n3313), .B1(n4690), .B2(n3322), .ZN(n4716)
         );
  OAI221_X1 U3141 ( .B1(n2840), .B2(n2712), .C1(n2713), .C2(n8310), .A(n6042), 
        .ZN(n4654) );
  AOI22_X1 U3142 ( .A1(n4717), .A2(n3328), .B1(n4690), .B2(n3325), .ZN(n6042)
         );
  OAI221_X1 U3143 ( .B1(n2413), .B2(n631), .C1(n2403), .C2(n459), .A(n5322), 
        .ZN(n3364) );
  AOI22_X1 U3144 ( .A1(n5280), .A2(n5323), .B1(n568), .B2(n5324), .ZN(n5322)
         );
  OAI221_X1 U3146 ( .B1(n2438), .B2(n631), .C1(n2400), .C2(n3358), .A(n5985), 
        .ZN(n3323) );
  AOI22_X1 U3148 ( .A1(n4734), .A2(n4664), .B1(n568), .B2(n5986), .ZN(n5985)
         );
  INV_X1 U3149 ( .A(HWDATA[17]), .ZN(n2679) );
  INV_X1 U3150 ( .A(HWDATA[19]), .ZN(n2686) );
  OAI222_X1 U3151 ( .A1(n439), .A2(n1804), .B1(n3881), .B2(n448), .C1(n243), 
        .C2(n4364), .ZN(n3424) );
  INV_X1 U3152 ( .A(HWDATA[20]), .ZN(n2689) );
  INV_X1 U3153 ( .A(HWDATA[21]), .ZN(n2691) );
  OAI221_X1 U3154 ( .B1(n2717), .B2(n4411), .C1(n4412), .C2(n2724), .A(n4413), 
        .ZN(n302) );
  AOI22_X1 U3155 ( .A1(n4150), .A2(n4414), .B1(n4415), .B2(n4416), .ZN(n4413)
         );
  AOI22_X1 U3156 ( .A1(n5070), .A2(n1520), .B1(n5771), .B2(n1642), .ZN(n4561)
         );
  NAND2_X1 U3157 ( .A1(n1419), .A2(n3282), .ZN(n1376) );
  NAND4_X1 U3158 ( .A1(n3283), .A2(n3284), .A3(n3285), .A4(n1978), .ZN(n3282)
         );
  OAI21_X1 U3159 ( .B1(n524), .B2(n963), .A(n3286), .ZN(n3284) );
  NAND3_X1 U3160 ( .A1(n1430), .A2(n2510), .A3(n1996), .ZN(n3286) );
  OAI221_X1 U3161 ( .B1(n2432), .B2(n3358), .C1(n2436), .C2(n459), .A(n5497), 
        .ZN(n3319) );
  AOI22_X1 U3162 ( .A1(n568), .A2(n5498), .B1(n4763), .B2(n5499), .ZN(n5497)
         );
  OAI221_X1 U3163 ( .B1(n2370), .B2(n3358), .C1(n2384), .C2(n459), .A(n5339), 
        .ZN(n3366) );
  AOI22_X1 U3164 ( .A1(n568), .A2(n4646), .B1(n4763), .B2(n5340), .ZN(n5339)
         );
  OAI221_X1 U3165 ( .B1(n2390), .B2(n3347), .C1(n2392), .C2(n3358), .A(n5289), 
        .ZN(n3321) );
  AOI22_X1 U3166 ( .A1(n568), .A2(n4664), .B1(n4763), .B2(n5290), .ZN(n5289)
         );
  OAI221_X1 U3167 ( .B1(n2462), .B2(n3347), .C1(n2460), .C2(n631), .A(n5279), 
        .ZN(n3378) );
  AOI22_X1 U3168 ( .A1(n5280), .A2(n5281), .B1(n568), .B2(n5283), .ZN(n5279)
         );
  AOI222_X1 U3169 ( .A1(n5316), .A2(n3019), .B1(n5318), .B2(n3015), .C1(n5320), 
        .C2(n5321), .ZN(n5315) );
  OAI221_X1 U3170 ( .B1(n2462), .B2(n3358), .C1(n2460), .C2(n459), .A(n5490), 
        .ZN(n3379) );
  AOI22_X1 U3171 ( .A1(n629), .A2(n5283), .B1(n568), .B2(n5343), .ZN(n5490) );
  AOI22_X1 U3172 ( .A1(n5294), .A2(n1520), .B1(n5019), .B2(n1642), .ZN(n6485)
         );
  NOR2_X1 U3173 ( .A1(n6498), .A2(n6503), .ZN(n4763) );
  NOR2_X1 U3174 ( .A1(n5173), .A2(n5174), .ZN(n4400) );
  NOR2_X1 U3175 ( .A1(n904), .A2(n903), .ZN(n4844) );
  INV_X1 U3176 ( .A(n220), .ZN(n1852) );
  NAND3_X1 U3177 ( .A1(HADDR[5]), .A2(HADDR[11]), .A3(n175), .ZN(n170) );
  AOI22_X1 U3178 ( .A1(HADDR[2]), .A2(n176), .B1(n316), .B2(n1791), .ZN(n175)
         );
  NAND2_X1 U3179 ( .A1(n955), .A2(n365), .ZN(n176) );
  INV_X1 U3180 ( .A(n164), .ZN(n1791) );
  NOR2_X1 U3181 ( .A1(n2595), .A2(n5194), .ZN(n4612) );
  INV_X1 U3182 ( .A(HWDATA[24]), .ZN(n2632) );
  NOR3_X1 U3183 ( .A1(n202), .A2(n961), .A3(n2154), .ZN(n2152) );
  NOR2_X1 U3184 ( .A1(n5194), .A2(n5622), .ZN(n4407) );
  AOI22_X1 U3185 ( .A1(n4206), .A2(n4207), .B1(n7374), .B2(n963), .ZN(Crohu6)
         );
  NOR4_X1 U3186 ( .A1(n4208), .A2(n4209), .A3(n4210), .A4(n4211), .ZN(n4207)
         );
  NOR4_X1 U3187 ( .A1(n4224), .A2(n4225), .A3(n1932), .A4(n2904), .ZN(n4206)
         );
  AOI22_X1 U3188 ( .A1(n3785), .A2(n6154), .B1(n4454), .B2(n2226), .ZN(n5900)
         );
  OAI221_X1 U3189 ( .B1(n2458), .B2(n3347), .C1(n2459), .C2(n3358), .A(n5995), 
        .ZN(n5395) );
  AOI22_X1 U3190 ( .A1(n568), .A2(n5491), .B1(n4763), .B2(n5492), .ZN(n5995)
         );
  OAI221_X1 U3191 ( .B1(n4836), .B2(n2724), .C1(n2721), .C2(n2435), .A(n5599), 
        .ZN(n297) );
  AOI22_X1 U3192 ( .A1(n4148), .A2(n2385), .B1(n4415), .B2(n2398), .ZN(n5599)
         );
  NOR3_X1 U3193 ( .A1(n398), .A2(n1886), .A3(n1887), .ZN(n1861) );
  OAI221_X1 U3194 ( .B1(n2459), .B2(n3347), .C1(n2447), .C2(n3358), .A(n5949), 
        .ZN(n5674) );
  AOI22_X1 U3195 ( .A1(n568), .A2(n5492), .B1(n4763), .B2(n5281), .ZN(n5949)
         );
  OAI221_X1 U3196 ( .B1(n2403), .B2(n631), .C1(n2406), .C2(n459), .A(n6084), 
        .ZN(n3367) );
  AOI22_X1 U3197 ( .A1(n5280), .A2(n4646), .B1(n568), .B2(n5984), .ZN(n6084)
         );
  OAI221_X1 U3198 ( .B1(n4006), .B2(n442), .C1(n439), .C2(n1775), .A(n5044), 
        .ZN(n3415) );
  AOI211_X1 U3199 ( .C1(W4epw6), .C2(n5045), .A(Affpw6[8]), .B(n5046), .ZN(
        n5044) );
  NOR3_X1 U3200 ( .A1(n3791), .A2(n2549), .A3(W4epw6), .ZN(n5046) );
  OAI22_X1 U3201 ( .A1(n4446), .A2(n2294), .B1(n2550), .B2(n3791), .ZN(n5045)
         );
  OAI221_X1 U3202 ( .B1(n2367), .B2(n3358), .C1(n2370), .C2(n3347), .A(n6456), 
        .ZN(n3383) );
  AOI22_X1 U3203 ( .A1(n629), .A2(n5943), .B1(n568), .B2(n5340), .ZN(n6456) );
  OAI221_X1 U3204 ( .B1(n2451), .B2(n631), .C1(n2456), .C2(n459), .A(n6020), 
        .ZN(n5393) );
  AOI22_X1 U3205 ( .A1(n5280), .A2(n5499), .B1(n568), .B2(n5286), .ZN(n6020)
         );
  OAI221_X1 U3206 ( .B1(n2413), .B2(n3347), .C1(n2403), .C2(n3358), .A(n5471), 
        .ZN(n3363) );
  AOI22_X1 U3207 ( .A1(n629), .A2(n5324), .B1(n568), .B2(n5472), .ZN(n5471) );
  AOI221_X1 U3208 ( .B1(n1957), .B2(n1975), .C1(n3703), .C2(n2124), .A(n963), 
        .ZN(n1956) );
  INV_X1 U3209 ( .A(n1959), .ZN(n3703) );
  INV_X1 U3210 ( .A(HADDR[8]), .ZN(n1772) );
  OAI222_X1 U3211 ( .A1(n2700), .A2(n3968), .B1(n3873), .B2(n442), .C1(n439), 
        .C2(n1809), .ZN(n4249) );
  NOR4_X1 U3212 ( .A1(Affpw6[0]), .A2(n635), .A3(n4380), .A4(n4381), .ZN(n3433) );
  OAI21_X1 U3213 ( .B1(n4382), .B2(n4383), .A(n4384), .ZN(n4380) );
  OAI222_X1 U3214 ( .A1(n439), .A2(n1814), .B1(n2700), .B2(n5112), .C1(n3885), 
        .C2(n448), .ZN(n4381) );
  NOR2_X1 U3215 ( .A1(n6447), .A2(n6445), .ZN(n4559) );
  OAI221_X1 U3216 ( .B1(n4180), .B2(n4153), .C1(n439), .C2(n1783), .A(n5177), 
        .ZN(n3417) );
  AOI211_X1 U3217 ( .C1(S2epw6), .C2(n5178), .A(Affpw6[7]), .B(n5179), .ZN(
        n5177) );
  NOR3_X1 U3218 ( .A1(n3792), .A2(n2549), .A3(S2epw6), .ZN(n5179) );
  AND2_X1 U3219 ( .A1(n1412), .A2(n3503), .ZN(n716) );
  XNOR2_X1 U3220 ( .A(n6509), .B(n6485), .ZN(n6498) );
  NAND2_X1 U3221 ( .A1(n254), .A2(n6503), .ZN(n6509) );
  NOR2_X1 U3222 ( .A1(n1000), .A2(n741), .ZN(n876) );
  AOI211_X1 U3223 ( .C1(n1763), .C2(n3512), .A(n3513), .B(n2593), .ZN(n3491)
         );
  OAI221_X1 U3224 ( .B1(n57), .B2(n3714), .C1(n266), .C2(n3858), .A(n3531), 
        .ZN(n3512) );
  OAI22_X1 U3225 ( .A1(n2124), .A2(n3516), .B1(n878), .B2(n2752), .ZN(n3513)
         );
  OAI21_X1 U3226 ( .B1(n266), .B2(n1482), .A(n505), .ZN(n3531) );
  AOI21_X1 U3227 ( .B1(n2154), .B2(n407), .A(HMASTER), .ZN(n203) );
  NAND2_X1 U3228 ( .A1(n1371), .A2(n4152), .ZN(n3872) );
  NOR2_X1 U3229 ( .A1(n4142), .A2(\Aphpw6[2] ), .ZN(\add_3107/B[1] ) );
  NAND3_X1 U3230 ( .A1(n4253), .A2(n3811), .A3(Qbfpw6_1), .ZN(n4252) );
  NAND3_X1 U3231 ( .A1(n1366), .A2(n2394), .A3(n5196), .ZN(n1361) );
  AND3_X1 U3232 ( .A1(n2393), .A2(n4144), .A3(n3911), .ZN(n5196) );
  NOR3_X1 U3233 ( .A1(n152), .A2(n946), .A3(n4149), .ZN(n151) );
  OAI222_X1 U3234 ( .A1(n538), .A2(n4756), .B1(n2733), .B2(n963), .C1(n267), 
        .C2(N701), .ZN(Qrohu6) );
  NOR3_X1 U3236 ( .A1(n2734), .A2(n2735), .A3(n2736), .ZN(n2733) );
  OAI211_X1 U3237 ( .C1(n2744), .C2(n4507), .A(n2746), .B(n2747), .ZN(n2734)
         );
  OAI22_X1 U3238 ( .A1(n5309), .A2(n6133), .B1(n6134), .B2(n2787), .ZN(n6110)
         );
  AOI22_X1 U3239 ( .A1(n5303), .A2(n6135), .B1(n3659), .B2(n6137), .ZN(n6134)
         );
  AOI221_X1 U3240 ( .B1(n5311), .B2(n4437), .C1(n5310), .C2(n6139), .A(n6140), 
        .ZN(n6133) );
  OAI221_X1 U3241 ( .B1(n8312), .B2(n2965), .C1(n8174), .C2(n1020), .A(n1021), 
        .ZN(n1018) );
  OAI221_X1 U3242 ( .B1(n2390), .B2(n631), .C1(n2392), .C2(n3347), .A(n6406), 
        .ZN(n3360) );
  AOI22_X1 U3243 ( .A1(n5280), .A2(n5324), .B1(n568), .B2(n5290), .ZN(n6406)
         );
  NAND4_X1 U3244 ( .A1(n5931), .A2(n5932), .A3(n5933), .A4(n5934), .ZN(n1228)
         );
  AOI222_X1 U3245 ( .A1(n2882), .A2(n8228), .B1(n2988), .B2(n8234), .C1(n2886), 
        .C2(n8236), .ZN(n5933) );
  AOI221_X1 U3246 ( .B1(n2985), .B2(n8232), .C1(n2884), .C2(n8230), .A(n5936), 
        .ZN(n5934) );
  AOI222_X1 U3247 ( .A1(n2852), .A2(n8237), .B1(n2978), .B2(n8233), .C1(n2866), 
        .C2(n8239), .ZN(n5932) );
  NAND4_X1 U3248 ( .A1(n5502), .A2(n5503), .A3(n5504), .A4(n5505), .ZN(n900)
         );
  AOI221_X1 U3249 ( .B1(n2985), .B2(n8198), .C1(n2884), .C2(n8199), .A(n5524), 
        .ZN(n5504) );
  AOI211_X1 U3250 ( .C1(n2858), .C2(n8200), .A(n5508), .B(n5509), .ZN(n5505)
         );
  AOI221_X1 U3251 ( .B1(n2866), .B2(n8203), .C1(n2852), .C2(n8201), .A(n5525), 
        .ZN(n5503) );
  NAND4_X1 U3252 ( .A1(n4845), .A2(n4846), .A3(n4847), .A4(n4848), .ZN(n904)
         );
  NOR4_X1 U3254 ( .A1(HWDATA[27]), .A2(HWDATA[25]), .A3(HWDATA[18]), .A4(
        HWDATA[16]), .ZN(n4847) );
  NOR4_X1 U3255 ( .A1(HWDATA[31]), .A2(HWDATA[30]), .A3(HWDATA[29]), .A4(
        HWDATA[28]), .ZN(n4848) );
  NOR4_X1 U3257 ( .A1(n2691), .A2(n2689), .A3(n2686), .A4(n2679), .ZN(n4845)
         );
  OAI221_X1 U3258 ( .B1(n2459), .B2(n631), .C1(n2447), .C2(n459), .A(n5488), 
        .ZN(n4731) );
  AOI22_X1 U3259 ( .A1(n5280), .A2(n5489), .B1(n568), .B2(n5281), .ZN(n5488)
         );
  INV_X1 U3260 ( .A(SLEEPING), .ZN(n5237) );
  NAND2_X1 U3261 ( .A1(n1144), .A2(n354), .ZN(n1966) );
  OAI22_X1 U3262 ( .A1(n4446), .A2(n2304), .B1(n2550), .B2(n3817), .ZN(n5132)
         );
  INV_X1 U3263 ( .A(n3817), .ZN(n2304) );
  OAI22_X1 U3264 ( .A1(n4446), .A2(n2310), .B1(n2550), .B2(n3792), .ZN(n5178)
         );
  INV_X1 U3265 ( .A(n3792), .ZN(n2310) );
  AOI21_X1 U3266 ( .B1(n3571), .B2(n1924), .A(n1916), .ZN(n1914) );
  NOR3_X1 U3267 ( .A1(n4386), .A2(n3822), .A3(n4254), .ZN(n4382) );
  AOI211_X1 U3268 ( .C1(n3960), .C2(n762), .A(n2819), .B(n8335), .ZN(Pvuhu6)
         );
  INV_X1 U3269 ( .A(n2824), .ZN(n3960) );
  OAI211_X1 U3270 ( .C1(n2821), .C2(n8293), .A(n906), .B(n2823), .ZN(n2819) );
  AOI211_X1 U3271 ( .C1(n3985), .C2(n762), .A(n2221), .B(n8337), .ZN(Ztuhu6)
         );
  OAI211_X1 U3272 ( .C1(n2223), .C2(n8287), .A(n906), .B(n2225), .ZN(n2221) );
  AOI211_X1 U3273 ( .C1(n3961), .C2(n762), .A(n4469), .B(n8343), .ZN(Bpthu6)
         );
  OAI211_X1 U3274 ( .C1(n3613), .C2(n8249), .A(n897), .B(n3619), .ZN(n4469) );
  AOI211_X1 U3275 ( .C1(n3978), .C2(n762), .A(n3155), .B(n8338), .ZN(Ltuhu6)
         );
  OAI211_X1 U3276 ( .C1(n3157), .C2(n8226), .A(n906), .B(n3159), .ZN(n3155) );
  AOI211_X1 U3277 ( .C1(n3975), .C2(n762), .A(n4037), .B(n8347), .ZN(Enthu6)
         );
  OAI211_X1 U3278 ( .C1(n3627), .C2(n5198), .A(n897), .B(n3633), .ZN(n4037) );
  AOI211_X1 U3279 ( .C1(n3972), .C2(n762), .A(n4842), .B(n8351), .ZN(Asthu6)
         );
  INV_X1 U3280 ( .A(n4843), .ZN(n3972) );
  OAI211_X1 U3281 ( .C1(n3927), .C2(n5193), .A(n897), .B(n3933), .ZN(n4842) );
  AOI211_X1 U3282 ( .C1(n3946), .C2(n762), .A(n3485), .B(n8340), .ZN(Jsuhu6)
         );
  OAI211_X1 U3283 ( .C1(n3487), .C2(n5134), .A(n897), .B(n3489), .ZN(n3485) );
  AOI211_X1 U3284 ( .C1(n3973), .C2(n762), .A(n3088), .B(n8355), .ZN(Mivhu6)
         );
  OAI211_X1 U3285 ( .C1(n3090), .C2(n4839), .A(n897), .B(n3092), .ZN(n3088) );
  AOI211_X1 U3286 ( .C1(n3951), .C2(n762), .A(n2966), .B(n8349), .ZN(Osthu6)
         );
  OAI211_X1 U3287 ( .C1(n2968), .C2(n4281), .A(n906), .B(n2970), .ZN(n2966) );
  AOI211_X1 U3288 ( .C1(n3988), .C2(n762), .A(n4274), .B(n8354), .ZN(Cmthu6)
         );
  INV_X1 U3289 ( .A(n4276), .ZN(n3988) );
  OAI211_X1 U3290 ( .C1(n3665), .C2(n3268), .A(n897), .B(n3671), .ZN(n4274) );
  AOI211_X1 U3291 ( .C1(n3990), .C2(n762), .A(n2467), .B(n8341), .ZN(Vruhu6)
         );
  INV_X1 U3292 ( .A(n2472), .ZN(n3990) );
  OAI211_X1 U3293 ( .C1(n2469), .C2(n8286), .A(n906), .B(n2471), .ZN(n2467) );
  AOI211_X1 U3294 ( .C1(n3955), .C2(n762), .A(n2461), .B(n8348), .ZN(Vsthu6)
         );
  OAI211_X1 U3296 ( .C1(n2463), .C2(n8238), .A(n906), .B(n2465), .ZN(n2461) );
  AOI211_X1 U3297 ( .C1(n3954), .C2(n762), .A(n2600), .B(n8352), .ZN(Trthu6)
         );
  OAI211_X1 U3298 ( .C1(n2602), .C2(n5209), .A(n906), .B(n2604), .ZN(n2600) );
  AOI211_X1 U3299 ( .C1(n3977), .C2(n762), .A(n2257), .B(n8342), .ZN(Zgthu6)
         );
  OAI211_X1 U3300 ( .C1(n2259), .C2(n5129), .A(n906), .B(n2261), .ZN(n2257) );
  AOI211_X1 U3301 ( .C1(n3957), .C2(n762), .A(n2352), .B(n8339), .ZN(Xsuhu6)
         );
  INV_X1 U3302 ( .A(n2357), .ZN(n3957) );
  OAI211_X1 U3303 ( .C1(n2354), .C2(n5128), .A(n906), .B(n2356), .ZN(n2352) );
  AOI211_X1 U3304 ( .C1(n762), .C2(n3193), .A(n3194), .B(n8346), .ZN(Lnthu6)
         );
  OAI21_X1 U3305 ( .B1(n3196), .B2(n8290), .A(n3198), .ZN(n3194) );
  NAND2_X1 U3306 ( .A1(n897), .A2(n3199), .ZN(n3193) );
  AOI211_X1 U3307 ( .C1(n762), .C2(n3856), .A(n3857), .B(n8350), .ZN(Hsthu6)
         );
  OAI21_X1 U3308 ( .B1(n3859), .B2(n8289), .A(n3861), .ZN(n3857) );
  NAND2_X1 U3309 ( .A1(n897), .A2(n3862), .ZN(n3856) );
  AOI211_X1 U3310 ( .C1(n762), .C2(n3552), .A(n3553), .B(n8332), .ZN(J6vhu6)
         );
  OAI21_X1 U3311 ( .B1(n3555), .B2(n8288), .A(n3557), .ZN(n3553) );
  NAND2_X1 U3312 ( .A1(n897), .A2(n3558), .ZN(n3552) );
  AOI211_X1 U3313 ( .C1(n762), .C2(n2520), .A(n2521), .B(n8336), .ZN(Uuuhu6)
         );
  OAI21_X1 U3314 ( .B1(n2523), .B2(n8202), .A(n2525), .ZN(n2521) );
  NAND2_X1 U3315 ( .A1(n897), .A2(n2526), .ZN(n2520) );
  AOI211_X1 U3316 ( .C1(n762), .C2(n3536), .A(n3537), .B(n8353), .ZN(Jmthu6)
         );
  OAI21_X1 U3317 ( .B1(n3539), .B2(n5216), .A(n3541), .ZN(n3537) );
  NAND2_X1 U3318 ( .A1(n897), .A2(n3542), .ZN(n3536) );
  INV_X1 U3319 ( .A(n2480), .ZN(n1889) );
  OAI21_X1 U3320 ( .B1(n6423), .B2(n5564), .A(n5572), .ZN(n4397) );
  AOI21_X1 U3321 ( .B1(n3836), .B2(n3835), .A(n6454), .ZN(n6423) );
  NOR4_X1 U3322 ( .A1(n5775), .A2(n4133), .A3(n8175), .A4(n4694), .ZN(n6454)
         );
  AOI21_X1 U3323 ( .B1(n5065), .B2(n6529), .A(n6533), .ZN(n5921) );
  NOR3_X1 U3324 ( .A1(n1149), .A2(n999), .A3(n3397), .ZN(n1139) );
  OAI21_X1 U3325 ( .B1(n3885), .B2(n3763), .A(n5904), .ZN(n2386) );
  NAND3_X1 U3326 ( .A1(n80), .A2(n5312), .A3(n52), .ZN(n5904) );
  OAI221_X1 U3327 ( .B1(n2111), .B2(n3620), .C1(n7381), .C2(n1376), .A(n1408), 
        .ZN(n7936) );
  AOI222_X1 U3328 ( .A1(n2119), .A2(n8298), .B1(n1410), .B2(n1411), .C1(n1412), 
        .C2(n801), .ZN(n1408) );
  OAI22_X1 U3329 ( .A1(n2549), .A2(n2535), .B1(n2550), .B2(n5156), .ZN(n5155)
         );
  NOR2_X1 U3330 ( .A1(n4826), .A2(n522), .ZN(n1730) );
  INV_X1 U3331 ( .A(n2893), .ZN(n4188) );
  INV_X1 U3332 ( .A(n6503), .ZN(n3351) );
  OAI22_X1 U3333 ( .A1(n2549), .A2(G3epw6), .B1(n2550), .B2(n2533), .ZN(n4796)
         );
  INV_X1 U3334 ( .A(G3epw6), .ZN(n2533) );
  OAI221_X1 U3335 ( .B1(n1640), .B2(n961), .C1(n7355), .C2(N701), .A(n1641), 
        .ZN(n7944) );
  AND3_X1 U3336 ( .A1(n1644), .A2(n1645), .A3(n1646), .ZN(n1640) );
  NAND3_X1 U3337 ( .A1(n1642), .A2(n228), .A3(n1643), .ZN(n1641) );
  AND4_X1 U3338 ( .A1(n3757), .A2(n3122), .A3(n447), .A4(n1452), .ZN(n1645) );
  OAI221_X1 U3339 ( .B1(n1707), .B2(n961), .C1(n228), .C2(N701), .A(n1708), 
        .ZN(n7946) );
  AND2_X1 U3340 ( .A1(n1710), .A2(n1711), .ZN(n1707) );
  OAI211_X1 U3341 ( .C1(n536), .C2(n4826), .A(n808), .B(n1643), .ZN(n1708) );
  AOI221_X1 U3342 ( .B1(n1628), .B2(n1724), .C1(n1725), .C2(n230), .A(n2128), 
        .ZN(n1710) );
  INV_X1 U3343 ( .A(n1576), .ZN(n2694) );
  AOI22_X1 U3344 ( .A1(n3793), .A2(n2745), .B1(n2332), .B2(n4254), .ZN(n4510)
         );
  INV_X1 U3345 ( .A(n3793), .ZN(n2332) );
  OAI22_X1 U3346 ( .A1(n2549), .A2(n3797), .B1(n2537), .B2(n4331), .ZN(n4327)
         );
  NOR2_X1 U3347 ( .A1(n2280), .A2(n4253), .ZN(n4331) );
  AOI22_X1 U3348 ( .A1(Qbfpw6_1), .A2(n4254), .B1(n4255), .B2(n4256), .ZN(
        n4251) );
  INV_X1 U3349 ( .A(n6154), .ZN(n2226) );
  OAI22_X1 U3350 ( .A1(n450), .A2(n5270), .B1(n8299), .B2(n1997), .ZN(n8034)
         );
  OAI22_X1 U3351 ( .A1(n450), .A2(n4701), .B1(n8312), .B2(n1997), .ZN(n8022)
         );
  OAI22_X1 U3352 ( .A1(n451), .A2(n4700), .B1(n8313), .B2(n1997), .ZN(n8021)
         );
  OAI22_X1 U3353 ( .A1(n451), .A2(n3673), .B1(n8314), .B2(n1997), .ZN(n8035)
         );
  AOI22_X1 U3354 ( .A1(n2226), .A2(n4459), .B1(n6154), .B2(n8200), .ZN(n6159)
         );
  AOI21_X1 U3355 ( .B1(n2550), .B2(Qbfpw6[30]), .A(n3798), .ZN(n5424) );
  AOI21_X1 U3356 ( .B1(n2549), .B2(n5094), .A(n3794), .ZN(n5091) );
  AND2_X1 U3357 ( .A1(Ntkbx6[7]), .A2(n3477), .ZN(K5ihu6) );
  OAI22_X1 U3358 ( .A1(n697), .A2(n1780), .B1(n696), .B2(n4811), .ZN(n3477) );
  AND2_X1 U3359 ( .A1(Ntkbx6[4]), .A2(n3148), .ZN(M1ihu6) );
  OAI22_X1 U3360 ( .A1(n701), .A2(n1793), .B1(n696), .B2(n4783), .ZN(n3148) );
  NAND2_X1 U3361 ( .A1(n1755), .A2(n1576), .ZN(n3522) );
  OAI211_X1 U3362 ( .C1(n3459), .C2(n4538), .A(n4539), .B(n4540), .ZN(n4537)
         );
  OAI221_X1 U3363 ( .B1(n4541), .B2(n4542), .C1(n228), .C2(n4538), .A(n517), 
        .ZN(n4540) );
  NAND3_X1 U3364 ( .A1(n4538), .A2(n516), .A3(n4551), .ZN(n4539) );
  NAND2_X1 U3365 ( .A1(n4557), .A2(n4558), .ZN(n4538) );
  AOI21_X1 U3366 ( .B1(Qbfpw6_0), .B2(n4253), .A(n4385), .ZN(n4383) );
  AOI21_X1 U3367 ( .B1(n2549), .B2(n4386), .A(n3822), .ZN(n4385) );
  INV_X1 U3368 ( .A(n4143), .ZN(n2363) );
  AOI21_X1 U3369 ( .B1(n1219), .B2(n883), .A(n877), .ZN(n1218) );
  AND2_X1 U3370 ( .A1(Ntkbx6[3]), .A2(n4113), .ZN(E0ihu6) );
  OAI22_X1 U3371 ( .A1(n697), .A2(n1798), .B1(n4787), .B2(n2297), .ZN(n4113)
         );
  INV_X1 U3372 ( .A(n3022), .ZN(n1913) );
  AOI21_X1 U3373 ( .B1(n2732), .B2(n3802), .A(n2539), .ZN(n5108) );
  INV_X1 U3374 ( .A(Qbfpw6[28]), .ZN(n2539) );
  NOR2_X1 U3375 ( .A1(n2602), .A2(n2942), .ZN(n7263) );
  INV_X1 U3376 ( .A(n3657), .ZN(n2942) );
  OAI211_X1 U3377 ( .C1(n8352), .C2(n5209), .A(n3658), .B(n2604), .ZN(n3657)
         );
  OAI21_X1 U3378 ( .B1(n3769), .B2(n672), .A(n5210), .ZN(n3658) );
  NOR2_X1 U3379 ( .A1(n3927), .A2(n2770), .ZN(H4phu6) );
  INV_X1 U3380 ( .A(n3929), .ZN(n2770) );
  OAI211_X1 U3381 ( .C1(n8351), .C2(n5193), .A(n3932), .B(n3933), .ZN(n3929)
         );
  OAI21_X1 U3382 ( .B1(n2776), .B2(n672), .A(n5197), .ZN(n3932) );
  NOR2_X1 U3383 ( .A1(n3555), .A2(n2648), .ZN(Qyohu6) );
  INV_X1 U3384 ( .A(n3747), .ZN(n2648) );
  OAI211_X1 U3385 ( .C1(n8332), .C2(n8288), .A(n3748), .B(n3557), .ZN(n3747)
         );
  OAI21_X1 U3386 ( .B1(n2649), .B2(n672), .A(n3037), .ZN(n3748) );
  AND2_X1 U3387 ( .A1(Nvkbx6[4]), .A2(n5103), .ZN(Alkhu6) );
  OAI22_X1 U3388 ( .A1(n733), .A2(n4783), .B1(n736), .B2(n1793), .ZN(n5103) );
  AND2_X1 U3389 ( .A1(Nvkbx6[3]), .A2(n2677), .ZN(Sjkhu6) );
  OAI22_X1 U3390 ( .A1(n2264), .A2(n4787), .B1(n736), .B2(n1798), .ZN(n2677)
         );
  AND2_X1 U3391 ( .A1(Nvkbx6[5]), .A2(n3782), .ZN(Imkhu6) );
  OAI22_X1 U3392 ( .A1(n2264), .A2(n4782), .B1(n736), .B2(n1788), .ZN(n3782)
         );
  AND3_X1 U3393 ( .A1(n840), .A2(n2096), .A3(n842), .ZN(n819) );
  NAND3_X1 U3394 ( .A1(n843), .A2(n844), .A3(n883), .ZN(n842) );
  INV_X1 U3395 ( .A(n6162), .ZN(n2227) );
  INV_X1 U3396 ( .A(n4636), .ZN(n2708) );
  OAI22_X1 U3397 ( .A1(n2382), .A2(n3114), .B1(n3116), .B2(n2584), .ZN(Xdvhu6)
         );
  INV_X1 U3398 ( .A(n2386), .ZN(n3116) );
  INV_X1 U3399 ( .A(n2382), .ZN(n2584) );
  NOR2_X1 U3400 ( .A1(n961), .A2(n2590), .ZN(n2382) );
  OAI22_X1 U3401 ( .A1(n4111), .A2(n1364), .B1(n1369), .B2(n4116), .ZN(n7923)
         );
  AOI21_X1 U3402 ( .B1(n1351), .B2(n1371), .A(n4112), .ZN(n1369) );
  OAI22_X1 U3403 ( .A1(n536), .A2(N701), .B1(n1546), .B2(n961), .ZN(n7942) );
  NOR4_X1 U3404 ( .A1(n1547), .A2(n1548), .A3(n1549), .A4(n1550), .ZN(n1546)
         );
  OAI221_X1 U3405 ( .B1(n4685), .B2(n1482), .C1(n4205), .C2(n3709), .A(n4215), 
        .ZN(n1550) );
  NAND4_X1 U3406 ( .A1(n1630), .A2(n2268), .A3(n3805), .A4(n4616), .ZN(n1547)
         );
  NOR2_X1 U3407 ( .A1(n3090), .A2(n1829), .ZN(n7268) );
  INV_X1 U3408 ( .A(n3636), .ZN(n1829) );
  OAI211_X1 U3409 ( .C1(n8355), .C2(n4839), .A(n3637), .B(n3092), .ZN(n3636)
         );
  OAI21_X1 U3410 ( .B1(n1831), .B2(n672), .A(n4001), .ZN(n3637) );
  NOR2_X1 U3411 ( .A1(n3196), .A2(n2660), .ZN(Uwdpw6) );
  INV_X1 U3412 ( .A(n3584), .ZN(n2660) );
  OAI211_X1 U3413 ( .C1(n8346), .C2(n8290), .A(n3585), .B(n3198), .ZN(n3584)
         );
  OAI21_X1 U3414 ( .B1(n339), .B2(n672), .A(n3930), .ZN(n3585) );
  NOR2_X1 U3415 ( .A1(n3627), .A2(n2652), .ZN(n7266) );
  INV_X1 U3416 ( .A(n3629), .ZN(n2652) );
  OAI211_X1 U3417 ( .C1(n8347), .C2(n5198), .A(n3632), .B(n3633), .ZN(n3629)
         );
  OAI21_X1 U3418 ( .B1(n335), .B2(n672), .A(n4010), .ZN(n3632) );
  NOR2_X1 U3419 ( .A1(n3157), .A2(n2688), .ZN(n7260) );
  INV_X1 U3420 ( .A(n3674), .ZN(n2688) );
  OAI211_X1 U3421 ( .C1(n8338), .C2(n8226), .A(n3675), .B(n3159), .ZN(n3674)
         );
  OAI21_X1 U3422 ( .B1(n2689), .B2(n672), .A(n8227), .ZN(n3675) );
  NOR2_X1 U3423 ( .A1(n2469), .A2(n2678), .ZN(n7265) );
  INV_X1 U3424 ( .A(n3651), .ZN(n2678) );
  OAI211_X1 U3425 ( .C1(n8341), .C2(n8286), .A(n3652), .B(n2471), .ZN(n3651)
         );
  OAI21_X1 U3426 ( .B1(n2679), .B2(n672), .A(n3310), .ZN(n3652) );
  NOR2_X1 U3427 ( .A1(n2463), .A2(n2943), .ZN(n7272) );
  INV_X1 U3428 ( .A(n3621), .ZN(n2943) );
  OAI211_X1 U3429 ( .C1(n8348), .C2(n8238), .A(n3622), .B(n2465), .ZN(n3621)
         );
  OAI21_X1 U3430 ( .B1(n4134), .B2(n672), .A(n8239), .ZN(n3622) );
  NOR2_X1 U3431 ( .A1(n2523), .A2(n2670), .ZN(Zzohu6) );
  INV_X1 U3432 ( .A(n3599), .ZN(n2670) );
  OAI211_X1 U3433 ( .C1(n8336), .C2(n8202), .A(n3600), .B(n2525), .ZN(n3599)
         );
  OAI21_X1 U3434 ( .B1(n2671), .B2(n672), .A(n8203), .ZN(n3600) );
  INV_X1 U3435 ( .A(n1996), .ZN(n4695) );
  INV_X1 U3436 ( .A(n4632), .ZN(n2443) );
  NOR2_X1 U3437 ( .A1(n2968), .A2(n2944), .ZN(n7273) );
  INV_X1 U3438 ( .A(n3594), .ZN(n2944) );
  OAI211_X1 U3439 ( .C1(n8349), .C2(n4281), .A(n3595), .B(n2970), .ZN(n3594)
         );
  OAI21_X1 U3440 ( .B1(n4126), .B2(n672), .A(n4293), .ZN(n3595) );
  OR4_X1 U3441 ( .A1(Affpw6[6]), .A2(n635), .A3(n4508), .A4(n4509), .ZN(n3428)
         );
  NOR3_X1 U3442 ( .A1(E2epw6), .A2(n2549), .A3(n3793), .ZN(n4508) );
  OAI222_X1 U3443 ( .A1(n4275), .A2(n442), .B1(n4510), .B2(n4511), .C1(n4154), 
        .C2(n1786), .ZN(n4509) );
  INV_X1 U3444 ( .A(n4836), .ZN(n2341) );
  INV_X1 U3445 ( .A(n4262), .ZN(n2351) );
  OAI21_X1 U3446 ( .B1(n5303), .B2(n2787), .A(n5305), .ZN(n5301) );
  OAI211_X1 U3447 ( .C1(n5306), .C2(n2788), .A(n5308), .B(n2787), .ZN(n5305)
         );
  OR3_X1 U3448 ( .A1(n5309), .A2(n5310), .A3(n5311), .ZN(n5308) );
  INV_X1 U3449 ( .A(n4411), .ZN(n2383) );
  INV_X1 U3450 ( .A(n5156), .ZN(n2535) );
  NAND2_X1 U3451 ( .A1(n6147), .A2(n4790), .ZN(n6109) );
  NAND3_X1 U3452 ( .A1(n3290), .A2(n6149), .A3(n5309), .ZN(n6147) );
  OAI22_X1 U3453 ( .A1(n3869), .A2(n3292), .B1(n3300), .B2(n5306), .ZN(n6149)
         );
  AND2_X1 U3454 ( .A1(n1891), .A2(n2977), .ZN(n398) );
  NAND2_X1 U3455 ( .A1(n5302), .A2(n6530), .ZN(n5919) );
  AND2_X1 U3456 ( .A1(n5174), .A2(n5173), .ZN(n5087) );
  INV_X1 U3457 ( .A(n797), .ZN(n3503) );
  NAND2_X1 U3458 ( .A1(n5312), .A2(n6534), .ZN(n5920) );
  NOR2_X1 U3459 ( .A1(Qbfpw6_3), .A2(n4256), .ZN(n4825) );
  INV_X1 U3460 ( .A(n3801), .ZN(n2293) );
  INV_X1 U3461 ( .A(n3797), .ZN(n2280) );
  BUF_X1 U3462 ( .A(n963), .Z(n961) );
  INV_X1 U3463 ( .A(n1426), .ZN(n3488) );
  INV_X1 U3464 ( .A(n4414), .ZN(n2429) );
  AND3_X1 U3465 ( .A1(n911), .A2(n2098), .A3(n1323), .ZN(n1293) );
  NOR3_X1 U3466 ( .A1(n1135), .A2(n1324), .A3(n1136), .ZN(n1323) );
  INV_X1 U3467 ( .A(n4840), .ZN(n2435) );
  INV_X1 U3468 ( .A(n3820), .ZN(n2316) );
  INV_X1 U3469 ( .A(n3791), .ZN(n2294) );
  INV_X1 U3470 ( .A(n3818), .ZN(n2312) );
  INV_X1 U3471 ( .A(n3819), .ZN(n2287) );
  BUF_X1 U3472 ( .A(n403), .Z(n731) );
  INV_X1 U3473 ( .A(n3806), .ZN(n2313) );
  NAND2_X1 U3474 ( .A1(n5388), .A2(n5389), .ZN(n3334) );
  NAND3_X1 U3475 ( .A1(n5390), .A2(n523), .A3(n3108), .ZN(n5389) );
  OAI21_X1 U3476 ( .B1(n228), .B2(n5391), .A(n2418), .ZN(n5388) );
  INV_X1 U3477 ( .A(n3821), .ZN(n2291) );
  INV_X1 U3478 ( .A(n5194), .ZN(n2464) );
  NAND2_X1 U3479 ( .A1(n1107), .A2(n1108), .ZN(n1050) );
  INV_X1 U3480 ( .A(n3807), .ZN(n2279) );
  AND2_X1 U3481 ( .A1(n4614), .A2(n4615), .ZN(n3442) );
  NAND3_X1 U3483 ( .A1(n2550), .A2(n2709), .A3(Qbfpw6_2), .ZN(n4615) );
  OAI22_X1 U3484 ( .A1(n2732), .A2(n4617), .B1(n2330), .B2(n4618), .ZN(n4614)
         );
  NOR2_X1 U3485 ( .A1(Qbfpw6_2), .A2(n4256), .ZN(n4618) );
  INV_X1 U3486 ( .A(n1413), .ZN(n3505) );
  AND2_X1 U3487 ( .A1(n2569), .A2(n454), .ZN(n213) );
  OAI221_X1 U3488 ( .B1(n455), .B2(n4546), .C1(n457), .C2(n5256), .A(n2548), 
        .ZN(n454) );
  AND4_X1 U3489 ( .A1(n1135), .A2(n1136), .A3(n1137), .A4(n2098), .ZN(n1107)
         );
  NAND2_X1 U3490 ( .A1(n911), .A2(n4046), .ZN(n1137) );
  NAND2_X1 U3491 ( .A1(n1777), .A2(n1778), .ZN(n7952) );
  OAI221_X1 U3492 ( .B1(n2644), .B2(n2818), .C1(n1781), .C2(n3851), .A(n3617), 
        .ZN(n1778) );
  INV_X1 U3493 ( .A(n5173), .ZN(n2582) );
  INV_X1 U3494 ( .A(n3808), .ZN(n2309) );
  INV_X1 U3495 ( .A(n3813), .ZN(n2282) );
  INV_X1 U3496 ( .A(n3812), .ZN(n2317) );
  INV_X1 U3497 ( .A(n3809), .ZN(n2286) );
  INV_X1 U3498 ( .A(n3810), .ZN(n2290) );
  INV_X1 U3499 ( .A(n3816), .ZN(n2283) );
  INV_X1 U3500 ( .A(n3815), .ZN(n2296) );
  INV_X1 U3501 ( .A(n3814), .ZN(n2320) );
  INV_X1 U3502 ( .A(n2430), .ZN(n4157) );
  AND3_X1 U3503 ( .A1(n4401), .A2(n4394), .A3(n4748), .ZN(n399) );
  INV_X1 U3504 ( .A(n6481), .ZN(n3112) );
  INV_X1 U3505 ( .A(n5903), .ZN(n2590) );
  INV_X1 U3506 ( .A(n5090), .ZN(n2298) );
  OAI22_X1 U3507 ( .A1(n5091), .A2(n5092), .B1(n3794), .B2(n5093), .ZN(n5090)
         );
  NAND2_X1 U3508 ( .A1(Qbfpw6_5), .A2(n2550), .ZN(n5093) );
  NOR2_X1 U3509 ( .A1(n2732), .A2(n5094), .ZN(n5092) );
  INV_X1 U3510 ( .A(n5107), .ZN(n2301) );
  OAI22_X1 U3511 ( .A1(n5108), .A2(n5109), .B1(n3802), .B2(n5110), .ZN(n5107)
         );
  NOR2_X1 U3512 ( .A1(n2549), .A2(n3802), .ZN(n5109) );
  NAND2_X1 U3513 ( .A1(n2550), .A2(Qbfpw6[28]), .ZN(n5110) );
  AND2_X1 U3514 ( .A1(Ntkbx6[1]), .A2(n2958), .ZN(Oxhhu6) );
  OAI22_X1 U3515 ( .A1(n4548), .A2(n2297), .B1(n701), .B2(n2959), .ZN(n2958)
         );
  AND2_X1 U3516 ( .A1(Nvkbx6[1]), .A2(n4283), .ZN(Chkhu6) );
  OAI22_X1 U3517 ( .A1(n733), .A2(n4548), .B1(n736), .B2(n2959), .ZN(n4283) );
  OR3_X1 U3518 ( .A1(n4824), .A2(n4254), .A3(n3796), .ZN(n4823) );
  INV_X1 U3519 ( .A(n1365), .ZN(n4111) );
  OR3_X1 U3520 ( .A1(n1343), .A2(n1002), .A3(n1278), .ZN(n1328) );
  AND2_X1 U3521 ( .A1(n5713), .A2(n5714), .ZN(n3438) );
  OAI22_X1 U3522 ( .A1(n5715), .A2(n2732), .B1(n5717), .B2(n3795), .ZN(n5713)
         );
  OR3_X1 U3523 ( .A1(n5715), .A2(n3795), .A3(n4254), .ZN(n5714) );
  NOR2_X1 U3524 ( .A1(Qbfpw6_4), .A2(n4256), .ZN(n5717) );
  AND2_X1 U3525 ( .A1(Qbfpw6[30]), .A2(n3798), .ZN(n5423) );
  AND2_X1 U3526 ( .A1(Ntkbx6[2]), .A2(n2401), .ZN(Wyhhu6) );
  OAI22_X1 U3527 ( .A1(n701), .A2(n1802), .B1(n2297), .B2(n4795), .ZN(n2401)
         );
  AND2_X1 U3528 ( .A1(Ntkbx6[5]), .A2(n2552), .ZN(U2ihu6) );
  OAI22_X1 U3529 ( .A1(n701), .A2(n1788), .B1(n2297), .B2(n4782), .ZN(n2552)
         );
  AND2_X1 U3530 ( .A1(Nvkbx6[2]), .A2(n3455), .ZN(Kikhu6) );
  OAI22_X1 U3531 ( .A1(n2264), .A2(n4795), .B1(n734), .B2(n1802), .ZN(n3455)
         );
  AND2_X1 U3532 ( .A1(Nvkbx6[7]), .A2(n2308), .ZN(Yokhu6) );
  OAI22_X1 U3533 ( .A1(n2264), .A2(n4811), .B1(n736), .B2(n1780), .ZN(n2308)
         );
  NOR2_X1 U3534 ( .A1(n3487), .A2(n2666), .ZN(n7264) );
  INV_X1 U3535 ( .A(n3646), .ZN(n2666) );
  OAI211_X1 U3536 ( .C1(n8340), .C2(n5134), .A(n3647), .B(n3489), .ZN(n3646)
         );
  OAI21_X1 U3537 ( .B1(n2667), .B2(n672), .A(n4061), .ZN(n3647) );
  NOR2_X1 U3538 ( .A1(n2259), .A2(n2663), .ZN(n7267) );
  INV_X1 U3539 ( .A(n3641), .ZN(n2663) );
  OAI211_X1 U3540 ( .C1(n8342), .C2(n5129), .A(n3642), .B(n2261), .ZN(n3641)
         );
  OAI21_X1 U3541 ( .B1(n2664), .B2(n672), .A(n4005), .ZN(n3642) );
  NOR2_X1 U3542 ( .A1(n2821), .A2(n2675), .ZN(n7270) );
  INV_X1 U3543 ( .A(n3605), .ZN(n2675) );
  OAI211_X1 U3544 ( .C1(n8335), .C2(n8293), .A(n3606), .B(n2823), .ZN(n3605)
         );
  OAI21_X1 U3545 ( .B1(n2676), .B2(n672), .A(n8294), .ZN(n3606) );
  NOR2_X1 U3546 ( .A1(n2354), .A2(n2684), .ZN(n7262) );
  INV_X1 U3547 ( .A(n3662), .ZN(n2684) );
  OAI211_X1 U3548 ( .C1(n8339), .C2(n5128), .A(n3663), .B(n2356), .ZN(n3662)
         );
  OAI21_X1 U3549 ( .B1(n2686), .B2(n672), .A(n3870), .ZN(n3663) );
  NOR2_X1 U3550 ( .A1(n2223), .A2(n2690), .ZN(n7269) );
  INV_X1 U3551 ( .A(n3609), .ZN(n2690) );
  OAI211_X1 U3552 ( .C1(n8337), .C2(n8287), .A(n3610), .B(n2225), .ZN(n3609)
         );
  OAI21_X1 U3553 ( .B1(n2691), .B2(n672), .A(n3669), .ZN(n3610) );
  NOR2_X1 U3554 ( .A1(n3539), .A2(n2949), .ZN(V4phu6) );
  INV_X1 U3555 ( .A(n3589), .ZN(n2949) );
  OAI211_X1 U3556 ( .C1(n8353), .C2(n5216), .A(n3590), .B(n3541), .ZN(n3589)
         );
  OAI21_X1 U3557 ( .B1(n905), .B2(n672), .A(n3030), .ZN(n3590) );
  NOR2_X1 U3558 ( .A1(n3665), .A2(n2938), .ZN(n7254) );
  INV_X1 U3559 ( .A(n3667), .ZN(n2938) );
  OAI211_X1 U3560 ( .C1(n8354), .C2(n3268), .A(n3670), .B(n3671), .ZN(n3667)
         );
  OAI21_X1 U3561 ( .B1(n700), .B2(n672), .A(n3276), .ZN(n3670) );
  INV_X1 U3562 ( .A(n1213), .ZN(n2828) );
  INV_X1 U3563 ( .A(n2172), .ZN(n2651) );
  INV_X1 U3564 ( .A(n2074), .ZN(n3520) );
  AOI22_X1 U3565 ( .A1(n8298), .A2(n4695), .B1(n1411), .B2(n451), .ZN(n2074)
         );
  OAI21_X1 U3566 ( .B1(n619), .B2(n4029), .A(n3223), .ZN(n2705) );
  OAI21_X1 U3567 ( .B1(n1856), .B2(n1325), .A(n1857), .ZN(n4729) );
  OAI21_X1 U3568 ( .B1(n4182), .B2(n5980), .A(n5981), .ZN(n4714) );
  NAND3_X1 U3569 ( .A1(n844), .A2(n1277), .A3(n1183), .ZN(n5981) );
  NAND2_X1 U3570 ( .A1(n1325), .A2(n5406), .ZN(n2202) );
  OAI21_X1 U3571 ( .B1(n1856), .B2(n1325), .A(n5545), .ZN(n4730) );
  INV_X1 U3572 ( .A(n1893), .ZN(n2976) );
  NOR3_X1 U3573 ( .A1(n2057), .A2(n579), .A3(n2056), .ZN(n2665) );
  NAND3_X1 U3574 ( .A1(n4694), .A2(n8175), .A3(n6040), .ZN(n6038) );
  NOR2_X1 U3575 ( .A1(n2015), .A2(n4033), .ZN(n542) );
  NOR4_X1 U3576 ( .A1(n2057), .A2(n579), .A3(n4032), .A4(n4035), .ZN(n642) );
  NAND2_X1 U3577 ( .A1(n3634), .A2(HWDATA[15]), .ZN(n1835) );
  NOR2_X1 U3578 ( .A1(n4329), .A2(n4406), .ZN(n1345) );
  NOR2_X1 U3579 ( .A1(n2262), .A2(n2699), .ZN(n518) );
  OAI21_X1 U3580 ( .B1(n1763), .B2(n5219), .A(n2731), .ZN(n4153) );
  NAND3_X1 U3581 ( .A1(n1182), .A2(n4054), .A3(n4306), .ZN(n988) );
  INV_X1 U3582 ( .A(n4705), .ZN(n2712) );
  OAI21_X1 U3583 ( .B1(n1763), .B2(n5219), .A(n2731), .ZN(n448) );
  OAI21_X1 U3584 ( .B1(n1763), .B2(n5219), .A(n2731), .ZN(n442) );
  NAND4_X1 U3585 ( .A1(n5406), .A2(n4410), .A3(n4160), .A4(n4182), .ZN(n4788)
         );
  INV_X1 U3586 ( .A(n4691), .ZN(n2713) );
  NOR3_X1 U3587 ( .A1(n1565), .A2(n52), .A3(n4084), .ZN(n4213) );
  NOR3_X1 U3588 ( .A1(n4214), .A2(n2933), .A3(n4588), .ZN(n4212) );
  OAI21_X1 U3589 ( .B1(n5042), .B2(n1493), .A(n4216), .ZN(n4214) );
  INV_X1 U3590 ( .A(n5345), .ZN(n2825) );
  INV_X1 U3591 ( .A(HWDATA[7]), .ZN(n4134) );
  INV_X1 U3592 ( .A(HWDATA[6]), .ZN(n4126) );
  NOR2_X1 U3593 ( .A1(n4637), .A2(n3099), .ZN(n57) );
  NOR2_X1 U3594 ( .A1(n101), .A2(n99), .ZN(n97) );
  NAND2_X1 U3595 ( .A1(n1969), .A2(n844), .ZN(n1006) );
  NAND4_X1 U3596 ( .A1(n1504), .A2(n493), .A3(n524), .A4(n2731), .ZN(n4261) );
  NAND2_X1 U3597 ( .A1(n2132), .A2(n844), .ZN(n989) );
  NOR3_X1 U3598 ( .A1(n3083), .A2(n5070), .A3(n4261), .ZN(n4342) );
  NOR3_X1 U3599 ( .A1(n2698), .A2(n1939), .A3(n2262), .ZN(n70) );
  NAND2_X1 U3600 ( .A1(n3634), .A2(HWDATA[2]), .ZN(n905) );
  NAND2_X1 U3601 ( .A1(n1969), .A2(n1182), .ZN(n985) );
  NOR3_X1 U3602 ( .A1(n3712), .A2(n3763), .A3(n3083), .ZN(n3049) );
  AOI221_X1 U3603 ( .B1(n3121), .B2(n2866), .C1(n8137), .C2(n2852), .A(n4714), 
        .ZN(n1180) );
  NAND2_X1 U3604 ( .A1(n5406), .A2(n5972), .ZN(n2197) );
  NOR2_X1 U3605 ( .A1(n5042), .A2(n470), .ZN(n2933) );
  AOI221_X1 U3606 ( .B1(n8296), .B2(n2866), .C1(n8295), .C2(n2852), .A(n2856), 
        .ZN(n1158) );
  AOI221_X1 U3607 ( .B1(n3037), .B2(n2866), .C1(n8147), .C2(n2852), .A(n2856), 
        .ZN(n1085) );
  NOR2_X1 U3608 ( .A1(n4054), .A2(n4405), .ZN(n1277) );
  NOR2_X1 U3609 ( .A1(n3882), .A2(n3470), .ZN(n1274) );
  NAND2_X1 U3610 ( .A1(n3634), .A2(HWDATA[1]), .ZN(n700) );
  NOR3_X1 U3611 ( .A1(n4187), .A2(n875), .A3(n2256), .ZN(n3188) );
  NAND4_X1 U3612 ( .A1(n3077), .A2(n1462), .A3(n228), .A4(n7381), .ZN(n1458)
         );
  NAND2_X1 U3613 ( .A1(n5545), .A2(n5971), .ZN(n2195) );
  NAND4_X1 U3614 ( .A1(n90), .A2(n88), .A3(n1594), .A4(n4635), .ZN(n1518) );
  AOI222_X1 U3615 ( .A1(n2488), .A2(n4932), .B1(n2489), .B2(n4855), .C1(n1698), 
        .C2(n464), .ZN(n2487) );
  OAI221_X1 U3616 ( .B1(n2873), .B2(n2607), .C1(n3831), .C2(n4633), .A(n2874), 
        .ZN(n2872) );
  AOI222_X1 U3617 ( .A1(n1627), .A2(n2562), .B1(n2875), .B2(n4932), .C1(n2876), 
        .C2(n2124), .ZN(n2874) );
  INV_X1 U3618 ( .A(HWDATA[16]), .ZN(n2664) );
  OAI221_X1 U3619 ( .B1(n2367), .B2(n387), .C1(n2360), .C2(n459), .A(n5341), 
        .ZN(n3371) );
  AOI22_X1 U3620 ( .A1(n629), .A2(n5342), .B1(n5280), .B2(n5343), .ZN(n5341)
         );
  INV_X1 U3621 ( .A(HWDATA[18]), .ZN(n2667) );
  NAND2_X1 U3622 ( .A1(n5483), .A2(n5406), .ZN(n2199) );
  NAND3_X1 U3623 ( .A1(n2961), .A2(n3634), .A3(HALTED), .ZN(n397) );
  INV_X1 U3624 ( .A(HWDATA[4]), .ZN(n2776) );
  INV_X1 U3625 ( .A(HWDATA[0]), .ZN(n1831) );
  AOI222_X1 U3626 ( .A1(n429), .A2(n428), .B1(n1673), .B2(n449), .C1(n1674), 
        .C2(n1675), .ZN(n1664) );
  OAI21_X1 U3627 ( .B1(n1686), .B2(n1687), .A(n1688), .ZN(n1673) );
  OAI22_X1 U3628 ( .A1(n1676), .A2(n3547), .B1(n1678), .B2(n2243), .ZN(n1675)
         );
  NAND4_X1 U3629 ( .A1(n519), .A2(n1684), .A3(n1595), .A4(n475), .ZN(n1688) );
  NOR2_X1 U3630 ( .A1(n4187), .A2(n270), .ZN(n1762) );
  NAND2_X1 U3631 ( .A1(n1325), .A2(n2969), .ZN(n1009) );
  INV_X1 U3632 ( .A(HWDATA[28]), .ZN(n2650) );
  OAI221_X1 U3633 ( .B1(n265), .B2(n504), .C1(n3804), .C2(n4749), .A(n4585), 
        .ZN(n810) );
  NOR3_X1 U3634 ( .A1(n4586), .A2(n3165), .A3(n1660), .ZN(n4585) );
  NOR4_X1 U3635 ( .A1(n482), .A2(n230), .A3(n4628), .A4(n4205), .ZN(n4586) );
  INV_X1 U3636 ( .A(HWDATA[25]), .ZN(n2644) );
  NOR3_X1 U3637 ( .A1(n1945), .A2(n4507), .A3(n4187), .ZN(n1512) );
  AOI221_X1 U3638 ( .B1(n4313), .B2(n476), .C1(n4314), .C2(n470), .A(n4315), 
        .ZN(n4312) );
  NOR3_X1 U3639 ( .A1(n230), .A2(n3749), .A3(n516), .ZN(n4315) );
  OAI21_X1 U3640 ( .B1(n1926), .B2(n2696), .A(n4319), .ZN(n4313) );
  OAI21_X1 U3641 ( .B1(n4566), .B2(n1925), .A(n4316), .ZN(n4314) );
  INV_X1 U3642 ( .A(HWDATA[10]), .ZN(n2653) );
  INV_X1 U3643 ( .A(HWDATA[11]), .ZN(n2655) );
  INV_X1 U3644 ( .A(HWDATA[12]), .ZN(n2654) );
  INV_X1 U3645 ( .A(HWDATA[13]), .ZN(n2657) );
  NOR3_X1 U3646 ( .A1(n4028), .A2(n620), .A3(n3144), .ZN(n586) );
  INV_X1 U3647 ( .A(HWDATA[3]), .ZN(n3769) );
  INV_X1 U3648 ( .A(HWDATA[5]), .ZN(n4072) );
  NOR4_X1 U3649 ( .A1(n4993), .A2(n4732), .A3(n3682), .A4(n4978), .ZN(n2588)
         );
  NOR3_X1 U3650 ( .A1(n4119), .A2(n1324), .A3(n4118), .ZN(n2394) );
  AOI221_X1 U3651 ( .B1(n2563), .B2(n1763), .C1(n2564), .C2(n4263), .A(n2565), 
        .ZN(n2557) );
  OAI221_X1 U3652 ( .B1(n2566), .B2(n254), .C1(n270), .C2(n2266), .A(n2567), 
        .ZN(n2565) );
  OAI221_X1 U3653 ( .B1(n2568), .B2(n1572), .C1(n529), .C2(n3730), .A(n2570), 
        .ZN(n2564) );
  NOR2_X1 U3654 ( .A1(n1761), .A2(n1462), .ZN(n2566) );
  AOI221_X1 U3655 ( .B1(n70), .B2(n1465), .C1(n1466), .C2(n4635), .A(n1468), 
        .ZN(n1440) );
  OAI211_X1 U3656 ( .C1(n1493), .C2(n5037), .A(n1494), .B(n1495), .ZN(n1465)
         );
  OAI211_X1 U3657 ( .C1(n2277), .C2(n1939), .A(n1486), .B(n1487), .ZN(n1466)
         );
  OAI221_X1 U3658 ( .B1(n4608), .B2(n1470), .C1(n1471), .C2(n2547), .A(n1473), 
        .ZN(n1468) );
  NAND2_X1 U3659 ( .A1(n5406), .A2(n5971), .ZN(n2198) );
  INV_X1 U3660 ( .A(HWDATA[29]), .ZN(n2649) );
  NAND3_X1 U3661 ( .A1(n6547), .A2(n6548), .A3(n6549), .ZN(n6531) );
  AOI222_X1 U3662 ( .A1(n1540), .A2(n1620), .B1(n496), .B2(n3189), .C1(n4298), 
        .C2(n1642), .ZN(n6547) );
  NOR4_X1 U3663 ( .A1(n6550), .A2(n6551), .A3(n3165), .A4(n6552), .ZN(n6549)
         );
  AOI221_X1 U3664 ( .B1(n1520), .B2(n6556), .C1(n417), .C2(n6557), .A(n6558), 
        .ZN(n6548) );
  AOI221_X1 U3665 ( .B1(n1462), .B2(n1496), .C1(n1497), .C2(n4263), .A(n1498), 
        .ZN(n1439) );
  NAND3_X1 U3666 ( .A1(n1534), .A2(n4693), .A3(n1535), .ZN(n1496) );
  OAI221_X1 U3667 ( .B1(n3732), .B2(n4608), .C1(n3860), .C2(n4229), .A(n1531), 
        .ZN(n1497) );
  OAI222_X1 U3668 ( .A1(n1499), .A2(n2572), .B1(n270), .B2(n1501), .C1(n1502), 
        .C2(n2524), .ZN(n1498) );
  NAND3_X1 U3669 ( .A1(n5570), .A2(n5577), .A3(n5578), .ZN(n4439) );
  NAND3_X1 U3670 ( .A1(n2722), .A2(n8175), .A3(n5574), .ZN(n5578) );
  NAND4_X1 U3671 ( .A1(n2135), .A2(n1269), .A3(n1270), .A4(n994), .ZN(n1059)
         );
  OR2_X1 U3672 ( .A1(n1248), .A2(n4054), .ZN(n1269) );
  NAND3_X1 U3673 ( .A1(n1277), .A2(n3913), .A3(n1274), .ZN(n1270) );
  INV_X1 U3674 ( .A(n1278), .ZN(n2135) );
  NAND2_X1 U3675 ( .A1(n5972), .A2(n5545), .ZN(n2200) );
  AOI221_X1 U3676 ( .B1(n4908), .B2(n3025), .C1(n1624), .C2(n3074), .A(n3075), 
        .ZN(n3073) );
  INV_X1 U3677 ( .A(n4253), .ZN(n2732) );
  OAI221_X1 U3678 ( .B1(n2991), .B2(n3699), .C1(n2993), .C2(n2994), .A(n2995), 
        .ZN(n2505) );
  AOI22_X1 U3679 ( .A1(n2996), .A2(n2997), .B1(n3698), .B2(n2999), .ZN(n2995)
         );
  INV_X1 U3680 ( .A(n3000), .ZN(n3698) );
  OAI222_X1 U3681 ( .A1(n538), .A2(n3760), .B1(n4670), .B2(n1518), .C1(n3804), 
        .C2(n4749), .ZN(n1541) );
  NAND2_X1 U3682 ( .A1(n674), .A2(HWDATA[28]), .ZN(n3448) );
  NOR2_X1 U3683 ( .A1(n5042), .A2(n7514), .ZN(n1587) );
  OAI222_X1 U3684 ( .A1(n6553), .A2(n4265), .B1(n6554), .B2(n3766), .C1(n6555), 
        .C2(n4190), .ZN(n6550) );
  AOI21_X1 U3685 ( .B1(n4298), .B2(n266), .A(n4581), .ZN(n6555) );
  AOI21_X1 U3686 ( .B1(n1566), .B2(n7282), .A(n3829), .ZN(n6554) );
  AOI22_X1 U3687 ( .A1(n1723), .A2(n5013), .B1(n1951), .B2(n7374), .ZN(n6553)
         );
  OAI222_X1 U3688 ( .A1(n554), .A2(n555), .B1(n556), .B2(n557), .C1(n558), 
        .C2(n559), .ZN(n553) );
  OAI21_X1 U3689 ( .B1(n4932), .B2(n3761), .A(n3966), .ZN(n3025) );
  AOI211_X1 U3690 ( .C1(n1488), .C2(n1666), .A(n1667), .B(n1668), .ZN(n1665)
         );
  NOR3_X1 U3691 ( .A1(n3838), .A2(n266), .A3(n2594), .ZN(n1668) );
  OAI22_X1 U3692 ( .A1(n476), .A2(n2262), .B1(n5037), .B2(n3625), .ZN(n1666)
         );
  AOI211_X1 U3693 ( .C1(n1584), .C2(n3517), .A(n3518), .B(n3519), .ZN(n3516)
         );
  OAI21_X1 U3694 ( .B1(n3529), .B2(n4187), .A(n2267), .ZN(n3517) );
  OAI221_X1 U3695 ( .B1(n3521), .B2(n3522), .C1(n3523), .C2(n2277), .A(n3524), 
        .ZN(n3518) );
  NAND4_X1 U3696 ( .A1(n3911), .A2(n4046), .A3(n4118), .A4(n5195), .ZN(n4137)
         );
  NOR2_X1 U3698 ( .A1(n911), .A2(n4115), .ZN(n5195) );
  NAND2_X1 U3699 ( .A1(n5257), .A2(n6492), .ZN(n5387) );
  OAI211_X1 U3700 ( .C1(n1539), .C2(n505), .A(n4250), .B(n4650), .ZN(n6492) );
  AOI211_X1 U3702 ( .C1(n485), .C2(n55), .A(n56), .B(n517), .ZN(n53) );
  NAND3_X1 U3703 ( .A1(n228), .A2(n266), .A3(n57), .ZN(n55) );
  OAI21_X1 U3704 ( .B1(n5735), .B2(n2601), .A(n2731), .ZN(n5426) );
  INV_X1 U3705 ( .A(n5737), .ZN(n2601) );
  AOI21_X1 U3706 ( .B1(n878), .B2(n1761), .A(n5738), .ZN(n5737) );
  NAND2_X1 U3707 ( .A1(n5406), .A2(n1856), .ZN(n1894) );
  NAND2_X1 U3708 ( .A1(n3582), .A2(HWDATA[16]), .ZN(n2261) );
  NAND2_X1 U3709 ( .A1(n3582), .A2(HWDATA[18]), .ZN(n3489) );
  NAND2_X1 U3710 ( .A1(n674), .A2(HWDATA[12]), .ZN(n3753) );
  NOR2_X1 U3711 ( .A1(n548), .A2(n3201), .ZN(n2046) );
  NAND2_X1 U3712 ( .A1(n674), .A2(HWDATA[29]), .ZN(n3557) );
  NAND2_X1 U3713 ( .A1(n674), .A2(HWDATA[25]), .ZN(n2830) );
  NAND2_X1 U3714 ( .A1(n3582), .A2(HWDATA[23]), .ZN(n2823) );
  NAND2_X1 U3715 ( .A1(n674), .A2(HWDATA[20]), .ZN(n3159) );
  NAND2_X1 U3716 ( .A1(n3582), .A2(HWDATA[21]), .ZN(n2225) );
  NAND2_X1 U3717 ( .A1(n3582), .A2(HWDATA[17]), .ZN(n2471) );
  NAND2_X1 U3718 ( .A1(n674), .A2(HWDATA[8]), .ZN(n3633) );
  NAND2_X1 U3719 ( .A1(n674), .A2(HWDATA[19]), .ZN(n2356) );
  NAND2_X1 U3720 ( .A1(n3582), .A2(HWDATA[22]), .ZN(n2525) );
  NAND2_X1 U3721 ( .A1(n3582), .A2(HWDATA[9]), .ZN(n3198) );
  NOR2_X1 U3722 ( .A1(n1948), .A2(n4670), .ZN(n1607) );
  NOR4_X1 U3723 ( .A1(n1658), .A2(n1659), .A3(n1660), .A4(n1661), .ZN(n1644)
         );
  AOI211_X1 U3724 ( .C1(n4738), .C2(n1662), .A(n7374), .B(n7375), .ZN(n1659)
         );
  AOI21_X1 U3725 ( .B1(n1664), .B2(n1665), .A(n4512), .ZN(n1658) );
  NAND2_X1 U3726 ( .A1(n1663), .A2(n875), .ZN(n1662) );
  NAND2_X1 U3727 ( .A1(n5668), .A2(n5545), .ZN(n2193) );
  NOR2_X1 U3728 ( .A1(n3894), .A2(Jshpw6[4]), .ZN(n939) );
  OAI21_X1 U3729 ( .B1(n3243), .B2(n4670), .A(n3238), .ZN(n2849) );
  NOR2_X1 U3730 ( .A1(n527), .A2(n2157), .ZN(n2155) );
  NAND2_X1 U3731 ( .A1(n674), .A2(HWDATA[10]), .ZN(n2669) );
  NAND2_X1 U3732 ( .A1(n674), .A2(HWDATA[11]), .ZN(n2241) );
  NAND2_X1 U3733 ( .A1(n674), .A2(HWDATA[13]), .ZN(n3035) );
  NOR2_X1 U3734 ( .A1(n4572), .A2(n4993), .ZN(n1683) );
  NAND4_X1 U3736 ( .A1(n1907), .A2(n1576), .A3(n1908), .A4(n2262), .ZN(n1687)
         );
  NAND2_X1 U3737 ( .A1(n4670), .A2(n5042), .ZN(n1739) );
  XNOR2_X1 U3738 ( .A(n3000), .B(n2999), .ZN(n2997) );
  NAND2_X1 U3739 ( .A1(n5483), .A2(n5545), .ZN(n2196) );
  OAI211_X1 U3740 ( .C1(n7514), .C2(n4670), .A(n5037), .B(n4669), .ZN(n2773)
         );
  OAI221_X1 U3741 ( .B1(n2437), .B2(n3347), .C1(n2438), .C2(n3358), .A(n5327), 
        .ZN(n3312) );
  AOI22_X1 U3742 ( .A1(n568), .A2(n5328), .B1(n4763), .B2(n5329), .ZN(n5327)
         );
  NAND2_X1 U3743 ( .A1(n5668), .A2(n5406), .ZN(n2194) );
  INV_X1 U3744 ( .A(n1419), .ZN(n2131) );
  XNOR2_X1 U3745 ( .A(n2996), .B(n2997), .ZN(n2993) );
  OAI221_X1 U3746 ( .B1(n3623), .B2(n2907), .C1(n4233), .C2(n4512), .A(n4234), 
        .ZN(n4224) );
  NOR3_X1 U3747 ( .A1(n4238), .A2(n489), .A3(n4239), .ZN(n4233) );
  AOI222_X1 U3748 ( .A1(n4235), .A2(n429), .B1(n1620), .B2(n4236), .C1(n3630), 
        .C2(n2894), .ZN(n4234) );
  AND3_X1 U3749 ( .A1(n3188), .A2(n7381), .A3(n1456), .ZN(n4239) );
  OAI221_X1 U3750 ( .B1(n1740), .B2(n56), .C1(n1741), .C2(n508), .A(n1742), 
        .ZN(n1735) );
  OAI21_X1 U3751 ( .B1(n1743), .B2(n1612), .A(n1744), .ZN(n1742) );
  AOI21_X1 U3752 ( .B1(n1747), .B2(n1748), .A(n1749), .ZN(n1740) );
  AOI211_X1 U3753 ( .C1(n82), .C2(n266), .A(n1745), .B(n1746), .ZN(n1741) );
  NAND2_X1 U3754 ( .A1(n3582), .A2(HWDATA[7]), .ZN(n2465) );
  NAND2_X1 U3755 ( .A1(n674), .A2(HWDATA[3]), .ZN(n2604) );
  NAND2_X1 U3756 ( .A1(n3582), .A2(HWDATA[4]), .ZN(n3933) );
  NAND2_X1 U3757 ( .A1(n3582), .A2(HWDATA[6]), .ZN(n2970) );
  NAND2_X1 U3758 ( .A1(n3582), .A2(HWDATA[0]), .ZN(n3092) );
  NAND2_X1 U3759 ( .A1(n3582), .A2(HWDATA[5]), .ZN(n3861) );
  OAI221_X1 U3760 ( .B1(n2360), .B2(n3358), .C1(n2365), .C2(n459), .A(n5535), 
        .ZN(n3372) );
  AOI22_X1 U3761 ( .A1(n629), .A2(n5536), .B1(n568), .B2(n5537), .ZN(n5535) );
  OAI221_X1 U3762 ( .B1(n2442), .B2(n3347), .C1(n2437), .C2(n3358), .A(n5500), 
        .ZN(n3313) );
  AOI22_X1 U3763 ( .A1(n629), .A2(n5328), .B1(n568), .B2(n5501), .ZN(n5500) );
  NOR3_X1 U3764 ( .A1(n4555), .A2(n4670), .A3(n5002), .ZN(n2583) );
  NAND2_X1 U3765 ( .A1(n3725), .A2(n5390), .ZN(n4726) );
  NAND2_X1 U3766 ( .A1(n610), .A2(n2054), .ZN(n555) );
  INV_X1 U3767 ( .A(n4526), .ZN(n2719) );
  OAI211_X1 U3768 ( .C1(n2277), .C2(n4187), .A(n3267), .B(n2242), .ZN(n3263)
         );
  NAND3_X1 U3769 ( .A1(n1584), .A2(n4670), .A3(n3269), .ZN(n3267) );
  INV_X1 U3770 ( .A(n2916), .ZN(n2242) );
  INV_X1 U3771 ( .A(n1592), .ZN(n4672) );
  NOR2_X1 U3772 ( .A1(n1926), .A2(n3549), .ZN(n1456) );
  NAND4_X1 U3773 ( .A1(n2893), .A2(n1612), .A3(n3181), .A4(n90), .ZN(n3176) );
  OAI21_X1 U3774 ( .B1(n4054), .B2(n1282), .A(n1023), .ZN(n1278) );
  OAI21_X1 U3775 ( .B1(n1589), .B2(n464), .A(n470), .ZN(n79) );
  OAI21_X1 U3776 ( .B1(n2498), .B2(n4187), .A(n2250), .ZN(n2842) );
  INV_X1 U3777 ( .A(n544), .ZN(n3180) );
  NAND3_X1 U3778 ( .A1(n1539), .A2(n56), .A3(n37), .ZN(n1630) );
  NAND3_X1 U3779 ( .A1(n4572), .A2(n5042), .A3(n2585), .ZN(n1495) );
  OAI21_X1 U3780 ( .B1(n5025), .B2(n3966), .A(n2738), .ZN(n3075) );
  NOR2_X1 U3781 ( .A1(n3269), .A2(n475), .ZN(n5025) );
  NAND2_X1 U3782 ( .A1(n2876), .A2(n4187), .ZN(n3186) );
  NAND3_X1 U3783 ( .A1(n469), .A2(n2696), .A3(n471), .ZN(n258) );
  NAND3_X1 U3784 ( .A1(n472), .A2(n464), .A3(n473), .ZN(n471) );
  NAND4_X1 U3785 ( .A1(n2124), .A2(n474), .A3(n4910), .A4(n4932), .ZN(n469) );
  OAI21_X1 U3786 ( .B1(n3247), .B2(n4932), .A(n3000), .ZN(n3246) );
  INV_X1 U3787 ( .A(n1020), .ZN(n3481) );
  OAI21_X1 U3789 ( .B1(n3245), .B2(n4987), .A(n2994), .ZN(n3244) );
  INV_X1 U3790 ( .A(n548), .ZN(n4015) );
  AOI211_X1 U3791 ( .C1(n1744), .C2(n1752), .A(n2769), .B(n1737), .ZN(n2768)
         );
  AND3_X1 U3792 ( .A1(n2771), .A2(n476), .A3(n1685), .ZN(n2769) );
  OAI211_X1 U3793 ( .C1(n5042), .C2(n1948), .A(n270), .B(n2772), .ZN(n2771) );
  AOI21_X1 U3794 ( .B1(n2773), .B2(n464), .A(n2774), .ZN(n2772) );
  NAND3_X1 U3795 ( .A1(n3211), .A2(n4187), .A3(n518), .ZN(n3209) );
  INV_X1 U3796 ( .A(n2846), .ZN(n2272) );
  OAI22_X1 U3797 ( .A1(n3638), .A2(n6130), .B1(n6131), .B2(n6132), .ZN(n6112)
         );
  NAND2_X1 U3798 ( .A1(n1346), .A2(n4405), .ZN(n1284) );
  NAND2_X1 U3799 ( .A1(n3243), .A2(n4670), .ZN(n3238) );
  OAI22_X1 U3800 ( .A1(n485), .A2(n412), .B1(n3507), .B2(n56), .ZN(n3506) );
  AOI22_X1 U3801 ( .A1(n3508), .A2(n513), .B1(n3509), .B2(n1761), .ZN(n3507)
         );
  NOR2_X1 U3802 ( .A1(n265), .A2(n3838), .ZN(n3508) );
  NAND2_X1 U3803 ( .A1(n824), .A2(n1371), .ZN(n2085) );
  NAND2_X1 U3804 ( .A1(n847), .A2(n1371), .ZN(n2081) );
  NAND2_X1 U3805 ( .A1(n854), .A2(n1371), .ZN(n2079) );
  NAND2_X1 U3806 ( .A1(n863), .A2(n1371), .ZN(n2077) );
  OAI22_X1 U3807 ( .A1(n3837), .A2(n3746), .B1(n4226), .B2(n56), .ZN(n4225) );
  AOI21_X1 U3808 ( .B1(n1952), .B2(n4227), .A(n4228), .ZN(n4226) );
  OAI21_X1 U3809 ( .B1(n266), .B2(n4610), .A(n1470), .ZN(n4227) );
  NOR2_X1 U3810 ( .A1(n4024), .A2(n3200), .ZN(n2053) );
  NAND2_X1 U3811 ( .A1(n2893), .A2(n1538), .ZN(n2738) );
  NAND2_X1 U3812 ( .A1(n663), .A2(n2168), .ZN(n530) );
  AOI22_X1 U3813 ( .A1(n3062), .A2(n6125), .B1(n5321), .B2(n6126), .ZN(n6123)
         );
  INV_X1 U3814 ( .A(n5390), .ZN(n2444) );
  NOR2_X1 U3815 ( .A1(n3186), .A2(n3074), .ZN(n2898) );
  NAND3_X1 U3816 ( .A1(n56), .A2(n463), .A3(n1567), .ZN(n3498) );
  OAI21_X1 U3817 ( .B1(n3504), .B2(n4187), .A(n2251), .ZN(n3500) );
  AOI21_X1 U3818 ( .B1(n473), .B2(n470), .A(n2767), .ZN(n3504) );
  NOR2_X1 U3819 ( .A1(n532), .A2(n1820), .ZN(n527) );
  INV_X1 U3820 ( .A(n531), .ZN(n1820) );
  OAI21_X1 U3821 ( .B1(n4572), .B2(n5042), .A(n7381), .ZN(n3262) );
  INV_X1 U3822 ( .A(n648), .ZN(n3223) );
  AOI22_X1 U3823 ( .A1(n3550), .A2(n693), .B1(n808), .B2(n4826), .ZN(n3218) );
  NOR2_X1 U3824 ( .A1(n2849), .A2(n4579), .ZN(n3236) );
  INV_X1 U3825 ( .A(n2848), .ZN(n4579) );
  NAND2_X1 U3826 ( .A1(n3481), .A2(n1144), .ZN(n1023) );
  OAI21_X1 U3827 ( .B1(n2676), .B2(n892), .A(n1842), .ZN(n7974) );
  OAI21_X1 U3828 ( .B1(n891), .B2(n2676), .A(n8292), .ZN(n1842) );
  OAI21_X1 U3829 ( .B1(n356), .B2(n892), .A(n1839), .ZN(n7973) );
  OAI21_X1 U3830 ( .B1(n891), .B2(n356), .A(n8150), .ZN(n1839) );
  INV_X1 U3831 ( .A(n2159), .ZN(n3136) );
  OAI221_X1 U3832 ( .B1(n56), .B2(n3746), .C1(n3804), .C2(n4608), .A(n3257), 
        .ZN(n3256) );
  AOI21_X1 U3833 ( .B1(n878), .B2(n1620), .A(n3217), .ZN(n3257) );
  AOI22_X1 U3834 ( .A1(n415), .A2(n1937), .B1(n1938), .B2(n693), .ZN(n1933) );
  OAI21_X1 U3835 ( .B1(n878), .B2(n1994), .A(n56), .ZN(n1937) );
  AOI22_X1 U3836 ( .A1(n1674), .A2(n3174), .B1(n3175), .B2(n4932), .ZN(n3168)
         );
  NAND3_X1 U3837 ( .A1(n3176), .A2(n3177), .A3(n3178), .ZN(n3174) );
  NAND3_X1 U3838 ( .A1(n2848), .A2(n1918), .A3(n3179), .ZN(n3177) );
  NAND3_X1 U3839 ( .A1(n473), .A2(n230), .A3(n519), .ZN(n3178) );
  OAI21_X1 U3840 ( .B1(n3561), .B2(n5772), .A(n2731), .ZN(n4154) );
  AOI22_X1 U3841 ( .A1(n5773), .A2(n5774), .B1(n692), .B2(n272), .ZN(n5772) );
  AOI21_X1 U3842 ( .B1(n5776), .B2(n7355), .A(n491), .ZN(n5773) );
  NOR2_X1 U3843 ( .A1(n5775), .A2(n2562), .ZN(n5774) );
  NAND2_X1 U3844 ( .A1(n3247), .A2(n4932), .ZN(n3000) );
  INV_X1 U3845 ( .A(n3288), .ZN(n2969) );
  NOR2_X1 U3846 ( .A1(n3952), .A2(n5797), .ZN(n2170) );
  AOI21_X1 U3847 ( .B1(n2113), .B2(n4673), .A(n2500), .ZN(n5797) );
  INV_X1 U3848 ( .A(n663), .ZN(n3156) );
  INV_X1 U3849 ( .A(n903), .ZN(n2856) );
  OAI211_X1 U3850 ( .C1(n1762), .C2(n3549), .A(n449), .B(n529), .ZN(n4319) );
  INV_X1 U3851 ( .A(n655), .ZN(n3208) );
  OAI21_X1 U3852 ( .B1(n4134), .B2(n892), .A(n1845), .ZN(n7975) );
  OAI21_X1 U3853 ( .B1(n891), .B2(n4134), .A(n8237), .ZN(n1845) );
  OAI21_X1 U3854 ( .B1(n4126), .B2(n892), .A(n1833), .ZN(n7971) );
  OAI21_X1 U3855 ( .B1(n891), .B2(n4126), .A(n8149), .ZN(n1833) );
  NAND2_X1 U3856 ( .A1(n1613), .A2(n1457), .ZN(n2378) );
  OAI21_X1 U3857 ( .B1(n2671), .B2(n894), .A(n1830), .ZN(n7970) );
  OAI21_X1 U3858 ( .B1(n891), .B2(n2671), .A(n8201), .ZN(n1830) );
  OAI211_X1 U3859 ( .C1(n523), .C2(n3625), .A(n1598), .B(n482), .ZN(n1578) );
  NAND3_X1 U3860 ( .A1(n1599), .A2(n5225), .A3(n7282), .ZN(n1598) );
  OAI21_X1 U3861 ( .B1(n349), .B2(n894), .A(n907), .ZN(n7881) );
  OAI21_X1 U3862 ( .B1(n891), .B2(n349), .A(n8135), .ZN(n907) );
  INV_X1 U3863 ( .A(n3687), .ZN(n2818) );
  OAI21_X1 U3864 ( .B1(n332), .B2(n894), .A(n1827), .ZN(n7969) );
  OAI21_X1 U3865 ( .B1(n891), .B2(n332), .A(n8257), .ZN(n1827) );
  NAND2_X1 U3866 ( .A1(n3245), .A2(n4987), .ZN(n2994) );
  OAI221_X1 U3867 ( .B1(n2524), .B2(n3727), .C1(n504), .C2(n3746), .A(n506), 
        .ZN(n487) );
  AOI21_X1 U3868 ( .B1(n507), .B2(n230), .A(n509), .ZN(n506) );
  NAND3_X1 U3869 ( .A1(n510), .A2(n511), .A3(n512), .ZN(n507) );
  NAND4_X1 U3871 ( .A1(n518), .A2(n519), .A3(n93), .A4(n449), .ZN(n510) );
  INV_X1 U3872 ( .A(n1595), .ZN(n5047) );
  AND2_X1 U3873 ( .A1(n5972), .A2(n2969), .ZN(n2201) );
  INV_X1 U3874 ( .A(n4267), .ZN(n2723) );
  NAND4_X1 U3875 ( .A1(n966), .A2(n4145), .A3(n967), .A4(n968), .ZN(n965) );
  NOR3_X1 U3876 ( .A1(n944), .A2(n152), .A3(n4402), .ZN(n968) );
  OAI21_X1 U3877 ( .B1(n922), .B2(n3886), .A(n8253), .ZN(n966) );
  AOI22_X1 U3878 ( .A1(n939), .A2(n3886), .B1(n918), .B2(Jshpw6[4]), .ZN(n967)
         );
  INV_X1 U3879 ( .A(n2446), .ZN(n3007) );
  INV_X1 U3880 ( .A(n1000), .ZN(n3479) );
  OAI21_X1 U3881 ( .B1(n352), .B2(n894), .A(n1797), .ZN(n7958) );
  OAI21_X1 U3882 ( .B1(n891), .B2(n352), .A(n8295), .ZN(n1797) );
  NOR2_X1 U3883 ( .A1(n4029), .A2(n3201), .ZN(n2704) );
  NAND3_X1 U3884 ( .A1(n5032), .A2(n3271), .A3(n5033), .ZN(n4304) );
  NAND3_X1 U3885 ( .A1(n1594), .A2(n4672), .A3(n4317), .ZN(n5032) );
  AOI21_X1 U3886 ( .B1(n518), .B2(n2921), .A(n3270), .ZN(n5033) );
  AOI21_X1 U3887 ( .B1(n4015), .B2(n562), .A(n551), .ZN(n560) );
  OAI211_X1 U3888 ( .C1(n3201), .C2(n3225), .A(n3204), .B(n566), .ZN(n562) );
  AND3_X1 U3889 ( .A1(n555), .A2(n3215), .A3(n558), .ZN(n566) );
  INV_X1 U3890 ( .A(n4834), .ZN(n2700) );
  OAI21_X1 U3891 ( .B1(n894), .B2(n1835), .A(n1836), .ZN(n7972) );
  OAI21_X1 U3892 ( .B1(n891), .B2(n1835), .A(n8240), .ZN(n1836) );
  OAI21_X1 U3893 ( .B1(n892), .B2(n905), .A(n1789), .ZN(n7955) );
  OAI21_X1 U3894 ( .B1(n891), .B2(n905), .A(n8142), .ZN(n1789) );
  INV_X1 U3895 ( .A(n1755), .ZN(n2267) );
  NAND2_X1 U3896 ( .A1(n1672), .A2(n2262), .ZN(n1670) );
  OAI21_X1 U3897 ( .B1(n2679), .B2(n894), .A(n1848), .ZN(n7976) );
  OAI21_X1 U3898 ( .B1(n891), .B2(n2679), .A(n8151), .ZN(n1848) );
  OAI21_X1 U3899 ( .B1(n2686), .B2(n894), .A(n1800), .ZN(n7959) );
  OAI21_X1 U3900 ( .B1(n703), .B2(n2686), .A(n8143), .ZN(n1800) );
  OAI21_X1 U3901 ( .B1(n2689), .B2(n894), .A(n1810), .ZN(n7963) );
  OAI21_X1 U3902 ( .B1(n703), .B2(n2689), .A(n8225), .ZN(n1810) );
  OAI21_X1 U3903 ( .B1(n2691), .B2(n894), .A(n1821), .ZN(n7967) );
  OAI21_X1 U3904 ( .B1(n703), .B2(n2691), .A(n8148), .ZN(n1821) );
  OAI21_X1 U3907 ( .B1(n700), .B2(n892), .A(n702), .ZN(n7851) );
  OAI21_X1 U3908 ( .B1(n891), .B2(n700), .A(n8134), .ZN(n702) );
  INV_X1 U3909 ( .A(n619), .ZN(n3225) );
  OAI21_X1 U3910 ( .B1(n2776), .B2(n894), .A(n1813), .ZN(n7964) );
  OAI21_X1 U3911 ( .B1(n703), .B2(n2776), .A(n8146), .ZN(n1813) );
  OAI21_X1 U3912 ( .B1(n2650), .B2(n894), .A(n1807), .ZN(n7962) );
  OAI21_X1 U3913 ( .B1(n703), .B2(n2650), .A(n8278), .ZN(n1807) );
  OAI21_X1 U3914 ( .B1(n3769), .B2(n894), .A(n1803), .ZN(n7960) );
  OAI21_X1 U3915 ( .B1(n703), .B2(n3769), .A(n8144), .ZN(n1803) );
  OAI21_X1 U3916 ( .B1(n2649), .B2(n894), .A(n1818), .ZN(n7966) );
  OAI21_X1 U3917 ( .B1(n703), .B2(n2649), .A(n8147), .ZN(n1818) );
  AOI21_X1 U3918 ( .B1(n2845), .B2(n2846), .A(n2847), .ZN(n2844) );
  XNOR2_X1 U3919 ( .A(n2848), .B(n2849), .ZN(n2845) );
  OAI21_X1 U3920 ( .B1(n2667), .B2(n892), .A(n1787), .ZN(n7954) );
  OAI21_X1 U3921 ( .B1(n891), .B2(n2667), .A(n8141), .ZN(n1787) );
  OAI21_X1 U3922 ( .B1(n2664), .B2(n894), .A(n1773), .ZN(n7950) );
  OAI21_X1 U3923 ( .B1(n891), .B2(n2664), .A(n8139), .ZN(n1773) );
  OAI21_X1 U3924 ( .B1(n2632), .B2(n892), .A(n1768), .ZN(n7948) );
  OAI21_X1 U3925 ( .B1(n891), .B2(n2632), .A(n8137), .ZN(n1768) );
  OAI21_X1 U3926 ( .B1(n1831), .B2(n894), .A(n1765), .ZN(n7947) );
  OAI21_X1 U3927 ( .B1(n891), .B2(n1831), .A(n8136), .ZN(n1765) );
  INV_X1 U3928 ( .A(n2151), .ZN(n2858) );
  NAND3_X1 U3929 ( .A1(n1732), .A2(n1733), .A3(n1734), .ZN(n1725) );
  AOI222_X1 U3930 ( .A1(n1761), .A2(n693), .B1(n1762), .B2(n1685), .C1(n1763), 
        .C2(n1620), .ZN(n1732) );
  AOI221_X1 U3931 ( .B1(n1750), .B2(n529), .C1(n1751), .C2(n1752), .A(n1753), 
        .ZN(n1733) );
  NOR4_X1 U3932 ( .A1(n1735), .A2(n1736), .A3(n1613), .A4(n1737), .ZN(n1734)
         );
  NAND2_X1 U3933 ( .A1(n4222), .A2(n480), .ZN(n259) );
  NAND4_X1 U3934 ( .A1(n4341), .A2(n4932), .A3(n7355), .A4(n481), .ZN(n480) );
  NOR2_X1 U3935 ( .A1(n508), .A2(n449), .ZN(n481) );
  NOR2_X1 U3936 ( .A1(n4512), .A2(n56), .ZN(n61) );
  INV_X1 U3937 ( .A(n1744), .ZN(n2696) );
  INV_X1 U3938 ( .A(n1698), .ZN(n2235) );
  INV_X1 U3939 ( .A(n2921), .ZN(n1967) );
  NAND3_X1 U3940 ( .A1(n4559), .A2(n4560), .A3(n4561), .ZN(n4558) );
  OAI21_X1 U3941 ( .B1(n4562), .B2(n4563), .A(n1642), .ZN(n4560) );
  OAI221_X1 U3942 ( .B1(n47), .B2(n254), .C1(n49), .C2(n463), .A(n51), .ZN(n38) );
  AOI21_X1 U3943 ( .B1(SLEEPHOLDACKn), .B2(n2502), .A(n2124), .ZN(n49) );
  AOI21_X1 U3944 ( .B1(n61), .B2(n62), .A(n63), .ZN(n47) );
  NOR2_X1 U3945 ( .A1(n52), .A2(n53), .ZN(n51) );
  INV_X1 U3946 ( .A(n938), .ZN(n4146) );
  NAND2_X1 U3947 ( .A1(n1595), .A2(n4669), .ZN(n1593) );
  INV_X1 U3948 ( .A(n4530), .ZN(n2507) );
  NAND2_X1 U3949 ( .A1(n4322), .A2(n3209), .ZN(n2374) );
  NAND4_X1 U3950 ( .A1(n90), .A2(n4323), .A3(n5047), .A4(n4635), .ZN(n4322) );
  NAND2_X1 U3951 ( .A1(n5042), .A2(n475), .ZN(n4323) );
  INV_X1 U3952 ( .A(n1083), .ZN(n3439) );
  NAND2_X1 U3953 ( .A1(n4033), .A2(n4036), .ZN(n641) );
  AND2_X1 U3954 ( .A1(n3582), .A2(HWDATA[14]), .ZN(n2532) );
  AND2_X1 U3955 ( .A1(n3582), .A2(HWDATA[27]), .ZN(n4023) );
  AND2_X1 U3956 ( .A1(n3582), .A2(HWDATA[30]), .ZN(n2681) );
  AND2_X1 U3957 ( .A1(n3582), .A2(HWDATA[31]), .ZN(n2796) );
  AND2_X1 U3958 ( .A1(n3582), .A2(HWDATA[26]), .ZN(n2422) );
  NAND2_X1 U3959 ( .A1(n5973), .A2(n4160), .ZN(n1638) );
  AND2_X1 U3960 ( .A1(n3582), .A2(HWDATA[24]), .ZN(n3758) );
  INV_X1 U3961 ( .A(n41), .ZN(n1947) );
  AND2_X1 U3962 ( .A1(n5978), .A2(n4182), .ZN(n5668) );
  NAND3_X1 U3963 ( .A1(n2740), .A2(n2073), .A3(n2741), .ZN(n2735) );
  NAND4_X1 U3964 ( .A1(n2742), .A2(n2743), .A3(n1952), .A4(n56), .ZN(n2741) );
  NAND4_X1 U3965 ( .A1(n2571), .A2(n1951), .A3(n3550), .A4(n4263), .ZN(n2740)
         );
  OR4_X1 U3966 ( .A1(n1660), .A2(n2898), .A3(n2875), .A4(n2899), .ZN(n2889) );
  OR4_X1 U3967 ( .A1(n1686), .A2(n4978), .A3(n7514), .A4(n270), .ZN(n2951) );
  AND3_X1 U3968 ( .A1(n4410), .A2(n4182), .A3(n1857), .ZN(n5973) );
  NAND3_X1 U3969 ( .A1(n67), .A2(n3186), .A3(n2598), .ZN(n4208) );
  INV_X1 U3970 ( .A(n3175), .ZN(n2598) );
  INV_X1 U3971 ( .A(n2876), .ZN(n3757) );
  NAND2_X1 U3972 ( .A1(n1857), .A2(n5978), .ZN(n5980) );
  INV_X1 U3973 ( .A(n1324), .ZN(n4046) );
  INV_X1 U3974 ( .A(n957), .ZN(n4149) );
  INV_X1 U3975 ( .A(n3240), .ZN(n3699) );
  AND3_X1 U3976 ( .A1(n1595), .A2(n4670), .A3(n1948), .ZN(n2774) );
  AND3_X1 U3977 ( .A1(n5483), .A2(n4459), .A3(n2969), .ZN(n5481) );
  INV_X1 U3978 ( .A(n4557), .ZN(n3082) );
  AND2_X1 U3979 ( .A1(n5545), .A2(n3634), .ZN(n5544) );
  INV_X1 U3980 ( .A(n1695), .ZN(n2238) );
  AOI221_X1 U3981 ( .B1(n4978), .B2(n1697), .C1(n5042), .C2(n1698), .A(n1699), 
        .ZN(n1695) );
  NAND2_X1 U3982 ( .A1(n559), .A2(n3216), .ZN(n574) );
  AND2_X1 U3983 ( .A1(n3894), .A2(n920), .ZN(n940) );
  OR2_X1 U3984 ( .A1(n699), .A2(n400), .ZN(n7850) );
  AND3_X1 U3985 ( .A1(n897), .A2(n4673), .A3(n698), .ZN(n400) );
  INV_X1 U3986 ( .A(n1183), .ZN(n4333) );
  NAND3_X1 U3987 ( .A1(n844), .A2(n4054), .A3(n4306), .ZN(n984) );
  INV_X1 U3988 ( .A(n420), .ZN(n824) );
  INV_X1 U3989 ( .A(n431), .ZN(n809) );
  NAND3_X1 U3990 ( .A1(n1182), .A2(n1345), .A3(n1311), .ZN(n125) );
  NOR3_X1 U3991 ( .A1(n3226), .A2(n4029), .A3(n3208), .ZN(n591) );
  NAND2_X1 U3992 ( .A1(n1086), .A2(n1182), .ZN(n990) );
  NOR2_X1 U3993 ( .A1(n636), .A2(n4015), .ZN(n609) );
  NAND2_X1 U3994 ( .A1(n2132), .A2(n1182), .ZN(n1004) );
  NAND3_X1 U3995 ( .A1(n1287), .A2(n4405), .A3(n1182), .ZN(n113) );
  NAND3_X1 U3996 ( .A1(n844), .A2(n1277), .A3(n1345), .ZN(n992) );
  NOR2_X1 U3997 ( .A1(n1247), .A2(n4301), .ZN(n1074) );
  NAND2_X1 U3998 ( .A1(n1086), .A2(n844), .ZN(n1005) );
  NOR2_X1 U3999 ( .A1(n4137), .A2(n1108), .ZN(n2434) );
  NOR2_X1 U4000 ( .A1(n1247), .A2(n4330), .ZN(n1066) );
  OAI221_X1 U4001 ( .B1(n4749), .B2(n3705), .C1(n265), .C2(n2603), .A(n4080), 
        .ZN(n1932) );
  INV_X1 U4002 ( .A(n2089), .ZN(n2883) );
  INV_X1 U4003 ( .A(n2097), .ZN(n2987) );
  INV_X1 U4004 ( .A(n2105), .ZN(n2897) );
  INV_X1 U4005 ( .A(n2095), .ZN(n2992) );
  INV_X1 U4006 ( .A(n2101), .ZN(n2989) );
  INV_X1 U4007 ( .A(n2093), .ZN(n2885) );
  INV_X1 U4008 ( .A(n2099), .ZN(n2983) );
  INV_X1 U4009 ( .A(n2091), .ZN(n2906) );
  AOI21_X1 U4010 ( .B1(n4187), .B2(n1538), .A(n5029), .ZN(n3028) );
  AND3_X1 U4011 ( .A1(n1442), .A2(n2262), .A3(n3527), .ZN(n5029) );
  NAND4_X1 U4012 ( .A1(n1183), .A2(n844), .A3(n4405), .A4(n4054), .ZN(n827) );
  AOI21_X1 U4013 ( .B1(n1684), .B2(n3211), .A(n1918), .ZN(n1701) );
  AOI211_X1 U4014 ( .C1(n3201), .C2(n657), .A(n591), .B(n658), .ZN(n652) );
  AOI211_X1 U4015 ( .C1(n3201), .C2(n3223), .A(n655), .B(n656), .ZN(n653) );
  AOI211_X1 U4016 ( .C1(n2806), .C2(n1706), .A(n2807), .B(n2808), .ZN(n2805)
         );
  NOR3_X1 U4017 ( .A1(n3571), .A2(n2806), .A3(n5065), .ZN(n2808) );
  NAND4_X1 U4018 ( .A1(n3692), .A2(n3693), .A3(n3694), .A4(n3695), .ZN(n1890)
         );
  NOR3_X1 U4019 ( .A1(n3708), .A2(Tzfpw6[20]), .A3(Tzfpw6[12]), .ZN(n3692) );
  NOR4_X1 U4020 ( .A1(n3704), .A2(Tzfpw6[1]), .A3(Tzfpw6[10]), .A4(Tzfpw6[16]), 
        .ZN(n3693) );
  NOR4_X1 U4021 ( .A1(n3700), .A2(Tzfpw6[8]), .A3(Tzfpw6[11]), .A4(Tzfpw6[19]), 
        .ZN(n3694) );
  NAND3_X1 U4022 ( .A1(n1023), .A2(n827), .A3(n1181), .ZN(n999) );
  OAI21_X1 U4023 ( .B1(n1182), .B2(n844), .A(n843), .ZN(n1181) );
  AOI21_X1 U4024 ( .B1(n1325), .B2(n1854), .A(n389), .ZN(n703) );
  NAND3_X1 U4025 ( .A1(n3439), .A2(n1277), .A3(n1346), .ZN(n991) );
  OAI221_X1 U4026 ( .B1(n2605), .B2(n1482), .C1(n3749), .C2(n4749), .A(n1901), 
        .ZN(n1899) );
  AOI22_X1 U4027 ( .A1(n1902), .A2(n3837), .B1(n878), .B2(n1539), .ZN(n1901)
         );
  INV_X1 U4028 ( .A(n1903), .ZN(n2605) );
  NOR2_X1 U4029 ( .A1(n1284), .A2(n4054), .ZN(n1086) );
  AOI21_X1 U4030 ( .B1(n529), .B2(n3549), .A(n1462), .ZN(n2381) );
  NOR3_X1 U4031 ( .A1(n4987), .A2(n5047), .A3(n4672), .ZN(n3179) );
  AOI21_X1 U4033 ( .B1(n1310), .B2(n3405), .A(n1347), .ZN(n1313) );
  AOI211_X1 U4034 ( .C1(n1348), .C2(n1284), .A(n3478), .B(n3915), .ZN(n1347)
         );
  OR2_X1 U4035 ( .A1(n1246), .A2(n4405), .ZN(n1348) );
  OAI21_X1 U4036 ( .B1(n1283), .B2(n1309), .A(n1313), .ZN(n1002) );
  NAND3_X1 U4037 ( .A1(n4405), .A2(n3913), .A3(n1274), .ZN(n1272) );
  NAND3_X1 U4038 ( .A1(n1183), .A2(n4405), .A3(n1304), .ZN(n993) );
  NOR2_X1 U4039 ( .A1(n3225), .A2(n4029), .ZN(n2048) );
  NOR2_X1 U4040 ( .A1(n1000), .A2(n4140), .ZN(n1435) );
  INV_X1 U4041 ( .A(n2137), .ZN(n3460) );
  INV_X1 U4042 ( .A(n2141), .ZN(n3454) );
  OAI21_X1 U4043 ( .B1(n1624), .B2(n2662), .A(n2233), .ZN(n1700) );
  NAND2_X1 U4044 ( .A1(n4222), .A2(n4633), .ZN(n2662) );
  NAND4_X1 U4045 ( .A1(n3077), .A2(n1442), .A3(n270), .A4(n2262), .ZN(n3076)
         );
  NOR2_X1 U4046 ( .A1(n1283), .A2(n1284), .ZN(n1073) );
  NAND2_X1 U4047 ( .A1(n833), .A2(n1371), .ZN(n2083) );
  NAND2_X1 U4048 ( .A1(n809), .A2(n1371), .ZN(n2087) );
  OAI22_X1 U4049 ( .A1(n3873), .A2(n354), .B1(n3329), .B2(n3712), .ZN(n4457)
         );
  OAI22_X1 U4050 ( .A1(n4932), .A2(n1458), .B1(n1459), .B2(n5225), .ZN(n1443)
         );
  AOI22_X1 U4051 ( .A1(n1461), .A2(n1462), .B1(n1463), .B2(n4512), .ZN(n1459)
         );
  NOR2_X1 U4052 ( .A1(n1464), .A2(n516), .ZN(n1461) );
  NOR2_X1 U4053 ( .A1(n597), .A2(n4017), .ZN(n639) );
  INV_X1 U4054 ( .A(n601), .ZN(n4017) );
  NAND2_X1 U4055 ( .A1(n2201), .A2(n3634), .ZN(n2123) );
  OAI211_X1 U4056 ( .C1(n4932), .C2(n516), .A(n3706), .B(n2867), .ZN(n2861) );
  AOI21_X1 U4057 ( .B1(n7375), .B2(n254), .A(n2868), .ZN(n2867) );
  INV_X1 U4058 ( .A(n2870), .ZN(n3706) );
  AOI21_X1 U4059 ( .B1(n479), .B2(n3686), .A(n521), .ZN(n2868) );
  NOR2_X1 U4060 ( .A1(Tzfpw6[0]), .A2(n1890), .ZN(n1887) );
  OAI22_X1 U4061 ( .A1(n2895), .A2(n3714), .B1(n2896), .B2(n4602), .ZN(n2890)
         );
  AOI21_X1 U4062 ( .B1(n521), .B2(n4826), .A(n536), .ZN(n2896) );
  AOI22_X1 U4063 ( .A1(n474), .A2(n1974), .B1(n1663), .B2(n875), .ZN(n2895) );
  AOI21_X1 U4064 ( .B1(n1948), .B2(n4670), .A(n1607), .ZN(n1946) );
  AOI22_X1 U4065 ( .A1(n2571), .A2(n4826), .B1(n513), .B2(n1520), .ZN(n2570)
         );
  NAND2_X1 U4066 ( .A1(n118), .A2(n1371), .ZN(n1963) );
  NOR2_X1 U4067 ( .A1(n592), .A2(n622), .ZN(n644) );
  OAI21_X1 U4068 ( .B1(n4795), .B2(n1482), .A(n4364), .ZN(n2862) );
  NAND3_X1 U4069 ( .A1(n4555), .A2(n4670), .A3(n7514), .ZN(n4216) );
  INV_X1 U4070 ( .A(n1907), .ZN(n3625) );
  INV_X1 U4071 ( .A(n2106), .ZN(n2865) );
  NOR2_X1 U4072 ( .A1(n3197), .A2(n593), .ZN(n643) );
  OR3_X1 U4073 ( .A1(n1703), .A2(n7514), .A3(n4187), .ZN(n1702) );
  AOI21_X1 U4074 ( .B1(n1457), .B2(n473), .A(n1704), .ZN(n1703) );
  AOI22_X1 U4075 ( .A1(n1760), .A2(n1751), .B1(n1584), .B2(n2262), .ZN(n4217)
         );
  NAND3_X1 U4076 ( .A1(n433), .A2(n434), .A3(n435), .ZN(n411) );
  OAI222_X1 U4077 ( .A1(n523), .A2(n4610), .B1(n4237), .B2(n3714), .C1(n266), 
        .C2(n3860), .ZN(n434) );
  OAI21_X1 U4078 ( .B1(n3549), .B2(n3525), .A(n529), .ZN(n3524) );
  AND2_X1 U4079 ( .A1(n2233), .A2(n3249), .ZN(n2489) );
  OAI22_X1 U4080 ( .A1(n477), .A2(n3766), .B1(n2915), .B2(n4229), .ZN(n3249)
         );
  NOR2_X1 U4081 ( .A1(n4548), .A2(n529), .ZN(n1431) );
  AND2_X1 U4082 ( .A1(n3441), .A2(n1287), .ZN(n1070) );
  INV_X1 U4083 ( .A(n647), .ZN(n3191) );
  AOI21_X1 U4084 ( .B1(n598), .B2(n555), .A(n4022), .ZN(n647) );
  NAND3_X1 U4085 ( .A1(n237), .A2(n3549), .A3(n2894), .ZN(n4311) );
  INV_X1 U4086 ( .A(n472), .ZN(n4725) );
  NOR2_X1 U4087 ( .A1(n1183), .A2(n1345), .ZN(n1246) );
  NAND3_X1 U4088 ( .A1(n7514), .A2(n464), .A3(n1576), .ZN(n1720) );
  INV_X1 U4089 ( .A(n2192), .ZN(n3471) );
  INV_X1 U4090 ( .A(n2144), .ZN(n3473) );
  INV_X1 U4091 ( .A(n2112), .ZN(n3002) );
  INV_X1 U4092 ( .A(n610), .ZN(n3226) );
  NAND2_X1 U4093 ( .A1(n636), .A2(n662), .ZN(n605) );
  OAI21_X1 U4094 ( .B1(n1083), .B2(n4053), .A(n1085), .ZN(n1082) );
  INV_X1 U4095 ( .A(n1086), .ZN(n4053) );
  NAND2_X1 U4096 ( .A1(n2048), .A2(n4024), .ZN(n558) );
  NAND2_X1 U4097 ( .A1(n557), .A2(n558), .ZN(n657) );
  INV_X1 U4098 ( .A(n2562), .ZN(n3803) );
  NAND3_X1 U4099 ( .A1(n470), .A2(n4993), .A3(n2454), .ZN(n2453) );
  INV_X1 U4100 ( .A(n2108), .ZN(n3419) );
  AND2_X1 U4101 ( .A1(n1310), .A2(n1311), .ZN(n843) );
  NAND2_X1 U4102 ( .A1(n5294), .A2(n5293), .ZN(n2501) );
  INV_X1 U4103 ( .A(n1346), .ZN(n4301) );
  NAND2_X1 U4104 ( .A1(n3441), .A2(n1346), .ZN(n1282) );
  OR4_X1 U4105 ( .A1(n1756), .A2(n2275), .A3(n475), .A4(n7381), .ZN(n2917) );
  INV_X1 U4106 ( .A(n1391), .ZN(n4052) );
  INV_X1 U4107 ( .A(n1379), .ZN(n4117) );
  INV_X1 U4108 ( .A(n1245), .ZN(n3443) );
  OAI22_X1 U4109 ( .A1(n1246), .A2(n1247), .B1(n1248), .B2(n1249), .ZN(n1245)
         );
  NAND2_X1 U4110 ( .A1(n4054), .A2(n4406), .ZN(n1249) );
  INV_X1 U4111 ( .A(n3077), .ZN(n4189) );
  INV_X1 U4112 ( .A(n1886), .ZN(n2977) );
  OR3_X1 U4113 ( .A1(n3208), .A2(n4028), .A3(n2049), .ZN(n598) );
  INV_X1 U4114 ( .A(n2843), .ZN(n3707) );
  INV_X1 U4115 ( .A(n595), .ZN(n3197) );
  INV_X1 U4116 ( .A(n987), .ZN(n3405) );
  INV_X1 U4117 ( .A(n2045), .ZN(n3215) );
  INV_X1 U4118 ( .A(n2057), .ZN(n4018) );
  INV_X1 U4119 ( .A(n1344), .ZN(n3478) );
  INV_X1 U4120 ( .A(n2127), .ZN(n2972) );
  INV_X1 U4121 ( .A(n552), .ZN(n1826) );
  AND2_X1 U4122 ( .A1(n2048), .A2(n655), .ZN(n622) );
  AND2_X1 U4123 ( .A1(n1857), .A2(n3634), .ZN(n1854) );
  INV_X1 U4124 ( .A(n662), .ZN(n3203) );
  AOI21_X1 U4125 ( .B1(n595), .B2(n3205), .A(n4022), .ZN(n614) );
  INV_X1 U4126 ( .A(n592), .ZN(n3205) );
  NAND2_X1 U4127 ( .A1(n3201), .A2(n4024), .ZN(n2063) );
  INV_X1 U4128 ( .A(n1303), .ZN(n3397) );
  AOI221_X1 U4129 ( .B1(n843), .B2(n1304), .C1(n1183), .C2(n3405), .A(n998), 
        .ZN(n1303) );
  INV_X1 U4130 ( .A(n1310), .ZN(n4330) );
  INV_X1 U4131 ( .A(n1290), .ZN(n3915) );
  INV_X1 U4132 ( .A(n557), .ZN(n3216) );
  INV_X1 U4133 ( .A(n3074), .ZN(n3684) );
  INV_X1 U4134 ( .A(n2149), .ZN(n4115) );
  NAND3_X1 U4135 ( .A1(n2058), .A2(n2059), .A3(n2060), .ZN(n8054) );
  OAI211_X1 U4137 ( .C1(n3223), .C2(n2063), .A(n4016), .B(n609), .ZN(n2058) );
  AOI22_X1 U4138 ( .A1(n666), .A2(n4028), .B1(n636), .B2(n4022), .ZN(n2060) );
  OAI211_X1 U4139 ( .C1(n2061), .C2(n2046), .A(n4024), .B(n648), .ZN(n2059) );
  INV_X1 U4140 ( .A(n603), .ZN(n3143) );
  BUF_X1 U4141 ( .A(n2103), .Z(n799) );
  INV_X1 U4142 ( .A(n1494), .ZN(n4588) );
  BUF_X1 U4143 ( .A(Fmdhu6), .Z(n956) );
  OAI221_X1 U4144 ( .B1(n4078), .B2(n4259), .C1(n7393), .C2(n2757), .A(n5100), 
        .ZN(n5099) );
  AOI22_X1 U4145 ( .A1(n4626), .A2(n5299), .B1(n4833), .B2(n5074), .ZN(n5100)
         );
  OAI22_X1 U4146 ( .A1(n3885), .A2(n4259), .B1(n7529), .B2(n4260), .ZN(n4392)
         );
  OAI221_X1 U4147 ( .B1(n3773), .B2(n4259), .C1(n7329), .C2(n2757), .A(n4832), 
        .ZN(n4831) );
  AOI22_X1 U4148 ( .A1(n4626), .A2(n5294), .B1(n4833), .B2(n5299), .ZN(n4832)
         );
  OAI221_X1 U4149 ( .B1(n7530), .B2(n4260), .C1(n3881), .C2(n4259), .A(n4625), 
        .ZN(n4624) );
  AOI22_X1 U4150 ( .A1(n4424), .A2(n4908), .B1(n4626), .B2(n5293), .ZN(n4625)
         );
  OAI22_X1 U4151 ( .A1(n659), .A2(n4940), .B1(n5181), .B2(n5182), .ZN(n3792)
         );
  OAI211_X1 U4152 ( .C1(n4176), .C2(n8112), .A(n2365), .B(n5183), .ZN(n5182)
         );
  OAI221_X1 U4153 ( .B1(n640), .B2(n4181), .C1(n2468), .C2(n6264), .A(n5184), 
        .ZN(n5181) );
  AOI222_X1 U4154 ( .A1(vis_r8_o[7]), .A2(n2336), .B1(vis_msp_o[5]), .B2(n2474), .C1(vis_r9_o[7]), .C2(n2338), .ZN(n5183) );
  OAI222_X1 U4155 ( .A1(n3873), .A2(n4259), .B1(n7326), .B2(n4260), .C1(n7359), 
        .C2(n2757), .ZN(n4257) );
  OAI221_X1 U4156 ( .B1(n3797), .B2(n3900), .C1(n1544), .C2(n661), .A(n3905), 
        .ZN(n199) );
  NAND2_X1 U4157 ( .A1(N5fpw6[30]), .A2(n669), .ZN(n3905) );
  NAND3_X1 U4158 ( .A1(n7343), .A2(n7284), .A3(n5722), .ZN(n4502) );
  OAI22_X1 U4159 ( .A1(n660), .A2(n4348), .B1(n4286), .B2(n4287), .ZN(n3811)
         );
  OAI211_X1 U4160 ( .C1(n4288), .C2(n8078), .A(n2458), .B(n4289), .ZN(n4287)
         );
  OAI221_X1 U4161 ( .B1(n646), .B2(n8129), .C1(n4291), .C2(n7922), .A(n4292), 
        .ZN(n4286) );
  AOI22_X1 U4162 ( .A1(vis_r12_o[1]), .A2(n4290), .B1(vis_r9_o[1]), .B2(n2338), 
        .ZN(n4289) );
  OAI22_X1 U4163 ( .A1(n659), .A2(n8167), .B1(n5719), .B2(n5720), .ZN(n3795)
         );
  OAI211_X1 U4164 ( .C1(n4176), .C2(n8124), .A(n2355), .B(n5721), .ZN(n5720)
         );
  OAI221_X1 U4165 ( .B1(n640), .B2(n3592), .C1(n2468), .C2(n2777), .A(n5727), 
        .ZN(n5719) );
  AOI222_X1 U4166 ( .A1(vis_r8_o[4]), .A2(n2336), .B1(vis_msp_o[2]), .B2(n2474), .C1(vis_r9_o[4]), .C2(n2338), .ZN(n5721) );
  OAI22_X1 U4167 ( .A1(n659), .A2(n8082), .B1(n5095), .B2(n5096), .ZN(n3794)
         );
  OAI211_X1 U4168 ( .C1(n4176), .C2(n4109), .A(n2347), .B(n5097), .ZN(n5096)
         );
  OAI221_X1 U4169 ( .B1(n640), .B2(n4086), .C1(n2468), .C2(n6229), .A(n5098), 
        .ZN(n5095) );
  AOI222_X1 U4170 ( .A1(vis_r8_o[5]), .A2(n2336), .B1(vis_msp_o[3]), .B2(n2474), .C1(vis_r9_o[5]), .C2(n2338), .ZN(n5097) );
  NOR2_X1 U4171 ( .A1(n5302), .A2(n7343), .ZN(n5723) );
  AOI22_X1 U4172 ( .A1(n650), .A2(n6676), .B1(n660), .B2(n4387), .ZN(n3822) );
  NAND2_X1 U4173 ( .A1(n4388), .A2(n4389), .ZN(n4387) );
  AOI221_X1 U4174 ( .B1(n2338), .B2(vis_r9_o[0]), .C1(n2336), .C2(vis_r8_o[0]), 
        .A(n4391), .ZN(n4388) );
  AOI221_X1 U4175 ( .B1(n2473), .B2(vis_r14_o[0]), .C1(n4290), .C2(
        vis_r12_o[0]), .A(n4390), .ZN(n4389) );
  OAI22_X1 U4176 ( .A1(n659), .A2(n8111), .B1(n4827), .B2(n4828), .ZN(n3796)
         );
  OAI211_X1 U4177 ( .C1(n4176), .C2(n8110), .A(n2460), .B(n4829), .ZN(n4828)
         );
  OAI221_X1 U4178 ( .B1(n640), .B2(n3774), .C1(n2468), .C2(n6260), .A(n4830), 
        .ZN(n4827) );
  AOI222_X1 U4179 ( .A1(vis_r8_o[3]), .A2(n2336), .B1(vis_msp_o[1]), .B2(n2474), .C1(vis_r9_o[3]), .C2(n2338), .ZN(n4829) );
  NOR2_X1 U4180 ( .A1(n7330), .A2(n7274), .ZN(n5770) );
  OAI22_X1 U4182 ( .A1(n7545), .A2(n660), .B1(n650), .B2(n4619), .ZN(n2709) );
  NOR3_X1 U4183 ( .A1(n4620), .A2(n4621), .A3(n4622), .ZN(n4619) );
  OAI22_X1 U4184 ( .A1(n4288), .A2(n8076), .B1(n4291), .B2(n8074), .ZN(n4622)
         );
  OAI222_X1 U4185 ( .A1(n4502), .A2(n5832), .B1(n4503), .B2(n6138), .C1(n646), 
        .C2(n8117), .ZN(n4621) );
  NOR4_X1 U4186 ( .A1(n3827), .A2(n2880), .A3(n7279), .A4(n3466), .ZN(n3826)
         );
  OAI21_X1 U4187 ( .B1(n491), .B2(n3173), .A(n3713), .ZN(n3827) );
  OAI21_X1 U4188 ( .B1(n7279), .B2(n5747), .A(n4452), .ZN(n4626) );
  AOI221_X1 U4189 ( .B1(n5753), .B2(n524), .C1(n4303), .C2(n266), .A(n5754), 
        .ZN(n5747) );
  AOI21_X1 U4190 ( .B1(n2754), .B2(n5755), .A(n7283), .ZN(n5753) );
  OAI22_X1 U4191 ( .A1(n477), .A2(n4193), .B1(n4265), .B2(n3732), .ZN(n5754)
         );
  NOR2_X1 U4193 ( .A1(n2466), .A2(n7520), .ZN(n5722) );
  NOR2_X1 U4194 ( .A1(n7520), .A2(n7382), .ZN(n5724) );
  AOI221_X1 U4195 ( .B1(vis_r14_o[7]), .B2(n2473), .C1(vis_r10_o[7]), .C2(
        n2322), .A(n650), .ZN(n5184) );
  AOI221_X1 U4196 ( .B1(vis_r14_o[3]), .B2(n2473), .C1(vis_r10_o[3]), .C2(
        n2322), .A(n654), .ZN(n4830) );
  AOI221_X1 U4198 ( .B1(vis_r14_o[4]), .B2(n2473), .C1(vis_r10_o[4]), .C2(
        n2322), .A(n654), .ZN(n5727) );
  AOI221_X1 U4199 ( .B1(vis_r14_o[5]), .B2(n2473), .C1(vis_r10_o[5]), .C2(
        n2322), .A(n650), .ZN(n5098) );
  NOR2_X1 U4200 ( .A1(n5304), .A2(n7284), .ZN(n5728) );
  NOR2_X1 U4201 ( .A1(n5312), .A2(n7360), .ZN(n5769) );
  NAND2_X1 U4202 ( .A1(n6510), .A2(n6511), .ZN(n5019) );
  AOI221_X1 U4203 ( .B1(vis_r5_o[1]), .B2(n582), .C1(vis_r4_o[1]), .C2(n581), 
        .A(n6512), .ZN(n6511) );
  AOI221_X1 U4204 ( .B1(vis_r6_o[1]), .B2(n576), .C1(vis_r1_o[1]), .C2(n575), 
        .A(n6513), .ZN(n6510) );
  OAI22_X1 U4205 ( .A1(n578), .A2(n4352), .B1(n4871), .B2(n6351), .ZN(n6512)
         );
  NOR4_X1 U4206 ( .A1(n428), .A2(n5731), .A3(n5732), .A4(n5733), .ZN(n4173) );
  OAI221_X1 U4207 ( .B1(n3714), .B2(n3232), .C1(n237), .C2(n3764), .A(n5734), 
        .ZN(n5733) );
  NOR3_X1 U4208 ( .A1(n3726), .A2(n7373), .A3(n272), .ZN(n5731) );
  AOI221_X1 U4209 ( .B1(n2730), .B2(n4519), .C1(n4424), .C2(n4987), .A(n4520), 
        .ZN(n4518) );
  OAI22_X1 U4210 ( .A1(n7527), .A2(n2546), .B1(n7400), .B2(n4452), .ZN(n4520)
         );
  NOR2_X1 U4211 ( .A1(n5313), .A2(n7394), .ZN(n5911) );
  NOR2_X1 U4212 ( .A1(n7360), .A2(n7394), .ZN(n5913) );
  OAI21_X1 U4213 ( .B1(n5761), .B2(n7279), .A(n4451), .ZN(n4833) );
  AOI222_X1 U4214 ( .A1(n5013), .A2(n5762), .B1(n529), .B2(n5763), .C1(n237), 
        .C2(n5764), .ZN(n5761) );
  OAI21_X1 U4215 ( .B1(n7373), .B2(n3732), .A(n3833), .ZN(n5763) );
  OAI21_X1 U4216 ( .B1(n228), .B2(n538), .A(n4245), .ZN(n5762) );
  NAND4_X1 U4217 ( .A1(n7343), .A2(n7520), .A3(n7284), .A4(n2466), .ZN(n6007)
         );
  NOR2_X1 U4218 ( .A1(n5291), .A2(n7330), .ZN(n6517) );
  NOR3_X1 U4219 ( .A1(n7343), .A2(n7284), .A3(n5307), .ZN(n6523) );
  NAND4_X1 U4220 ( .A1(n2618), .A2(n4989), .A3(n4990), .A4(n4991), .ZN(n4821)
         );
  NAND2_X1 U4221 ( .A1(n4864), .A2(n8111), .ZN(n4989) );
  AOI222_X1 U4222 ( .A1(vis_r10_o[3]), .A2(n617), .B1(vis_r11_o[3]), .B2(n4862), .C1(vis_r9_o[3]), .C2(n602), .ZN(n4990) );
  AOI221_X1 U4223 ( .B1(vis_r14_o[3]), .B2(n468), .C1(vis_r8_o[3]), .C2(n628), 
        .A(n4992), .ZN(n4991) );
  OAI221_X1 U4224 ( .B1(n7400), .B2(n2546), .C1(n3956), .C2(n4259), .A(n5746), 
        .ZN(n5740) );
  AOI22_X1 U4225 ( .A1(n4424), .A2(n4932), .B1(n4626), .B2(n3083), .ZN(n5746)
         );
  NAND3_X1 U4226 ( .A1(n5723), .A2(n2466), .A3(n7520), .ZN(n6006) );
  NAND3_X1 U4227 ( .A1(n7401), .A2(n5769), .A3(n5770), .ZN(n4859) );
  NAND3_X1 U4228 ( .A1(n7520), .A2(n5723), .A3(n7382), .ZN(n6002) );
  NAND3_X1 U4230 ( .A1(n7520), .A2(n2466), .A3(n5728), .ZN(n6001) );
  OAI211_X1 U4231 ( .C1(n4504), .C2(n5976), .A(n2462), .B(n4623), .ZN(n4620)
         );
  AOI22_X1 U4232 ( .A1(vis_psp_o[0]), .A2(n229), .B1(vis_r12_o[2]), .B2(n4290), 
        .ZN(n4623) );
  NAND2_X1 U4233 ( .A1(n6016), .A2(n6017), .ZN(n5281) );
  AOI221_X1 U4234 ( .B1(n561), .B2(vis_r2_o[1]), .C1(n550), .C2(vis_r0_o[1]), 
        .A(n6019), .ZN(n6016) );
  AOI221_X1 U4235 ( .B1(n5998), .B2(vis_r3_o[1]), .C1(n565), .C2(vis_r7_o[1]), 
        .A(n6018), .ZN(n6017) );
  OAI22_X1 U4236 ( .A1(n6479), .A2(n541), .B1(n5403), .B2(n540), .ZN(n6019) );
  AND4_X1 U4237 ( .A1(n4351), .A2(n5014), .A3(n5015), .A4(n5016), .ZN(n3873)
         );
  NAND2_X1 U4238 ( .A1(n4864), .A2(n4348), .ZN(n5014) );
  AOI22_X1 U4239 ( .A1(vis_r9_o[1]), .A2(n4863), .B1(vis_r10_o[1]), .B2(n4861), 
        .ZN(n5015) );
  AOI221_X1 U4240 ( .B1(vis_r8_o[1]), .B2(n628), .C1(vis_r11_o[1]), .C2(n615), 
        .A(n5017), .ZN(n5016) );
  AND4_X1 U4241 ( .A1(n2643), .A2(n5906), .A3(n5907), .A4(n5908), .ZN(n3885)
         );
  NAND2_X1 U4242 ( .A1(n6676), .A2(n599), .ZN(n5906) );
  AOI22_X1 U4243 ( .A1(vis_r9_o[0]), .A2(n4863), .B1(vis_r10_o[0]), .B2(n4861), 
        .ZN(n5907) );
  AOI221_X1 U4244 ( .B1(vis_r8_o[0]), .B2(n628), .C1(vis_r11_o[0]), .C2(n615), 
        .A(n5909), .ZN(n5908) );
  NAND3_X1 U4245 ( .A1(n5910), .A2(n7274), .A3(n7330), .ZN(n4871) );
  NAND3_X1 U4246 ( .A1(n7330), .A2(n7274), .A3(n5913), .ZN(n4870) );
  NAND3_X1 U4247 ( .A1(n7330), .A2(n7274), .A3(n5911), .ZN(n4876) );
  AOI21_X1 U4248 ( .B1(vis_r8_o[1]), .B2(n2336), .A(n654), .ZN(n4292) );
  AND4_X1 U4249 ( .A1(n2621), .A2(n4974), .A3(n4975), .A4(n4976), .ZN(n3881)
         );
  NAND2_X1 U4250 ( .A1(n599), .A2(n8168), .ZN(n4974) );
  AOI222_X1 U4251 ( .A1(vis_r10_o[2]), .A2(n4861), .B1(vis_r11_o[2]), .B2(
        n4862), .C1(vis_r9_o[2]), .C2(n602), .ZN(n4975) );
  AOI221_X1 U4252 ( .B1(vis_r14_o[2]), .B2(n468), .C1(vis_r8_o[2]), .C2(n628), 
        .A(n4977), .ZN(n4976) );
  NAND2_X1 U4253 ( .A1(n6012), .A2(n6013), .ZN(n4390) );
  AOI221_X1 U4254 ( .B1(n561), .B2(vis_r2_o[0]), .C1(n550), .C2(vis_r0_o[0]), 
        .A(n6015), .ZN(n6012) );
  AOI221_X1 U4255 ( .B1(n5998), .B2(vis_r3_o[0]), .C1(n565), .C2(vis_r7_o[0]), 
        .A(n6014), .ZN(n6013) );
  OAI22_X1 U4256 ( .A1(n3343), .A2(n541), .B1(n5366), .B2(n540), .ZN(n6015) );
  NAND2_X1 U4257 ( .A1(n5996), .A2(n5997), .ZN(n5492) );
  AOI221_X1 U4258 ( .B1(n561), .B2(vis_r2_o[2]), .C1(n550), .C2(vis_r0_o[2]), 
        .A(n6005), .ZN(n5996) );
  AOI221_X1 U4260 ( .B1(n5998), .B2(vis_r3_o[2]), .C1(n565), .C2(vis_r7_o[2]), 
        .A(n6000), .ZN(n5997) );
  OAI22_X1 U4261 ( .A1(n6537), .A2(n541), .B1(n5464), .B2(n540), .ZN(n6005) );
  AND3_X1 U4262 ( .A1(n5769), .A2(n7274), .A3(n7330), .ZN(n4873) );
  AND3_X1 U4263 ( .A1(n7382), .A2(n7520), .A3(n5728), .ZN(n6003) );
  INV_X1 U4264 ( .A(n4617), .ZN(Qbfpw6_2) );
  NOR3_X1 U4265 ( .A1(n3799), .A2(n3789), .A3(n2330), .ZN(Idfpw6[2]) );
  NOR3_X1 U4266 ( .A1(n3805), .A2(n7279), .A3(n522), .ZN(n3799) );
  AND2_X1 U4267 ( .A1(n6514), .A2(n6515), .ZN(n2643) );
  AOI221_X1 U4268 ( .B1(vis_r5_o[0]), .B2(n582), .C1(vis_r4_o[0]), .C2(n581), 
        .A(n6516), .ZN(n6515) );
  AOI221_X1 U4269 ( .B1(vis_r6_o[0]), .B2(n576), .C1(vis_r1_o[0]), .C2(n575), 
        .A(n6519), .ZN(n6514) );
  OAI22_X1 U4270 ( .A1(n578), .A2(n7578), .B1(n4871), .B2(n6378), .ZN(n6516)
         );
  AND2_X1 U4271 ( .A1(n6488), .A2(n6489), .ZN(n2621) );
  AOI221_X1 U4272 ( .B1(vis_r5_o[2]), .B2(n582), .C1(vis_r4_o[2]), .C2(n581), 
        .A(n6490), .ZN(n6489) );
  AOI221_X1 U4273 ( .B1(vis_r6_o[2]), .B2(n576), .C1(vis_r1_o[2]), .C2(n575), 
        .A(n6491), .ZN(n6488) );
  OAI22_X1 U4274 ( .A1(n578), .A2(n7370), .B1(n577), .B2(n4273), .ZN(n6490) );
  AND2_X1 U4275 ( .A1(n6448), .A2(n6449), .ZN(n2618) );
  AOI221_X1 U4276 ( .B1(vis_r5_o[3]), .B2(n582), .C1(vis_r4_o[3]), .C2(n581), 
        .A(n6450), .ZN(n6449) );
  AOI221_X1 U4277 ( .B1(vis_r6_o[3]), .B2(n576), .C1(vis_r1_o[3]), .C2(n575), 
        .A(n6451), .ZN(n6448) );
  OAI22_X1 U4278 ( .A1(n578), .A2(n7668), .B1(n577), .B2(n6365), .ZN(n6450) );
  AND2_X1 U4279 ( .A1(n6523), .A2(n7382), .ZN(n5998) );
  AND2_X1 U4280 ( .A1(n7330), .A2(n5291), .ZN(n5912) );
  NOR2_X1 U4281 ( .A1(n7532), .A2(n4354), .ZN(n1430) );
  OAI221_X1 U4282 ( .B1(n2757), .B2(n7527), .C1(n4259), .C2(n3278), .A(n2597), 
        .ZN(n4798) );
  AOI22_X1 U4283 ( .A1(n650), .A2(n6679), .B1(n660), .B2(n4513), .ZN(n3793) );
  OR3_X1 U4284 ( .A1(n4514), .A2(n4515), .A3(n4516), .ZN(n4513) );
  OAI22_X1 U4285 ( .A1(n4288), .A2(n4280), .B1(n4291), .B2(n8070), .ZN(n4516)
         );
  OAI222_X1 U4286 ( .A1(n4502), .A2(n5894), .B1(n4503), .B2(n6039), .C1(n646), 
        .C2(n8122), .ZN(n4515) );
  NOR2_X1 U4287 ( .A1(n479), .A2(n7492), .ZN(n1566) );
  OAI22_X1 U4288 ( .A1(n659), .A2(n8177), .B1(n4427), .B2(n4428), .ZN(n3813)
         );
  OAI211_X1 U4289 ( .C1(n4176), .C2(n8187), .A(n2390), .B(n4429), .ZN(n4428)
         );
  OAI221_X1 U4290 ( .B1(n640), .B2(n8184), .C1(n2468), .C2(n8181), .A(n4430), 
        .ZN(n4427) );
  AOI222_X1 U4291 ( .A1(vis_r8_o[18]), .A2(n2336), .B1(vis_msp_o[16]), .B2(
        n2474), .C1(vis_r9_o[18]), .C2(n2338), .ZN(n4429) );
  OAI22_X1 U4292 ( .A1(n659), .A2(n8224), .B1(n5610), .B2(n5611), .ZN(n3812)
         );
  OAI211_X1 U4293 ( .C1(n646), .C2(n3865), .A(n2400), .B(n5612), .ZN(n5611) );
  OAI221_X1 U4294 ( .B1(n640), .B2(n3864), .C1(n2468), .C2(n6239), .A(n5613), 
        .ZN(n5610) );
  AOI222_X1 U4295 ( .A1(vis_r8_o[19]), .A2(n2336), .B1(vis_msp_o[17]), .B2(
        n2474), .C1(vis_r9_o[19]), .C2(n2338), .ZN(n5612) );
  OAI22_X1 U4296 ( .A1(n659), .A2(n8116), .B1(n4483), .B2(n4484), .ZN(n3816)
         );
  OAI211_X1 U4297 ( .C1(n4176), .C2(n8115), .A(n2413), .B(n4485), .ZN(n4484)
         );
  OAI221_X1 U4298 ( .B1(n640), .B2(n3583), .C1(n2468), .C2(n2490), .A(n4486), 
        .ZN(n4483) );
  AOI222_X1 U4299 ( .A1(vis_r8_o[15]), .A2(n2336), .B1(vis_msp_o[13]), .B2(
        n2474), .C1(vis_r9_o[15]), .C2(n2338), .ZN(n4485) );
  OAI22_X1 U4300 ( .A1(n660), .A2(n4185), .B1(n5075), .B2(n5076), .ZN(n3815)
         );
  OAI211_X1 U4301 ( .C1(n4176), .C2(n8128), .A(n2397), .B(n5077), .ZN(n5076)
         );
  OAI221_X1 U4302 ( .B1(n640), .B2(n4003), .C1(n2468), .C2(n6218), .A(n5078), 
        .ZN(n5075) );
  AOI222_X1 U4303 ( .A1(vis_r8_o[16]), .A2(n2336), .B1(vis_msp_o[14]), .B2(
        n2474), .C1(vis_r9_o[16]), .C2(n2338), .ZN(n5077) );
  NAND3_X1 U4304 ( .A1(n5724), .A2(n5723), .A3(n7401), .ZN(n4504) );
  NOR2_X1 U4305 ( .A1(n476), .A2(n7510), .ZN(n1907) );
  NOR2_X1 U4306 ( .A1(n4635), .A2(n7399), .ZN(n3077) );
  OAI211_X1 U4307 ( .C1(n439), .C2(n1544), .A(n4325), .B(n4326), .ZN(n3409) );
  AOI22_X1 U4308 ( .A1(n2551), .A2(n3458), .B1(vis_apsr_o[3]), .B2(n4342), 
        .ZN(n4325) );
  AOI211_X1 U4309 ( .C1(n4327), .C2(n4328), .A(n635), .B(Affpw6[31]), .ZN(
        n4326) );
  NAND3_X1 U4310 ( .A1(n2550), .A2(D5epw6), .A3(n2280), .ZN(n4328) );
  NOR2_X1 U4311 ( .A1(n4670), .A2(n7505), .ZN(n2585) );
  NAND4_X1 U4312 ( .A1(n2637), .A2(n4898), .A3(n4899), .A4(n4900), .ZN(n4471)
         );
  NAND2_X1 U4313 ( .A1(n599), .A2(n8116), .ZN(n4898) );
  AOI222_X1 U4314 ( .A1(vis_r10_o[15]), .A2(n617), .B1(vis_r11_o[15]), .B2(
        n4862), .C1(vis_r9_o[15]), .C2(n602), .ZN(n4899) );
  AOI221_X1 U4315 ( .B1(vis_r14_o[15]), .B2(n5272), .C1(vis_r8_o[15]), .C2(
        n628), .A(n4901), .ZN(n4900) );
  NOR2_X1 U4316 ( .A1(n4354), .A2(n7493), .ZN(n1977) );
  AOI221_X1 U4317 ( .B1(vis_r14_o[10]), .B2(n2473), .C1(vis_r10_o[10]), .C2(
        n2322), .A(n654), .ZN(n4746) );
  AOI221_X1 U4318 ( .B1(vis_r14_o[11]), .B2(n2473), .C1(vis_r10_o[11]), .C2(
        n2322), .A(n650), .ZN(n5588) );
  AOI221_X1 U4319 ( .B1(vis_r14_o[14]), .B2(n2473), .C1(vis_r10_o[14]), .C2(
        n2322), .A(n650), .ZN(n5138) );
  AOI221_X1 U4320 ( .B1(vis_r14_o[8]), .B2(n2473), .C1(vis_r10_o[8]), .C2(
        n2322), .A(n654), .ZN(n5051) );
  AOI221_X1 U4321 ( .B1(vis_r14_o[13]), .B2(n2473), .C1(vis_r10_o[13]), .C2(
        n2322), .A(n650), .ZN(n5356) );
  AOI221_X1 U4322 ( .B1(vis_r14_o[12]), .B2(n2473), .C1(vis_r10_o[12]), .C2(
        n2322), .A(n654), .ZN(n4647) );
  AOI221_X1 U4323 ( .B1(vis_r14_o[18]), .B2(n2473), .C1(vis_r10_o[18]), .C2(
        n2322), .A(n654), .ZN(n4430) );
  AOI221_X1 U4324 ( .B1(vis_r14_o[19]), .B2(n2473), .C1(vis_r10_o[19]), .C2(
        n2322), .A(n650), .ZN(n5613) );
  AOI221_X1 U4325 ( .B1(vis_r14_o[15]), .B2(n2473), .C1(vis_r10_o[15]), .C2(
        n2322), .A(n654), .ZN(n4486) );
  AOI221_X1 U4326 ( .B1(vis_r14_o[17]), .B2(n2473), .C1(vis_r10_o[17]), .C2(
        n2322), .A(n650), .ZN(n5632) );
  AOI221_X1 U4327 ( .B1(vis_r14_o[16]), .B2(n2473), .C1(vis_r10_o[16]), .C2(
        n2322), .A(n654), .ZN(n5078) );
  NAND2_X1 U4328 ( .A1(n6093), .A2(n6094), .ZN(n5323) );
  AOI221_X1 U4329 ( .B1(vis_r2_o[13]), .B2(n6003), .C1(vis_r0_o[13]), .C2(n547), .A(n6096), .ZN(n6093) );
  AOI221_X1 U4330 ( .B1(vis_r3_o[13]), .B2(n567), .C1(vis_r7_o[13]), .C2(n5999), .A(n6095), .ZN(n6094) );
  OAI22_X1 U4331 ( .A1(n6006), .A2(n6595), .B1(n6007), .B2(n5334), .ZN(n6096)
         );
  NAND2_X1 U4332 ( .A1(n6469), .A2(n6470), .ZN(n5536) );
  AOI221_X1 U4333 ( .B1(vis_r2_o[8]), .B2(n561), .C1(vis_r0_o[8]), .C2(n547), 
        .A(n6472), .ZN(n6469) );
  AOI221_X1 U4334 ( .B1(vis_r3_o[8]), .B2(n567), .C1(vis_r7_o[8]), .C2(n565), 
        .A(n6471), .ZN(n6470) );
  OAI22_X1 U4335 ( .A1(n541), .A2(n6399), .B1(n540), .B2(n5370), .ZN(n6472) );
  NAND2_X1 U4336 ( .A1(n6085), .A2(n6086), .ZN(n5984) );
  AOI221_X1 U4337 ( .B1(vis_r2_o[15]), .B2(n6003), .C1(vis_r0_o[15]), .C2(n547), .A(n6088), .ZN(n6085) );
  AOI221_X1 U4338 ( .B1(vis_r3_o[15]), .B2(n567), .C1(vis_r7_o[15]), .C2(n5999), .A(n6087), .ZN(n6086) );
  OAI22_X1 U4339 ( .A1(n6006), .A2(n6585), .B1(n6007), .B2(n5317), .ZN(n6088)
         );
  NAND2_X1 U4340 ( .A1(n6089), .A2(n6090), .ZN(n4646) );
  AOI221_X1 U4341 ( .B1(vis_r2_o[12]), .B2(n6003), .C1(vis_r0_o[12]), .C2(n547), .A(n6092), .ZN(n6089) );
  AOI221_X1 U4342 ( .B1(vis_r3_o[12]), .B2(n567), .C1(vis_r7_o[12]), .C2(n5999), .A(n6091), .ZN(n6090) );
  OAI22_X1 U4343 ( .A1(n6006), .A2(n6526), .B1(n6007), .B2(n5449), .ZN(n6092)
         );
  NAND2_X1 U4344 ( .A1(n6457), .A2(n6458), .ZN(n5340) );
  AOI221_X1 U4345 ( .B1(vis_r2_o[11]), .B2(n6003), .C1(vis_r0_o[11]), .C2(n547), .A(n6460), .ZN(n6457) );
  AOI221_X1 U4346 ( .B1(vis_r3_o[11]), .B2(n567), .C1(vis_r7_o[11]), .C2(n5999), .A(n6459), .ZN(n6458) );
  OAI22_X1 U4347 ( .A1(n6006), .A2(n6425), .B1(n6007), .B2(n5372), .ZN(n6460)
         );
  XNOR2_X1 U4348 ( .A(n2545), .B(n5052), .ZN(W4epw6) );
  AOI221_X1 U4349 ( .B1(n2730), .B2(n4955), .C1(n4424), .C2(n4670), .A(n5053), 
        .ZN(n5052) );
  OAI22_X1 U4350 ( .A1(n7524), .A2(n4451), .B1(n7527), .B2(n4452), .ZN(n5053)
         );
  XNOR2_X1 U4351 ( .A(n2545), .B(n5185), .ZN(S2epw6) );
  AOI221_X1 U4352 ( .B1(n2730), .B2(n5186), .C1(n4424), .C2(n4993), .A(n5187), 
        .ZN(n5185) );
  OAI22_X1 U4353 ( .A1(n7506), .A2(n2546), .B1(n7356), .B2(n4452), .ZN(n5187)
         );
  XNOR2_X1 U4354 ( .A(n2545), .B(n4448), .ZN(Q5phu6) );
  AOI221_X1 U4355 ( .B1(n2730), .B2(n4449), .C1(n4424), .C2(n464), .A(n4450), 
        .ZN(n4448) );
  OAI22_X1 U4356 ( .A1(n7525), .A2(n4451), .B1(n7506), .B2(n4452), .ZN(n4450)
         );
  NAND4_X1 U4357 ( .A1(n2639), .A2(n5358), .A3(n5359), .A4(n5360), .ZN(n4878)
         );
  NAND2_X1 U4358 ( .A1(n4864), .A2(n3041), .ZN(n5358) );
  AOI222_X1 U4359 ( .A1(vis_r10_o[13]), .A2(n617), .B1(vis_r11_o[13]), .B2(
        n4862), .C1(vis_r9_o[13]), .C2(n602), .ZN(n5359) );
  AOI221_X1 U4360 ( .B1(vis_r14_o[13]), .B2(n5272), .C1(vis_r8_o[13]), .C2(
        n4856), .A(n5361), .ZN(n5360) );
  NAND2_X1 U4361 ( .A1(n6437), .A2(n6438), .ZN(n5550) );
  AOI221_X1 U4362 ( .B1(vis_r5_o[5]), .B2(n582), .C1(vis_r4_o[5]), .C2(n581), 
        .A(n6439), .ZN(n6438) );
  AOI221_X1 U4363 ( .B1(vis_r6_o[5]), .B2(n576), .C1(vis_r1_o[5]), .C2(n575), 
        .A(n6440), .ZN(n6437) );
  OAI22_X1 U4364 ( .A1(n578), .A2(n7600), .B1(n4871), .B2(n6331), .ZN(n6439)
         );
  NAND2_X1 U4365 ( .A1(n6426), .A2(n6427), .ZN(n5771) );
  AOI221_X1 U4366 ( .B1(vis_r5_o[4]), .B2(n582), .C1(vis_r4_o[4]), .C2(n581), 
        .A(n6428), .ZN(n6427) );
  AOI221_X1 U4367 ( .B1(vis_r6_o[4]), .B2(n576), .C1(vis_r1_o[4]), .C2(n575), 
        .A(n6429), .ZN(n6426) );
  OAI22_X1 U4368 ( .A1(n578), .A2(n7575), .B1(n577), .B2(n6349), .ZN(n6428) );
  NAND2_X1 U4369 ( .A1(n6433), .A2(n6434), .ZN(n4562) );
  AOI221_X1 U4370 ( .B1(vis_r5_o[6]), .B2(n582), .C1(vis_r4_o[6]), .C2(n581), 
        .A(n6435), .ZN(n6434) );
  AOI221_X1 U4371 ( .B1(vis_r6_o[6]), .B2(n576), .C1(vis_r1_o[6]), .C2(n575), 
        .A(n6436), .ZN(n6433) );
  OAI22_X1 U4372 ( .A1(n578), .A2(n7376), .B1(n4871), .B2(n6294), .ZN(n6435)
         );
  NAND2_X1 U4373 ( .A1(n6441), .A2(n6442), .ZN(n4563) );
  AOI221_X1 U4374 ( .B1(vis_r5_o[7]), .B2(n582), .C1(vis_r4_o[7]), .C2(n581), 
        .A(n6443), .ZN(n6442) );
  AOI221_X1 U4375 ( .B1(vis_r6_o[7]), .B2(n576), .C1(vis_r1_o[7]), .C2(n575), 
        .A(n6444), .ZN(n6441) );
  OAI22_X1 U4376 ( .A1(n578), .A2(n7695), .B1(n4871), .B2(n6377), .ZN(n6443)
         );
  NAND4_X1 U4377 ( .A1(n2640), .A2(n4852), .A3(n4853), .A4(n4854), .ZN(n4649)
         );
  NAND2_X1 U4378 ( .A1(n4864), .A2(n8103), .ZN(n4852) );
  AOI222_X1 U4379 ( .A1(vis_r10_o[12]), .A2(n617), .B1(vis_r11_o[12]), .B2(
        n615), .C1(vis_r9_o[12]), .C2(n4863), .ZN(n4853) );
  AOI221_X1 U4380 ( .B1(vis_r14_o[12]), .B2(n5272), .C1(vis_r8_o[12]), .C2(
        n4856), .A(n4857), .ZN(n4854) );
  NAND4_X1 U4381 ( .A1(n2641), .A2(n5590), .A3(n5591), .A4(n5592), .ZN(n4938)
         );
  NAND2_X1 U4382 ( .A1(n4864), .A2(n8163), .ZN(n5590) );
  AOI222_X1 U4383 ( .A1(vis_r10_o[11]), .A2(n617), .B1(vis_r11_o[11]), .B2(
        n615), .C1(vis_r9_o[11]), .C2(n4863), .ZN(n5591) );
  AOI221_X1 U4384 ( .B1(vis_r14_o[11]), .B2(n5272), .C1(vis_r8_o[11]), .C2(
        n4856), .A(n5593), .ZN(n5592) );
  NAND4_X1 U4385 ( .A1(n2638), .A2(n5140), .A3(n5141), .A4(n5142), .ZN(n4888)
         );
  NAND2_X1 U4386 ( .A1(n4864), .A2(n8252), .ZN(n5140) );
  AOI222_X1 U4387 ( .A1(vis_r10_o[14]), .A2(n617), .B1(vis_r11_o[14]), .B2(
        n615), .C1(vis_r9_o[14]), .C2(n4863), .ZN(n5141) );
  AOI221_X1 U4388 ( .B1(vis_r14_o[14]), .B2(n5272), .C1(vis_r8_o[14]), .C2(
        n4856), .A(n5143), .ZN(n5142) );
  NAND4_X1 U4389 ( .A1(n2612), .A2(n4928), .A3(n4929), .A4(n4930), .ZN(n4449)
         );
  NAND2_X1 U4390 ( .A1(n599), .A2(n8173), .ZN(n4928) );
  AOI222_X1 U4392 ( .A1(vis_r10_o[9]), .A2(n617), .B1(vis_r11_o[9]), .B2(n4862), .C1(vis_r9_o[9]), .C2(n602), .ZN(n4929) );
  AOI221_X1 U4393 ( .B1(vis_r14_o[9]), .B2(n468), .C1(vis_r8_o[9]), .C2(n4856), 
        .A(n4931), .ZN(n4930) );
  NAND4_X1 U4394 ( .A1(n2613), .A2(n5054), .A3(n5055), .A4(n5056), .ZN(n4955)
         );
  NAND2_X1 U4395 ( .A1(n4864), .A2(n4009), .ZN(n5054) );
  AOI222_X1 U4396 ( .A1(vis_r10_o[8]), .A2(n617), .B1(vis_r11_o[8]), .B2(n4862), .C1(vis_r9_o[8]), .C2(n602), .ZN(n5055) );
  AOI221_X1 U4397 ( .B1(vis_r14_o[8]), .B2(n468), .C1(vis_r8_o[8]), .C2(n4856), 
        .A(n5057), .ZN(n5056) );
  OAI22_X1 U4398 ( .A1(n7408), .A2(n659), .B1(n650), .B2(n5414), .ZN(n4447) );
  NOR3_X1 U4399 ( .A1(n5415), .A2(n5416), .A3(n5417), .ZN(n5414) );
  OAI22_X1 U4400 ( .A1(n4288), .A2(n8086), .B1(n4291), .B2(n8056), .ZN(n5417)
         );
  OAI222_X1 U4401 ( .A1(n4502), .A2(n5891), .B1(n4503), .B2(n6142), .C1(n646), 
        .C2(n8101), .ZN(n5416) );
  OAI222_X1 U4402 ( .A1(n7516), .A2(n2757), .B1(n3608), .B2(n4259), .C1(n7526), 
        .C2(n4451), .ZN(n4742) );
  OAI22_X1 U4403 ( .A1(n7332), .A2(n3459), .B1(n1542), .B2(n5257), .ZN(n2940)
         );
  INV_X1 U4404 ( .A(n3409), .ZN(n1542) );
  NAND4_X1 U4405 ( .A1(n7283), .A2(n4591), .A3(n4202), .A4(n3831), .ZN(n5221)
         );
  OAI22_X1 U4406 ( .A1(n659), .A2(n8171), .B1(n4743), .B2(n4744), .ZN(n3821)
         );
  OAI211_X1 U4407 ( .C1(n4176), .C2(n8113), .A(n2384), .B(n4745), .ZN(n4744)
         );
  OAI221_X1 U4408 ( .B1(n640), .B2(n3611), .C1(n2468), .C2(n6267), .A(n4746), 
        .ZN(n4743) );
  AOI222_X1 U4409 ( .A1(vis_r8_o[10]), .A2(n2336), .B1(vis_msp_o[8]), .B2(
        n2474), .C1(vis_r9_o[10]), .C2(n2338), .ZN(n4745) );
  OAI22_X1 U4410 ( .A1(n659), .A2(n8163), .B1(n5585), .B2(n5586), .ZN(n3820)
         );
  OAI211_X1 U4411 ( .C1(n646), .C2(n8126), .A(n2387), .B(n5587), .ZN(n5586) );
  OAI221_X1 U4412 ( .B1(n640), .B2(n3591), .C1(n2468), .C2(n6212), .A(n5588), 
        .ZN(n5585) );
  AOI222_X1 U4413 ( .A1(vis_r8_o[11]), .A2(n2336), .B1(vis_msp_o[9]), .B2(
        n2474), .C1(vis_r9_o[11]), .C2(n2338), .ZN(n5587) );
  OAI22_X1 U4414 ( .A1(n659), .A2(n8252), .B1(n5135), .B2(n5136), .ZN(n3817)
         );
  OAI211_X1 U4415 ( .C1(n4176), .C2(n8132), .A(n2403), .B(n5137), .ZN(n5136)
         );
  OAI221_X1 U4416 ( .B1(n640), .B2(n4167), .C1(n2468), .C2(n6225), .A(n5138), 
        .ZN(n5135) );
  AOI222_X1 U4417 ( .A1(vis_r8_o[14]), .A2(n2336), .B1(vis_msp_o[12]), .B2(
        n2474), .C1(vis_r9_o[14]), .C2(n2338), .ZN(n5137) );
  OAI22_X1 U4418 ( .A1(n659), .A2(n4009), .B1(n5048), .B2(n5049), .ZN(n3791)
         );
  OAI211_X1 U4419 ( .C1(n4176), .C2(n8125), .A(n2367), .B(n5050), .ZN(n5049)
         );
  OAI221_X1 U4422 ( .B1(n640), .B2(n4007), .C1(n2468), .C2(n6210), .A(n5051), 
        .ZN(n5048) );
  AOI222_X1 U4423 ( .A1(vis_r8_o[8]), .A2(n2336), .B1(vis_msp_o[6]), .B2(n2474), .C1(vis_r9_o[8]), .C2(n2338), .ZN(n5050) );
  OAI22_X1 U4424 ( .A1(n659), .A2(n3041), .B1(n5353), .B2(n5354), .ZN(n3818)
         );
  OAI211_X1 U4425 ( .C1(n4176), .C2(n8121), .A(n2406), .B(n5355), .ZN(n5354)
         );
  OAI221_X1 U4426 ( .B1(n640), .B2(n3588), .C1(n2468), .C2(n6183), .A(n5356), 
        .ZN(n5353) );
  AOI222_X1 U4427 ( .A1(vis_r8_o[13]), .A2(n2336), .B1(vis_msp_o[11]), .B2(
        n2474), .C1(vis_r9_o[13]), .C2(n2338), .ZN(n5355) );
  OAI22_X1 U4428 ( .A1(n659), .A2(n8103), .B1(n4643), .B2(n4644), .ZN(n3819)
         );
  OAI211_X1 U4429 ( .C1(n4176), .C2(n8102), .A(n2411), .B(n4645), .ZN(n4644)
         );
  OAI221_X1 U4430 ( .B1(n640), .B2(n4178), .C1(n2468), .C2(n6242), .A(n4647), 
        .ZN(n4643) );
  AOI222_X1 U4431 ( .A1(vis_r8_o[12]), .A2(n2336), .B1(vis_msp_o[10]), .B2(
        n2474), .C1(vis_r9_o[12]), .C2(n2338), .ZN(n4645) );
  OAI22_X1 U4432 ( .A1(n659), .A2(n3280), .B1(n5629), .B2(n5630), .ZN(n3814)
         );
  OAI211_X1 U4433 ( .C1(n646), .C2(n8109), .A(n2392), .B(n5631), .ZN(n5630) );
  OAI221_X1 U4434 ( .B1(n640), .B2(n3279), .C1(n2468), .C2(n6257), .A(n5632), 
        .ZN(n5629) );
  AOI222_X1 U4435 ( .A1(vis_r8_o[17]), .A2(n2336), .B1(vis_msp_o[15]), .B2(
        n2474), .C1(vis_r9_o[17]), .C2(n2338), .ZN(n5631) );
  OAI221_X1 U4436 ( .B1(n2905), .B2(n2726), .C1(n476), .C2(n2907), .A(n2908), 
        .ZN(n2900) );
  AOI22_X1 U4437 ( .A1(n88), .A2(n2909), .B1(n7492), .B2(n2910), .ZN(n2908) );
  AOI22_X1 U4438 ( .A1(n2920), .A2(n449), .B1(n2921), .B2(n2922), .ZN(n2905)
         );
  NAND3_X1 U4439 ( .A1(n2697), .A2(n2698), .A3(n2917), .ZN(n2909) );
  NAND4_X1 U4440 ( .A1(n2642), .A2(n4966), .A3(n4967), .A4(n4968), .ZN(n4747)
         );
  NAND2_X1 U4441 ( .A1(n599), .A2(n8171), .ZN(n4966) );
  AOI222_X1 U4442 ( .A1(vis_r10_o[10]), .A2(n617), .B1(vis_r11_o[10]), .B2(
        n4862), .C1(vis_r9_o[10]), .C2(n602), .ZN(n4967) );
  AOI221_X1 U4443 ( .B1(vis_r14_o[10]), .B2(n468), .C1(vis_r8_o[10]), .C2(
        n4856), .A(n4969), .ZN(n4968) );
  NAND4_X1 U4444 ( .A1(n5278), .A2(n4942), .A3(n4943), .A4(n4944), .ZN(n4519)
         );
  NAND2_X1 U4445 ( .A1(n6679), .A2(n599), .ZN(n4942) );
  AOI222_X1 U4446 ( .A1(vis_r10_o[6]), .A2(n617), .B1(vis_r11_o[6]), .B2(n4862), .C1(vis_r9_o[6]), .C2(n602), .ZN(n4943) );
  AOI221_X1 U4447 ( .B1(vis_r14_o[6]), .B2(n468), .C1(vis_r8_o[6]), .C2(n4856), 
        .A(n4945), .ZN(n4944) );
  NAND4_X1 U4448 ( .A1(n5273), .A2(n5188), .A3(n5189), .A4(n5190), .ZN(n5186)
         );
  NAND2_X1 U4449 ( .A1(n4864), .A2(n4940), .ZN(n5188) );
  AOI222_X1 U4450 ( .A1(vis_r10_o[7]), .A2(n617), .B1(vis_r11_o[7]), .B2(n4862), .C1(vis_r9_o[7]), .C2(n602), .ZN(n5189) );
  AOI221_X1 U4452 ( .B1(vis_r14_o[7]), .B2(n5272), .C1(vis_r8_o[7]), .C2(n4856), .A(n5191), .ZN(n5190) );
  NAND4_X1 U4453 ( .A1(n5277), .A2(n5546), .A3(n5547), .A4(n5548), .ZN(n5101)
         );
  NAND2_X1 U4454 ( .A1(n4864), .A2(n8082), .ZN(n5546) );
  AOI222_X1 U4455 ( .A1(vis_r10_o[5]), .A2(n617), .B1(vis_r11_o[5]), .B2(n615), 
        .C1(vis_r9_o[5]), .C2(n4863), .ZN(n5547) );
  AOI221_X1 U4456 ( .B1(vis_r14_o[5]), .B2(n5272), .C1(vis_r8_o[5]), .C2(n628), 
        .A(n5549), .ZN(n5548) );
  NOR2_X1 U4457 ( .A1(n7279), .A2(n4124), .ZN(Dqfhu6) );
  AOI211_X1 U4458 ( .C1(n1902), .C2(n3189), .A(n4125), .B(n2530), .ZN(n4124)
         );
  INV_X1 U4459 ( .A(n4127), .ZN(n2530) );
  OAI221_X1 U4460 ( .B1(n84), .B2(n4128), .C1(n524), .C2(n4129), .A(n4130), 
        .ZN(n4125) );
  NAND3_X1 U4461 ( .A1(n5420), .A2(n5421), .A3(n5422), .ZN(n3398) );
  OAI21_X1 U4462 ( .B1(n635), .B2(n5424), .A(n5425), .ZN(n5421) );
  AOI22_X1 U4463 ( .A1(n2551), .A2(n3297), .B1(Nxkbx6[31]), .B2(n438), .ZN(
        n5420) );
  AOI221_X1 U4464 ( .B1(vis_apsr_o[2]), .B2(n4342), .C1(n5423), .C2(n4253), 
        .A(Affpw6[30]), .ZN(n5422) );
  OAI211_X1 U4465 ( .C1(n4504), .C2(n5914), .A(n2370), .B(n5418), .ZN(n5415)
         );
  AOI22_X1 U4466 ( .A1(vis_psp_o[7]), .A2(n229), .B1(vis_r12_o[9]), .B2(n4290), 
        .ZN(n5418) );
  OAI211_X1 U4467 ( .C1(n4504), .C2(n5960), .A(n2360), .B(n4517), .ZN(n4514)
         );
  AOI22_X1 U4468 ( .A1(vis_psp_o[4]), .A2(n229), .B1(vis_r12_o[6]), .B2(n4290), 
        .ZN(n4517) );
  OAI22_X1 U4469 ( .A1(n2923), .A2(n476), .B1(n65), .B2(n2924), .ZN(n2922) );
  NAND2_X1 U4470 ( .A1(n7433), .A2(n4732), .ZN(n2924) );
  NOR3_X1 U4471 ( .A1(n2950), .A2(n7433), .A3(n1587), .ZN(n2923) );
  OAI21_X1 U4472 ( .B1(n5042), .B2(n4564), .A(n2951), .ZN(n2950) );
  AOI22_X1 U4473 ( .A1(n1724), .A2(n266), .B1(vis_apsr_o[1]), .B2(n4131), .ZN(
        n4129) );
  OAI21_X1 U4474 ( .B1(n7355), .B2(n522), .A(n4132), .ZN(n4131) );
  NAND3_X1 U4475 ( .A1(n7283), .A2(n538), .A3(n4133), .ZN(n4132) );
  AOI22_X1 U4476 ( .A1(n2940), .A2(n2941), .B1(n2610), .B2(vis_apsr_o[3]), 
        .ZN(n2939) );
  AND4_X1 U4477 ( .A1(n5282), .A2(n5765), .A3(n5766), .A4(n5767), .ZN(n3956)
         );
  NAND2_X1 U4478 ( .A1(n599), .A2(n8167), .ZN(n5765) );
  AOI222_X1 U4479 ( .A1(n617), .A2(vis_r10_o[4]), .B1(n4862), .B2(vis_r11_o[4]), .C1(n602), .C2(vis_r9_o[4]), .ZN(n5766) );
  AOI221_X1 U4480 ( .B1(n468), .B2(vis_r14_o[4]), .C1(n628), .C2(vis_r8_o[4]), 
        .A(n5768), .ZN(n5767) );
  NAND2_X1 U4482 ( .A1(n6465), .A2(n6466), .ZN(n5537) );
  AOI221_X1 U4483 ( .B1(vis_r2_o[9]), .B2(n561), .C1(vis_r0_o[9]), .C2(n547), 
        .A(n6468), .ZN(n6465) );
  AOI221_X1 U4484 ( .B1(vis_r3_o[9]), .B2(n567), .C1(vis_r7_o[9]), .C2(n565), 
        .A(n6467), .ZN(n6466) );
  OAI22_X1 U4485 ( .A1(n541), .A2(n6524), .B1(n540), .B2(n5428), .ZN(n6468) );
  NAND2_X1 U4486 ( .A1(n6520), .A2(n6521), .ZN(n5343) );
  AOI221_X1 U4487 ( .B1(n561), .B2(vis_r2_o[5]), .C1(n550), .C2(vis_r0_o[5]), 
        .A(n6525), .ZN(n6520) );
  AOI221_X1 U4488 ( .B1(n567), .B2(vis_r3_o[5]), .C1(n565), .C2(vis_r7_o[5]), 
        .A(n6522), .ZN(n6521) );
  OAI22_X1 U4489 ( .A1(n6487), .A2(n541), .B1(n5411), .B2(n540), .ZN(n6525) );
  NAND2_X1 U4490 ( .A1(n6499), .A2(n6500), .ZN(n5538) );
  AOI221_X1 U4491 ( .B1(n561), .B2(vis_r2_o[6]), .C1(n550), .C2(vis_r0_o[6]), 
        .A(n6502), .ZN(n6499) );
  AOI221_X1 U4492 ( .B1(n567), .B2(vis_r3_o[6]), .C1(n565), .C2(vis_r7_o[6]), 
        .A(n6501), .ZN(n6500) );
  OAI22_X1 U4493 ( .A1(n6394), .A2(n541), .B1(n5352), .B2(n540), .ZN(n6502) );
  NAND2_X1 U4494 ( .A1(n6494), .A2(n6495), .ZN(n5342) );
  AOI221_X1 U4495 ( .B1(n561), .B2(vis_r2_o[7]), .C1(n550), .C2(vis_r0_o[7]), 
        .A(n6497), .ZN(n6494) );
  AOI221_X1 U4496 ( .B1(n567), .B2(vis_r3_o[7]), .C1(n565), .C2(vis_r7_o[7]), 
        .A(n6496), .ZN(n6495) );
  OAI22_X1 U4497 ( .A1(n6571), .A2(n541), .B1(n5462), .B2(n540), .ZN(n6497) );
  NAND2_X1 U4498 ( .A1(n6505), .A2(n6506), .ZN(n5283) );
  AOI221_X1 U4499 ( .B1(n561), .B2(vis_r2_o[4]), .C1(n550), .C2(vis_r0_o[4]), 
        .A(n6508), .ZN(n6505) );
  AOI221_X1 U4500 ( .B1(n567), .B2(vis_r3_o[4]), .C1(n565), .C2(vis_r7_o[4]), 
        .A(n6507), .ZN(n6506) );
  OAI22_X1 U4501 ( .A1(n6586), .A2(n541), .B1(n5348), .B2(n540), .ZN(n6508) );
  NAND2_X1 U4502 ( .A1(n6008), .A2(n6009), .ZN(n5491) );
  AOI221_X1 U4503 ( .B1(n561), .B2(vis_r2_o[3]), .C1(n550), .C2(vis_r0_o[3]), 
        .A(n6011), .ZN(n6008) );
  AOI221_X1 U4504 ( .B1(n567), .B2(vis_r3_o[3]), .C1(n565), .C2(vis_r7_o[3]), 
        .A(n6010), .ZN(n6009) );
  OAI22_X1 U4505 ( .A1(n6570), .A2(n541), .B1(n5461), .B2(n540), .ZN(n6011) );
  AOI22_X1 U4506 ( .A1(n2947), .A2(n2941), .B1(n2610), .B2(n2948), .ZN(n2927)
         );
  XNOR2_X1 U4507 ( .A(vis_apsr_o[2]), .B(n93), .ZN(n2948) );
  XNOR2_X1 U4508 ( .A(n93), .B(n1543), .ZN(n2947) );
  OAI21_X1 U4509 ( .B1(n4795), .B2(n2510), .A(n1980), .ZN(n8014) );
  NAND3_X1 U4510 ( .A1(vis_pc_o[0]), .A2(n1981), .A3(n1430), .ZN(n1980) );
  AOI22_X1 U4511 ( .A1(n2887), .A2(n2888), .B1(n7279), .B2(n963), .ZN(Oxohu6)
         );
  NOR4_X1 U4512 ( .A1(n2889), .A2(n2890), .A3(n2891), .A4(n2892), .ZN(n2888)
         );
  NOR2_X1 U4513 ( .A1(n2900), .A2(n2125), .ZN(n2887) );
  AND4_X1 U4514 ( .A1(n476), .A2(n237), .A3(n2893), .A4(n2894), .ZN(n2891) );
  NAND2_X1 U4515 ( .A1(n6097), .A2(n6098), .ZN(n5945) );
  AOI221_X1 U4516 ( .B1(vis_r2_o[14]), .B2(n6003), .C1(vis_r0_o[14]), .C2(n547), .A(n6100), .ZN(n6097) );
  AOI221_X1 U4517 ( .B1(vis_r3_o[14]), .B2(n567), .C1(vis_r7_o[14]), .C2(n5999), .A(n6099), .ZN(n6098) );
  OAI22_X1 U4518 ( .A1(n6006), .A2(n6484), .B1(n6007), .B2(n5410), .ZN(n6100)
         );
  NAND2_X1 U4519 ( .A1(n6461), .A2(n6462), .ZN(n5943) );
  AOI221_X1 U4520 ( .B1(vis_r2_o[10]), .B2(n6003), .C1(vis_r0_o[10]), .C2(n547), .A(n6464), .ZN(n6461) );
  AOI221_X1 U4521 ( .B1(vis_r3_o[10]), .B2(n567), .C1(vis_r7_o[10]), .C2(n565), 
        .A(n6463), .ZN(n6462) );
  OAI22_X1 U4522 ( .A1(n541), .A2(n6574), .B1(n540), .B2(n5463), .ZN(n6464) );
  AND2_X1 U4523 ( .A1(n4933), .A2(n4934), .ZN(n2612) );
  AOI221_X1 U4524 ( .B1(vis_r6_o[9]), .B2(n4872), .C1(vis_r1_o[9]), .C2(n575), 
        .A(n4936), .ZN(n4933) );
  AOI221_X1 U4525 ( .B1(vis_r5_o[9]), .B2(n4867), .C1(vis_r4_o[9]), .C2(n581), 
        .A(n4935), .ZN(n4934) );
  OAI22_X1 U4526 ( .A1(n4875), .A2(n3341), .B1(n4876), .B2(n5523), .ZN(n4936)
         );
  AND2_X1 U4527 ( .A1(n4950), .A2(n4951), .ZN(n2628) );
  AOI221_X1 U4528 ( .B1(vis_r5_o[23]), .B2(n4867), .C1(vis_r4_o[23]), .C2(
        n4868), .A(n4952), .ZN(n4951) );
  AOI221_X1 U4529 ( .B1(vis_r6_o[23]), .B2(n4872), .C1(vis_r1_o[23]), .C2(
        n4873), .A(n4953), .ZN(n4950) );
  OAI22_X1 U4530 ( .A1(n4870), .A2(n7643), .B1(n4871), .B2(n6291), .ZN(n4952)
         );
  AND2_X1 U4531 ( .A1(n5705), .A2(n5706), .ZN(n2624) );
  AOI221_X1 U4532 ( .B1(vis_r6_o[27]), .B2(n576), .C1(vis_r1_o[27]), .C2(n4873), .A(n5708), .ZN(n5705) );
  AOI221_X1 U4533 ( .B1(vis_r5_o[27]), .B2(n582), .C1(vis_r4_o[27]), .C2(n4868), .A(n5707), .ZN(n5706) );
  OAI22_X1 U4534 ( .A1(n572), .A2(n7704), .B1(n4876), .B2(n5493), .ZN(n5708)
         );
  AND2_X1 U4535 ( .A1(n5377), .A2(n5378), .ZN(n2627) );
  AOI221_X1 U4537 ( .B1(vis_r6_o[24]), .B2(n4872), .C1(vis_r1_o[24]), .C2(
        n4873), .A(n5380), .ZN(n5377) );
  AOI221_X1 U4538 ( .B1(vis_r5_o[24]), .B2(n4867), .C1(vis_r4_o[24]), .C2(
        n4868), .A(n5379), .ZN(n5378) );
  OAI22_X1 U4539 ( .A1(n4875), .A2(n7818), .B1(n4876), .B2(n5470), .ZN(n5380)
         );
  AND2_X1 U4540 ( .A1(n4865), .A2(n4866), .ZN(n2640) );
  AOI221_X1 U4541 ( .B1(vis_r6_o[12]), .B2(n4872), .C1(vis_r1_o[12]), .C2(
        n4873), .A(n4874), .ZN(n4865) );
  AOI221_X1 U4542 ( .B1(vis_r5_o[12]), .B2(n4867), .C1(vis_r4_o[12]), .C2(
        n4868), .A(n4869), .ZN(n4866) );
  OAI22_X1 U4543 ( .A1(n4875), .A2(n4179), .B1(n4876), .B2(n5526), .ZN(n4874)
         );
  AND2_X1 U4544 ( .A1(n4924), .A2(n4925), .ZN(n2626) );
  AOI221_X1 U4545 ( .B1(vis_r5_o[25]), .B2(n4867), .C1(vis_r4_o[25]), .C2(
        n4868), .A(n4926), .ZN(n4925) );
  AOI221_X1 U4546 ( .B1(vis_r6_o[25]), .B2(n4872), .C1(vis_r1_o[25]), .C2(
        n4873), .A(n4927), .ZN(n4924) );
  OAI22_X1 U4547 ( .A1(n4870), .A2(n7571), .B1(n4871), .B2(n6313), .ZN(n4926)
         );
  AND2_X1 U4548 ( .A1(n5594), .A2(n5595), .ZN(n2641) );
  AOI221_X1 U4549 ( .B1(vis_r6_o[11]), .B2(n576), .C1(vis_r1_o[11]), .C2(n4873), .A(n5597), .ZN(n5594) );
  AOI221_X1 U4550 ( .B1(vis_r5_o[11]), .B2(n582), .C1(vis_r4_o[11]), .C2(n4868), .A(n5596), .ZN(n5595) );
  OAI22_X1 U4551 ( .A1(n572), .A2(n7790), .B1(n4876), .B2(n5606), .ZN(n5597)
         );
  AND2_X1 U4552 ( .A1(n5168), .A2(n5169), .ZN(n2629) );
  AOI221_X1 U4553 ( .B1(vis_r6_o[22]), .B2(n4872), .C1(vis_r1_o[22]), .C2(
        n4873), .A(n5171), .ZN(n5168) );
  AOI221_X1 U4554 ( .B1(vis_r5_o[22]), .B2(n4867), .C1(vis_r4_o[22]), .C2(
        n4868), .A(n5170), .ZN(n5169) );
  OAI22_X1 U4555 ( .A1(n4875), .A2(n7763), .B1(n4876), .B2(n5551), .ZN(n5171)
         );
  AND2_X1 U4556 ( .A1(n4962), .A2(n4963), .ZN(n2625) );
  AOI221_X1 U4557 ( .B1(vis_r6_o[26]), .B2(n4872), .C1(vis_r1_o[26]), .C2(
        n4873), .A(n4965), .ZN(n4962) );
  AOI221_X1 U4558 ( .B1(vis_r5_o[26]), .B2(n4867), .C1(vis_r4_o[26]), .C2(
        n4868), .A(n4964), .ZN(n4963) );
  OAI22_X1 U4559 ( .A1(n4875), .A2(n7784), .B1(n4876), .B2(n5556), .ZN(n4965)
         );
  AND2_X1 U4560 ( .A1(n5144), .A2(n5145), .ZN(n2638) );
  AOI221_X1 U4561 ( .B1(vis_r6_o[14]), .B2(n4872), .C1(vis_r1_o[14]), .C2(
        n4873), .A(n5147), .ZN(n5144) );
  AOI221_X1 U4562 ( .B1(vis_r5_o[14]), .B2(n4867), .C1(vis_r4_o[14]), .C2(
        n4868), .A(n5146), .ZN(n5145) );
  OAI22_X1 U4563 ( .A1(n4875), .A2(n7806), .B1(n4876), .B2(n5507), .ZN(n5147)
         );
  AND2_X1 U4564 ( .A1(n5058), .A2(n5059), .ZN(n2613) );
  AOI221_X1 U4565 ( .B1(vis_r6_o[8]), .B2(n4872), .C1(vis_r1_o[8]), .C2(n575), 
        .A(n5061), .ZN(n5058) );
  AOI221_X1 U4566 ( .B1(vis_r5_o[8]), .B2(n4867), .C1(vis_r4_o[8]), .C2(n581), 
        .A(n5060), .ZN(n5059) );
  OAI22_X1 U4567 ( .A1(n4875), .A2(n7787), .B1(n569), .B2(n5598), .ZN(n5061)
         );
  AND2_X1 U4568 ( .A1(n5362), .A2(n5363), .ZN(n2639) );
  AOI221_X1 U4569 ( .B1(vis_r6_o[13]), .B2(n4872), .C1(vis_r1_o[13]), .C2(
        n4873), .A(n5365), .ZN(n5362) );
  AOI221_X1 U4570 ( .B1(vis_r5_o[13]), .B2(n4867), .C1(vis_r4_o[13]), .C2(
        n4868), .A(n5364), .ZN(n5363) );
  OAI22_X1 U4571 ( .A1(n4875), .A2(n7778), .B1(n4876), .B2(n5584), .ZN(n5365)
         );
  AND2_X1 U4572 ( .A1(n4902), .A2(n4903), .ZN(n2637) );
  AOI221_X1 U4573 ( .B1(vis_r6_o[15]), .B2(n4872), .C1(vis_r1_o[15]), .C2(
        n4873), .A(n4905), .ZN(n4902) );
  AOI221_X1 U4574 ( .B1(vis_r5_o[15]), .B2(n4867), .C1(vis_r4_o[15]), .C2(
        n4868), .A(n4904), .ZN(n4903) );
  OAI22_X1 U4575 ( .A1(n4875), .A2(n7766), .B1(n4876), .B2(n5552), .ZN(n4905)
         );
  AND2_X1 U4576 ( .A1(n4970), .A2(n4971), .ZN(n2642) );
  AOI221_X1 U4577 ( .B1(vis_r6_o[10]), .B2(n4872), .C1(vis_r1_o[10]), .C2(
        n4873), .A(n4973), .ZN(n4970) );
  AOI221_X1 U4578 ( .B1(vis_r5_o[10]), .B2(n4867), .C1(vis_r4_o[10]), .C2(n581), .A(n4972), .ZN(n4971) );
  OAI22_X1 U4579 ( .A1(n4875), .A2(n7757), .B1(n4876), .B2(n5534), .ZN(n4973)
         );
  AND2_X1 U4580 ( .A1(n4883), .A2(n4884), .ZN(n2622) );
  AOI221_X1 U4581 ( .B1(vis_r5_o[29]), .B2(n4867), .C1(vis_r4_o[29]), .C2(
        n4868), .A(n4885), .ZN(n4884) );
  AOI221_X1 U4582 ( .B1(vis_r6_o[29]), .B2(n4872), .C1(vis_r1_o[29]), .C2(
        n4873), .A(n4886), .ZN(n4883) );
  OAI22_X1 U4583 ( .A1(n4870), .A2(n7341), .B1(n4871), .B2(n6289), .ZN(n4885)
         );
  AND2_X1 U4584 ( .A1(n4894), .A2(n4895), .ZN(n2619) );
  AOI221_X1 U4585 ( .B1(vis_r5_o[31]), .B2(n4867), .C1(vis_r4_o[31]), .C2(
        n4868), .A(n4896), .ZN(n4895) );
  AOI221_X1 U4586 ( .B1(vis_r6_o[31]), .B2(n4872), .C1(vis_r1_o[31]), .C2(
        n4873), .A(n4897), .ZN(n4894) );
  OAI22_X1 U4587 ( .A1(n4870), .A2(n7512), .B1(n4871), .B2(n2815), .ZN(n4896)
         );
  AND2_X1 U4588 ( .A1(n5121), .A2(n5122), .ZN(n2623) );
  AOI221_X1 U4589 ( .B1(vis_r6_o[28]), .B2(n4872), .C1(vis_r1_o[28]), .C2(
        n4873), .A(n5124), .ZN(n5121) );
  AOI221_X1 U4591 ( .B1(vis_r5_o[28]), .B2(n4867), .C1(vis_r4_o[28]), .C2(
        n4868), .A(n5123), .ZN(n5122) );
  OAI22_X1 U4592 ( .A1(n4875), .A2(n8268), .B1(n4876), .B2(n8274), .ZN(n5124)
         );
  AND2_X1 U4593 ( .A1(n5438), .A2(n5439), .ZN(n2620) );
  AOI221_X1 U4594 ( .B1(vis_r6_o[30]), .B2(n576), .C1(vis_r1_o[30]), .C2(n4873), .A(n5441), .ZN(n5438) );
  AOI221_X1 U4595 ( .B1(vis_r5_o[30]), .B2(n582), .C1(vis_r4_o[30]), .C2(n4868), .A(n5440), .ZN(n5439) );
  OAI22_X1 U4596 ( .A1(n572), .A2(n7793), .B1(n4876), .B2(n5541), .ZN(n5441)
         );
  NAND3_X1 U4597 ( .A1(n2562), .A2(n4512), .A3(n1540), .ZN(n5246) );
  OAI211_X1 U4598 ( .C1(n5248), .C2(n5249), .A(n82), .B(n517), .ZN(n5247) );
  NOR2_X1 U4599 ( .A1(n5231), .A2(n3721), .ZN(n5245) );
  AOI221_X1 U4600 ( .B1(n4166), .B2(n2262), .C1(n2730), .C2(n4168), .A(n4169), 
        .ZN(n4165) );
  OAI21_X1 U4601 ( .B1(n2757), .B2(n4171), .A(n2597), .ZN(n4169) );
  NAND2_X1 U4602 ( .A1(n6601), .A2(n7433), .ZN(n4171) );
  OAI211_X2 U4603 ( .C1(n7525), .C2(n7526), .A(n5644), .B(n5645), .ZN(n56) );
  AOI22_X1 U4604 ( .A1(n1706), .A2(n5070), .B1(n3551), .B2(n4506), .ZN(n5644)
         );
  AOI211_X1 U4605 ( .C1(n3099), .C2(n4637), .A(n5646), .B(n5647), .ZN(n5645)
         );
  AOI21_X1 U4606 ( .B1(n7525), .B2(n7526), .A(n7524), .ZN(n5647) );
  AOI221_X1 U4607 ( .B1(n4166), .B2(n475), .C1(n2730), .C2(n4941), .A(n5158), 
        .ZN(n5157) );
  OAI21_X1 U4608 ( .B1(n2757), .B2(n5159), .A(n2597), .ZN(n5158) );
  NAND2_X1 U4609 ( .A1(n6601), .A2(n270), .ZN(n5159) );
  OAI22_X1 U4610 ( .A1(n659), .A2(n3484), .B1(n5381), .B2(n5382), .ZN(n3806)
         );
  OAI211_X1 U4611 ( .C1(n4176), .C2(n3482), .A(n2419), .B(n5383), .ZN(n5382)
         );
  OAI221_X1 U4612 ( .B1(n640), .B2(n3596), .C1(n2468), .C2(n6234), .A(n5384), 
        .ZN(n5381) );
  AOI222_X1 U4613 ( .A1(vis_r8_o[24]), .A2(n2336), .B1(vis_msp_o[22]), .B2(
        n2474), .C1(vis_r9_o[24]), .C2(n2338), .ZN(n5383) );
  NAND3_X1 U4614 ( .A1(n7661), .A2(n7664), .A3(n7657), .ZN(n137) );
  NAND3_X1 U4615 ( .A1(n7450), .A2(n7655), .A3(n7429), .ZN(n138) );
  NAND4_X1 U4616 ( .A1(n7681), .A2(n7693), .A3(n7667), .A4(n151), .ZN(n136) );
  OAI222_X1 U4617 ( .A1(n3811), .A2(n3900), .B1(n4284), .B2(n242), .C1(n1809), 
        .C2(n661), .ZN(n443) );
  XNOR2_X1 U4618 ( .A(vis_pc_o[0]), .B(n1430), .ZN(n4284) );
  OAI211_X1 U4619 ( .C1(n6353), .C2(n6354), .A(n8106), .B(n8145), .ZN(n6125)
         );
  OR2_X1 U4620 ( .A1(n7586), .A2(n7574), .ZN(n6354) );
  AOI22_X1 U4621 ( .A1(n6356), .A2(n6702), .B1(n7622), .B2(n8230), .ZN(n6353)
         );
  OAI211_X1 U4622 ( .C1(n6339), .C2(n6322), .A(n8170), .B(n8169), .ZN(n6321)
         );
  AOI22_X1 U4623 ( .A1(n6340), .A2(n7613), .B1(n7614), .B2(n4433), .ZN(n6339)
         );
  AOI21_X1 U4624 ( .B1(n7612), .B2(n4434), .A(n7677), .ZN(n6340) );
  NOR3_X1 U4625 ( .A1(vis_ipsr_o[4]), .A2(vis_ipsr_o[5]), .A3(n5088), .ZN(
        n5862) );
  OAI21_X1 U4626 ( .B1(n6211), .B2(n6243), .A(n6244), .ZN(n6141) );
  OAI21_X1 U4627 ( .B1(n7601), .B2(n7280), .A(n6245), .ZN(n6244) );
  AOI22_X1 U4628 ( .A1(n6246), .A2(n6204), .B1(n6247), .B2(n2799), .ZN(n6243)
         );
  AOI21_X1 U4629 ( .B1(n3033), .B2(n6248), .A(n6201), .ZN(n6246) );
  OAI21_X1 U4630 ( .B1(n6345), .B2(n6346), .A(n6347), .ZN(n5321) );
  OAI21_X1 U4631 ( .B1(n7586), .B2(n7574), .A(n6125), .ZN(n6347) );
  AOI22_X1 U4632 ( .A1(n6348), .A2(n6326), .B1(n4460), .B2(n3063), .ZN(n6346)
         );
  INV_X1 U4633 ( .A(n6327), .ZN(n4460) );
  OAI22_X1 U4634 ( .A1(n659), .A2(n8204), .B1(n4812), .B2(n4813), .ZN(n3801)
         );
  OAI211_X1 U4635 ( .C1(n4176), .C2(n8120), .A(n2456), .B(n4814), .ZN(n4813)
         );
  OAI221_X1 U4636 ( .B1(n640), .B2(n3587), .C1(n2468), .C2(n6178), .A(n4815), 
        .ZN(n4812) );
  AOI222_X1 U4637 ( .A1(vis_r8_o[29]), .A2(n2336), .B1(vis_msp_o[27]), .B2(
        n2474), .C1(vis_r9_o[29]), .C2(n2338), .ZN(n4814) );
  OAI22_X1 U4638 ( .A1(n659), .A2(n8196), .B1(n5160), .B2(n5161), .ZN(n3808)
         );
  OAI211_X1 U4639 ( .C1(n4176), .C2(n8114), .A(n2437), .B(n5162), .ZN(n5161)
         );
  OAI221_X1 U4640 ( .B1(n640), .B2(n3581), .C1(n2468), .C2(n6271), .A(n5163), 
        .ZN(n5160) );
  AOI222_X1 U4641 ( .A1(vis_r8_o[22]), .A2(n2336), .B1(vis_msp_o[20]), .B2(
        n2474), .C1(vis_r9_o[22]), .C2(n2338), .ZN(n5162) );
  OAI22_X1 U4642 ( .A1(n659), .A2(n3672), .B1(n4604), .B2(n4605), .ZN(n3809)
         );
  OAI211_X1 U4643 ( .C1(n4176), .C2(n8130), .A(n2438), .B(n4606), .ZN(n4605)
         );
  OAI221_X1 U4644 ( .B1(n640), .B2(n3650), .C1(n2468), .C2(n6220), .A(n4607), 
        .ZN(n4604) );
  AOI222_X1 U4645 ( .A1(vis_r8_o[21]), .A2(n2336), .B1(vis_msp_o[19]), .B2(
        n2474), .C1(vis_r9_o[21]), .C2(n2338), .ZN(n4606) );
  OAI22_X1 U4646 ( .A1(n659), .A2(n8223), .B1(n4661), .B2(n4662), .ZN(n3810)
         );
  OAI211_X1 U4647 ( .C1(n4176), .C2(n8214), .A(n2440), .B(n4663), .ZN(n4662)
         );
  OAI221_X1 U4648 ( .B1(n640), .B2(n8211), .C1(n2468), .C2(n8208), .A(n4665), 
        .ZN(n4661) );
  AOI222_X1 U4649 ( .A1(vis_r8_o[20]), .A2(n2336), .B1(vis_msp_o[18]), .B2(
        n2474), .C1(vis_r9_o[20]), .C2(n2338), .ZN(n4663) );
  OAI21_X1 U4650 ( .B1(n6388), .B2(n6389), .A(n6390), .ZN(n6132) );
  OAI21_X1 U4651 ( .B1(n7572), .B2(n3645), .A(n6131), .ZN(n6390) );
  AOI22_X1 U4652 ( .A1(n6391), .A2(n6368), .B1(n6392), .B2(n4282), .ZN(n6389)
         );
  AOI21_X1 U4653 ( .B1(n3640), .B2(n6393), .A(n6367), .ZN(n6391) );
  OAI211_X1 U4654 ( .C1(n6254), .C2(n6255), .A(n2811), .B(n8135), .ZN(n6139)
         );
  NAND2_X1 U4655 ( .A1(n8150), .A2(n5192), .ZN(n6255) );
  AOI22_X1 U4656 ( .A1(n6256), .A2(n6776), .B1(n7620), .B2(n4468), .ZN(n6254)
         );
  OAI211_X1 U4657 ( .C1(n6235), .C2(n6236), .A(n3121), .B(n8137), .ZN(n6233)
         );
  OR2_X1 U4658 ( .A1(n7595), .A2(n7581), .ZN(n6236) );
  AOI22_X1 U4659 ( .A1(n6237), .A2(n7605), .B1(n7606), .B2(n8233), .ZN(n6235)
         );
  AOI21_X1 U4660 ( .B1(n6711), .B2(n8246), .A(n6778), .ZN(n6237) );
  NOR4_X1 U4661 ( .A1(n5828), .A2(n3940), .A3(n5830), .A4(n5831), .ZN(n5827)
         );
  OAI221_X1 U4663 ( .B1(n6759), .B2(n2824), .C1(n7675), .C2(n2526), .A(n3947), 
        .ZN(n5830) );
  OAI221_X1 U4664 ( .B1(n7637), .B2(n3958), .C1(n7552), .C2(n3612), .A(n3931), 
        .ZN(n5828) );
  OAI221_X1 U4665 ( .B1(n6776), .B2(n2800), .C1(n6775), .C2(n3449), .A(n3979), 
        .ZN(n5831) );
  OAI22_X1 U4666 ( .A1(n659), .A2(n8195), .B1(n4174), .B2(n4175), .ZN(n3807)
         );
  OAI211_X1 U4667 ( .C1(n646), .C2(n8131), .A(n2442), .B(n4177), .ZN(n4175) );
  OAI221_X1 U4668 ( .B1(n640), .B2(n3781), .C1(n2468), .C2(n6207), .A(n4183), 
        .ZN(n4174) );
  AOI222_X1 U4669 ( .A1(vis_r8_o[23]), .A2(n2336), .B1(vis_msp_o[21]), .B2(
        n2474), .C1(vis_r9_o[23]), .C2(n2338), .ZN(n4177) );
  NAND2_X1 U4670 ( .A1(n5852), .A2(n5853), .ZN(n5261) );
  NOR4_X1 U4671 ( .A1(n5881), .A2(n5882), .A3(n5883), .A4(n5884), .ZN(n5852)
         );
  NOR4_X1 U4672 ( .A1(n5854), .A2(n5855), .A3(n5856), .A4(n5857), .ZN(n5853)
         );
  OAI221_X1 U4673 ( .B1(n7619), .B2(n2685), .C1(n7620), .C2(n2800), .A(n5893), 
        .ZN(n5882) );
  AOI22_X1 U4674 ( .A1(n6126), .A2(n7624), .B1(n6777), .B2(n4465), .ZN(n6327)
         );
  NAND2_X1 U4675 ( .A1(n6601), .A2(n2806), .ZN(n1706) );
  AOI22_X1 U4676 ( .A1(n7331), .A2(n2224), .B1(n5456), .B2(n6160), .ZN(n5902)
         );
  AOI221_X1 U4677 ( .B1(n5345), .B2(n2161), .C1(n2858), .C2(n3785), .A(n5795), 
        .ZN(n5792) );
  OAI22_X1 U4678 ( .A1(n7563), .A2(n2197), .B1(n7612), .B2(n2195), .ZN(n5795)
         );
  INV_X1 U4679 ( .A(n2065), .ZN(n2161) );
  NOR4_X1 U4680 ( .A1(n7378), .A2(n3623), .A3(n3831), .A4(n4232), .ZN(n5248)
         );
  AOI22_X1 U4681 ( .A1(n6139), .A2(n6776), .B1(n2809), .B2(n7673), .ZN(n6201)
         );
  AOI221_X1 U4682 ( .B1(vis_r14_o[23]), .B2(n2473), .C1(vis_r10_o[23]), .C2(
        n2322), .A(n650), .ZN(n4183) );
  AOI221_X1 U4683 ( .B1(vis_r14_o[24]), .B2(n2473), .C1(vis_r10_o[24]), .C2(
        n2322), .A(n650), .ZN(n5384) );
  AOI221_X1 U4684 ( .B1(vis_r14_o[22]), .B2(n2473), .C1(vis_r10_o[22]), .C2(
        n2322), .A(n650), .ZN(n5163) );
  AOI221_X1 U4685 ( .B1(vis_r14_o[28]), .B2(n2473), .C1(vis_r10_o[28]), .C2(
        n2322), .A(n650), .ZN(n5116) );
  AOI221_X1 U4686 ( .B1(vis_r14_o[21]), .B2(n2473), .C1(vis_r10_o[21]), .C2(
        n2322), .A(n654), .ZN(n4607) );
  AOI221_X1 U4687 ( .B1(vis_r14_o[20]), .B2(n2473), .C1(vis_r10_o[20]), .C2(
        n2322), .A(n654), .ZN(n4665) );
  AOI221_X1 U4688 ( .B1(vis_r14_o[29]), .B2(n2473), .C1(vis_r10_o[29]), .C2(
        n2322), .A(n654), .ZN(n4815) );
  AOI221_X1 U4689 ( .B1(vis_r14_o[30]), .B2(n2473), .C1(vis_r10_o[30]), .C2(
        n2322), .A(n650), .ZN(n5432) );
  AOI221_X1 U4690 ( .B1(vis_r14_o[31]), .B2(n2473), .C1(vis_r10_o[31]), .C2(
        n2322), .A(n654), .ZN(n4340) );
  NAND2_X1 U4691 ( .A1(n6056), .A2(n6057), .ZN(n5986) );
  AOI221_X1 U4692 ( .B1(vis_r2_o[22]), .B2(n6003), .C1(vis_r0_o[22]), .C2(n547), .A(n6059), .ZN(n6056) );
  AOI221_X1 U4693 ( .B1(vis_r3_o[22]), .B2(n567), .C1(vis_r7_o[22]), .C2(n5999), .A(n6058), .ZN(n6057) );
  OAI22_X1 U4694 ( .A1(n6006), .A2(n6583), .B1(n6007), .B2(n2727), .ZN(n6059)
         );
  NAND2_X1 U4695 ( .A1(n6052), .A2(n6053), .ZN(n5445) );
  AOI221_X1 U4696 ( .B1(vis_r2_o[21]), .B2(n6003), .C1(vis_r0_o[21]), .C2(n547), .A(n6055), .ZN(n6052) );
  AOI221_X1 U4698 ( .B1(vis_r3_o[21]), .B2(n567), .C1(vis_r7_o[21]), .C2(n5999), .A(n6054), .ZN(n6053) );
  OAI22_X1 U4699 ( .A1(n6006), .A2(n6480), .B1(n6007), .B2(n5409), .ZN(n6055)
         );
  NAND3_X1 U4700 ( .A1(n8146), .A2(n5197), .A3(n6396), .ZN(n6131) );
  OR3_X1 U4701 ( .A1(n6397), .A2(n7572), .A3(n3645), .ZN(n6396) );
  AOI21_X1 U4702 ( .B1(n8228), .B2(n7556), .A(n6398), .ZN(n6397) );
  AOI211_X1 U4703 ( .C1(n8241), .C2(n7323), .A(n7639), .B(n8256), .ZN(n6398)
         );
  OAI211_X1 U4704 ( .C1(n6342), .C2(n6343), .A(n4010), .B(n8138), .ZN(n6338)
         );
  NAND2_X1 U4705 ( .A1(n8153), .A2(n3930), .ZN(n6343) );
  AOI22_X1 U4706 ( .A1(n6344), .A2(n6701), .B1(n7611), .B2(n8229), .ZN(n6342)
         );
  AOI21_X1 U4707 ( .B1(n7610), .B2(n8243), .A(n7638), .ZN(n6344) );
  NAND4_X1 U4708 ( .A1(n2629), .A2(n5164), .A3(n5165), .A4(n5166), .ZN(n4941)
         );
  NAND2_X1 U4709 ( .A1(n4864), .A2(n8196), .ZN(n5164) );
  AOI222_X1 U4710 ( .A1(vis_r10_o[22]), .A2(n617), .B1(vis_r11_o[22]), .B2(
        n615), .C1(vis_r9_o[22]), .C2(n4863), .ZN(n5165) );
  AOI221_X1 U4711 ( .B1(vis_r14_o[22]), .B2(n5272), .C1(vis_r8_o[22]), .C2(
        n4856), .A(n5167), .ZN(n5166) );
  NAND4_X1 U4712 ( .A1(n2634), .A2(n4911), .A3(n4912), .A4(n4913), .ZN(n4425)
         );
  NAND2_X1 U4713 ( .A1(n599), .A2(n8177), .ZN(n4911) );
  AOI222_X1 U4714 ( .A1(vis_r10_o[18]), .A2(n617), .B1(vis_r11_o[18]), .B2(
        n4862), .C1(vis_r9_o[18]), .C2(n602), .ZN(n4912) );
  AOI221_X1 U4715 ( .B1(vis_r14_o[18]), .B2(n5272), .C1(vis_r8_o[18]), .C2(
        n628), .A(n4914), .ZN(n4913) );
  NAND4_X1 U4716 ( .A1(n2633), .A2(n5614), .A3(n5615), .A4(n5616), .ZN(n4988)
         );
  NAND2_X1 U4717 ( .A1(n4864), .A2(n8224), .ZN(n5614) );
  AOI222_X1 U4718 ( .A1(vis_r10_o[19]), .A2(n4861), .B1(vis_r11_o[19]), .B2(
        n615), .C1(vis_r9_o[19]), .C2(n4863), .ZN(n5615) );
  AOI221_X1 U4719 ( .B1(vis_r14_o[19]), .B2(n5272), .C1(vis_r8_o[19]), .C2(
        n4856), .A(n5617), .ZN(n5616) );
  NAND4_X1 U4720 ( .A1(n2630), .A2(n5003), .A3(n5004), .A4(n5005), .ZN(n4603)
         );
  NAND2_X1 U4721 ( .A1(n4864), .A2(n3672), .ZN(n5003) );
  AOI222_X1 U4722 ( .A1(vis_r10_o[21]), .A2(n617), .B1(vis_r11_o[21]), .B2(
        n4862), .C1(vis_r9_o[21]), .C2(n602), .ZN(n5004) );
  AOI221_X1 U4723 ( .B1(vis_r14_o[21]), .B2(n468), .C1(vis_r8_o[21]), .C2(
        n4856), .A(n5006), .ZN(n5005) );
  NAND4_X1 U4724 ( .A1(n2631), .A2(n4994), .A3(n4995), .A4(n4996), .ZN(n4666)
         );
  NAND2_X1 U4725 ( .A1(n4864), .A2(n8223), .ZN(n4994) );
  AOI222_X1 U4726 ( .A1(vis_r10_o[20]), .A2(n617), .B1(vis_r11_o[20]), .B2(
        n4862), .C1(vis_r9_o[20]), .C2(n602), .ZN(n4995) );
  AOI221_X1 U4727 ( .B1(vis_r14_o[20]), .B2(n468), .C1(vis_r8_o[20]), .C2(
        n4856), .A(n4997), .ZN(n4996) );
  NAND4_X1 U4728 ( .A1(n2636), .A2(n5079), .A3(n5080), .A4(n5081), .ZN(n4909)
         );
  NAND2_X1 U4729 ( .A1(n4864), .A2(n4185), .ZN(n5079) );
  AOI222_X1 U4730 ( .A1(vis_r10_o[16]), .A2(n617), .B1(vis_r11_o[16]), .B2(
        n4862), .C1(vis_r9_o[16]), .C2(n602), .ZN(n5080) );
  AOI221_X1 U4731 ( .B1(vis_r14_o[16]), .B2(n468), .C1(vis_r8_o[16]), .C2(
        n4856), .A(n5082), .ZN(n5081) );
  AOI21_X1 U4732 ( .B1(n5796), .B2(n2171), .A(n2170), .ZN(n2065) );
  OAI22_X1 U4733 ( .A1(n5903), .A2(vis_primask_o), .B1(n2386), .B2(n2590), 
        .ZN(n5796) );
  NAND4_X1 U4734 ( .A1(n2627), .A2(n5373), .A3(n5374), .A4(n5375), .ZN(n4956)
         );
  NAND2_X1 U4735 ( .A1(n4864), .A2(n3484), .ZN(n5373) );
  AOI222_X1 U4736 ( .A1(vis_r10_o[24]), .A2(n617), .B1(vis_r11_o[24]), .B2(
        n615), .C1(vis_r9_o[24]), .C2(n4863), .ZN(n5374) );
  AOI221_X1 U4737 ( .B1(vis_r14_o[24]), .B2(n5272), .C1(vis_r8_o[24]), .C2(
        n4856), .A(n5376), .ZN(n5375) );
  NAND4_X1 U4738 ( .A1(n2626), .A2(n4920), .A3(n4921), .A4(n4922), .ZN(n4496)
         );
  NAND2_X1 U4739 ( .A1(n6680), .A2(n599), .ZN(n4920) );
  AOI222_X1 U4740 ( .A1(vis_r10_o[25]), .A2(n617), .B1(vis_r11_o[25]), .B2(
        n4862), .C1(vis_r9_o[25]), .C2(n602), .ZN(n4921) );
  AOI221_X1 U4741 ( .B1(vis_r14_o[25]), .B2(n5272), .C1(vis_r8_o[25]), .C2(
        n628), .A(n4923), .ZN(n4922) );
  NAND4_X1 U4742 ( .A1(n2625), .A2(n4958), .A3(n4959), .A4(n4960), .ZN(n4678)
         );
  NAND2_X1 U4743 ( .A1(n599), .A2(n8283), .ZN(n4958) );
  AOI222_X1 U4744 ( .A1(vis_r10_o[26]), .A2(n617), .B1(vis_r11_o[26]), .B2(
        n4862), .C1(vis_r9_o[26]), .C2(n602), .ZN(n4959) );
  AOI221_X1 U4745 ( .B1(vis_r14_o[26]), .B2(n468), .C1(vis_r8_o[26]), .C2(
        n4856), .A(n4961), .ZN(n4960) );
  AOI22_X1 U4746 ( .A1(n6338), .A2(n6701), .B1(n3928), .B2(n7638), .ZN(n6312)
         );
  OAI222_X1 U4747 ( .A1(n7613), .A2(n3579), .B1(n7638), .B2(n4039), .C1(n7623), 
        .C2(n4472), .ZN(n5841) );
  NAND3_X1 U4748 ( .A1(n5862), .A2(vis_ipsr_o[2]), .A3(n5798), .ZN(n1796) );
  NAND3_X1 U4749 ( .A1(n5255), .A2(vis_ipsr_o[2]), .A3(n5862), .ZN(n1781) );
  OAI22_X1 U4750 ( .A1(n7257), .A2(n5456), .B1(n2224), .B2(n6157), .ZN(n5821)
         );
  OAI22_X1 U4751 ( .A1(n7620), .A2(n2809), .B1(n7619), .B2(n6139), .ZN(n6248)
         );
  OAI22_X1 U4752 ( .A1(n7649), .A2(n659), .B1(n650), .B2(n5696), .ZN(n5695) );
  NOR3_X1 U4753 ( .A1(n5697), .A2(n5698), .A3(n5699), .ZN(n5696) );
  OAI22_X1 U4754 ( .A1(n4288), .A2(n8092), .B1(n4291), .B2(n8058), .ZN(n5699)
         );
  OAI222_X1 U4755 ( .A1(n4502), .A2(n5873), .B1(n4503), .B2(n6148), .C1(n646), 
        .C2(n8107), .ZN(n5698) );
  OAI22_X1 U4756 ( .A1(n7654), .A2(n659), .B1(n650), .B2(n4680), .ZN(n4679) );
  NOR3_X1 U4757 ( .A1(n4681), .A2(n4682), .A3(n4683), .ZN(n4680) );
  OAI22_X1 U4758 ( .A1(n4288), .A2(n8282), .B1(n4291), .B2(n8071), .ZN(n4683)
         );
  OAI222_X1 U4759 ( .A1(n4502), .A2(n5895), .B1(n4503), .B2(n6080), .C1(n646), 
        .C2(n8123), .ZN(n4682) );
  NOR2_X1 U4760 ( .A1(n2757), .A2(n6601), .ZN(n4166) );
  OAI22_X1 U4761 ( .A1(n7614), .A2(n4432), .B1(n7612), .B2(n6321), .ZN(n6335)
         );
  OAI221_X1 U4762 ( .B1(HADDR[4]), .B2(n1537), .C1(n7534), .C2(N701), .A(n128), 
        .ZN(n7734) );
  OAI22_X1 U4763 ( .A1(n7611), .A2(n3928), .B1(n7610), .B2(n6338), .ZN(n6337)
         );
  AOI22_X1 U4764 ( .A1(n6125), .A2(n6702), .B1(n3064), .B2(n7637), .ZN(n6326)
         );
  AOI22_X1 U4765 ( .A1(n6321), .A2(n7613), .B1(n4432), .B2(n7677), .ZN(n6309)
         );
  AOI22_X1 U4766 ( .A1(n6131), .A2(n7556), .B1(n7323), .B2(n3643), .ZN(n6392)
         );
  AOI22_X1 U4767 ( .A1(n6245), .A2(n7618), .B1(n6710), .B2(n3036), .ZN(n6247)
         );
  AOI22_X1 U4768 ( .A1(n4437), .A2(n7609), .B1(n7607), .B2(n6216), .ZN(n6231)
         );
  AOI22_X1 U4769 ( .A1(n6135), .A2(n7553), .B1(n7551), .B2(n3668), .ZN(n6263)
         );
  AOI22_X1 U4770 ( .A1(n4437), .A2(n7608), .B1(n6216), .B2(n7674), .ZN(n6222)
         );
  OAI221_X1 U4771 ( .B1(n7567), .B2(n4276), .C1(n7331), .C2(n1781), .A(n5885), 
        .ZN(n5884) );
  AOI22_X1 U4772 ( .A1(n3989), .A2(n8243), .B1(n3938), .B2(n3785), .ZN(n5885)
         );
  INV_X1 U4773 ( .A(n1796), .ZN(n3938) );
  OAI221_X1 U4774 ( .B1(n6711), .B2(n3778), .C1(n6710), .C2(n3449), .A(n5858), 
        .ZN(n5857) );
  AOI22_X1 U4775 ( .A1(n3967), .A2(n4454), .B1(n3951), .B2(n8159), .ZN(n5858)
         );
  INV_X1 U4776 ( .A(n1636), .ZN(n3967) );
  OAI221_X1 U4777 ( .B1(n7556), .B2(n3862), .C1(n7323), .C2(n4843), .A(n5890), 
        .ZN(n5883) );
  AOI22_X1 U4778 ( .A1(n3973), .A2(n8236), .B1(n3935), .B2(n4487), .ZN(n5890)
         );
  OAI221_X1 U4780 ( .B1(n7551), .B2(n3677), .C1(n7624), .C2(n4472), .A(n3948), 
        .ZN(n5856) );
  INV_X1 U4781 ( .A(n5866), .ZN(n3948) );
  OAI222_X1 U4782 ( .A1(n2472), .A2(n7562), .B1(n2426), .B2(n7607), .C1(n4121), 
        .C2(n7609), .ZN(n5866) );
  OAI221_X1 U4783 ( .B1(n7554), .B2(n2526), .C1(n7555), .C2(n2824), .A(n5871), 
        .ZN(n5855) );
  AOI22_X1 U4784 ( .A1(n3977), .A2(n8231), .B1(n3946), .B2(n4474), .ZN(n5871)
         );
  OAI221_X1 U4785 ( .B1(n7558), .B2(n3624), .C1(n7564), .C2(n2357), .A(n5874), 
        .ZN(n5854) );
  AOI222_X1 U4786 ( .A1(n3939), .A2(n4433), .B1(n3975), .B2(n8229), .C1(n3959), 
        .C2(n4434), .ZN(n5874) );
  OAI221_X1 U4787 ( .B1(n7606), .B2(n5838), .C1(n7618), .C2(n3558), .A(n5896), 
        .ZN(n5881) );
  AOI222_X1 U4788 ( .A1(n3985), .A2(n8242), .B1(n3954), .B2(n4482), .C1(n3971), 
        .C2(n8230), .ZN(n5896) );
  OAI221_X1 U4789 ( .B1(n4276), .B2(n7568), .C1(n1781), .C2(n7257), .A(n3937), 
        .ZN(n5845) );
  INV_X1 U4790 ( .A(n5847), .ZN(n3937) );
  OAI222_X1 U4791 ( .A1(n6701), .A2(n3199), .B1(n7670), .B2(n3542), .C1(n7679), 
        .C2(n1796), .ZN(n5847) );
  OAI22_X1 U4792 ( .A1(n659), .A2(n8261), .B1(n5113), .B2(n5114), .ZN(n3802)
         );
  OAI211_X1 U4793 ( .C1(n4176), .C2(n8269), .A(n2457), .B(n5115), .ZN(n5114)
         );
  OAI221_X1 U4794 ( .B1(n640), .B2(n8266), .C1(n2468), .C2(n8263), .A(n5116), 
        .ZN(n5113) );
  AOI222_X1 U4795 ( .A1(vis_r8_o[28]), .A2(n2336), .B1(vis_msp_o[26]), .B2(
        n2474), .C1(vis_r9_o[28]), .C2(n2338), .ZN(n5115) );
  OAI22_X1 U4796 ( .A1(n659), .A2(n2779), .B1(n5429), .B2(n5430), .ZN(n3798)
         );
  OAI211_X1 U4797 ( .C1(n646), .C2(n8108), .A(n2451), .B(n5431), .ZN(n5430) );
  OAI221_X1 U4798 ( .B1(n640), .B2(n3601), .C1(n2468), .C2(n6221), .A(n5432), 
        .ZN(n5429) );
  AOI222_X1 U4799 ( .A1(vis_r8_o[30]), .A2(n2336), .B1(vis_msp_o[28]), .B2(
        n2474), .C1(vis_r9_o[30]), .C2(n2338), .ZN(n5431) );
  OAI22_X1 U4800 ( .A1(n660), .A2(n2814), .B1(n4337), .B2(n4338), .ZN(n3797)
         );
  OAI211_X1 U4801 ( .C1(n4176), .C2(n8118), .A(n2447), .B(n4339), .ZN(n4338)
         );
  OAI221_X1 U4802 ( .B1(n640), .B2(n3593), .C1(n2468), .C2(n6253), .A(n4340), 
        .ZN(n4337) );
  AOI222_X1 U4803 ( .A1(vis_r8_o[31]), .A2(n2336), .B1(vis_msp_o[29]), .B2(
        n2474), .C1(vis_r9_o[31]), .C2(n2338), .ZN(n4339) );
  OAI221_X1 U4804 ( .B1(n1537), .B2(HADDR[8]), .C1(n7363), .C2(N701), .A(n128), 
        .ZN(n7735) );
  NAND4_X1 U4805 ( .A1(n2628), .A2(n4946), .A3(n4947), .A4(n4948), .ZN(n4168)
         );
  NAND2_X1 U4806 ( .A1(n599), .A2(n8195), .ZN(n4946) );
  AOI222_X1 U4807 ( .A1(vis_r10_o[23]), .A2(n617), .B1(vis_r11_o[23]), .B2(
        n4862), .C1(vis_r9_o[23]), .C2(n602), .ZN(n4947) );
  AOI221_X1 U4808 ( .B1(vis_r14_o[23]), .B2(n468), .C1(vis_r8_o[23]), .C2(
        n4856), .A(n4949), .ZN(n4948) );
  NAND4_X1 U4809 ( .A1(n2635), .A2(n4979), .A3(n4980), .A4(n4981), .ZN(n4800)
         );
  NAND2_X1 U4810 ( .A1(n4864), .A2(n3280), .ZN(n4979) );
  AOI222_X1 U4811 ( .A1(vis_r10_o[17]), .A2(n617), .B1(vis_r11_o[17]), .B2(
        n4862), .C1(vis_r9_o[17]), .C2(n602), .ZN(n4980) );
  AOI221_X1 U4812 ( .B1(vis_r14_o[17]), .B2(n468), .C1(vis_r8_o[17]), .C2(
        n4856), .A(n4982), .ZN(n4981) );
  NAND4_X1 U4813 ( .A1(n4141), .A2(n1840), .A3(n197), .A4(n198), .ZN(n187) );
  AND2_X1 U4814 ( .A1(N701), .A2(n203), .ZN(n197) );
  NOR4_X1 U4815 ( .A1(n199), .A2(n200), .A3(n201), .A4(n202), .ZN(n198) );
  NAND2_X1 U4816 ( .A1(n6048), .A2(n6049), .ZN(n4664) );
  AOI221_X1 U4817 ( .B1(vis_r2_o[20]), .B2(n6003), .C1(vis_r0_o[20]), .C2(n547), .A(n6051), .ZN(n6048) );
  AOI221_X1 U4818 ( .B1(vis_r3_o[20]), .B2(n567), .C1(vis_r7_o[20]), .C2(n5999), .A(n6050), .ZN(n6049) );
  OAI22_X1 U4819 ( .A1(n6006), .A2(n8221), .B1(n6007), .B2(n8209), .ZN(n6051)
         );
  OAI22_X1 U4820 ( .A1(n683), .A2(n8099), .B1(n2331), .B2(n2362), .ZN(Ecqhu6)
         );
  OAI22_X1 U4821 ( .A1(n683), .A2(n8093), .B1(n2205), .B2(n2362), .ZN(Lyphu6)
         );
  OAI22_X1 U4822 ( .A1(n683), .A2(n8091), .B1(n2327), .B2(n2362), .ZN(Meshu6)
         );
  OAI22_X1 U4823 ( .A1(n683), .A2(n8087), .B1(n2274), .B2(n2362), .ZN(P7qhu6)
         );
  OAI22_X1 U4824 ( .A1(n682), .A2(n8080), .B1(n2323), .B2(n2362), .ZN(Tgqhu6)
         );
  OAI22_X1 U4825 ( .A1(n767), .A2(n8073), .B1(n2340), .B2(n764), .ZN(D1qhu6)
         );
  OAI22_X1 U4826 ( .A1(n767), .A2(n8072), .B1(n2311), .B2(n2218), .ZN(Dnphu6)
         );
  OAI22_X1 U4827 ( .A1(n767), .A2(n8068), .B1(n2331), .B2(n764), .ZN(Haqhu6)
         );
  OAI22_X1 U4828 ( .A1(n768), .A2(n8062), .B1(n2205), .B2(n764), .ZN(Owphu6)
         );
  OAI22_X1 U4830 ( .A1(n768), .A2(n8061), .B1(n2327), .B2(n764), .ZN(Pcshu6)
         );
  OAI22_X1 U4831 ( .A1(n767), .A2(n8057), .B1(n2274), .B2(n2218), .ZN(S5qhu6)
         );
  OAI22_X1 U4832 ( .A1(n768), .A2(n8018), .B1(n2323), .B2(n2218), .ZN(Weqhu6)
         );
  OAI22_X1 U4833 ( .A1(n685), .A2(n6153), .B1(n2205), .B2(n684), .ZN(Hwphu6)
         );
  OAI22_X1 U4834 ( .A1(n685), .A2(n6152), .B1(n2327), .B2(n684), .ZN(Icshu6)
         );
  OAI22_X1 U4835 ( .A1(n685), .A2(n6144), .B1(n2274), .B2(n684), .ZN(L5qhu6)
         );
  OAI22_X1 U4836 ( .A1(n686), .A2(n6124), .B1(n2323), .B2(n2348), .ZN(Peqhu6)
         );
  OAI22_X1 U4837 ( .A1(n685), .A2(n6105), .B1(n2340), .B2(n2348), .ZN(W0qhu6)
         );
  OAI22_X1 U4838 ( .A1(n685), .A2(n6104), .B1(n2311), .B2(n2348), .ZN(Wmphu6)
         );
  OAI22_X1 U4839 ( .A1(n775), .A2(n5892), .B1(n2274), .B2(n2214), .ZN(E5qhu6)
         );
  OAI22_X1 U4840 ( .A1(n775), .A2(n5886), .B1(n2323), .B2(n771), .ZN(Ieqhu6)
         );
  OAI22_X1 U4841 ( .A1(n772), .A2(n5872), .B1(n2327), .B2(n2214), .ZN(Ofshu6)
         );
  OAI22_X1 U4842 ( .A1(n775), .A2(n5860), .B1(n2340), .B2(n2214), .ZN(P0qhu6)
         );
  OAI22_X1 U4843 ( .A1(n775), .A2(n5859), .B1(n2311), .B2(n2214), .ZN(Pmphu6)
         );
  OAI22_X1 U4844 ( .A1(n772), .A2(n5839), .B1(n2331), .B2(n2214), .ZN(T9qhu6)
         );
  OAI22_X1 U4845 ( .A1(n683), .A2(n4008), .B1(n2311), .B2(n2362), .ZN(Apphu6)
         );
  OAI22_X1 U4846 ( .A1(n775), .A2(n3614), .B1(n2205), .B2(n2214), .ZN(Awphu6)
         );
  OAI22_X1 U4847 ( .A1(n685), .A2(n3039), .B1(n2331), .B2(n2348), .ZN(Aaqhu6)
         );
  OAI22_X1 U4848 ( .A1(n682), .A2(n2816), .B1(n2340), .B2(n2362), .ZN(A3qhu6)
         );
  NAND4_X1 U4849 ( .A1(n5254), .A2(n455), .A3(n457), .A4(n3114), .ZN(n1599) );
  OAI221_X1 U4850 ( .B1(n3784), .B2(n4454), .C1(n4459), .C2(n5259), .A(n5260), 
        .ZN(n5254) );
  OAI21_X1 U4851 ( .B1(n7615), .B2(n5261), .A(n5262), .ZN(n5259) );
  AOI22_X1 U4852 ( .A1(n6126), .A2(n7623), .B1(n4465), .B2(n6735), .ZN(n6332)
         );
  NAND2_X1 U4853 ( .A1(n7527), .A2(n2807), .ZN(n3099) );
  OAI221_X1 U4854 ( .B1(n1544), .B2(n2513), .C1(n458), .C2(n3875), .A(n209), 
        .ZN(n7739) );
  AOI221_X1 U4855 ( .B1(n934), .B2(n211), .C1(Zsfpw6[30]), .C2(n931), .A(n213), 
        .ZN(n209) );
  NOR2_X1 U4856 ( .A1(n5105), .A2(vis_ipsr_o[5]), .ZN(n5888) );
  NOR2_X1 U4857 ( .A1(n5126), .A2(vis_ipsr_o[4]), .ZN(n5879) );
  OAI22_X1 U4858 ( .A1(n7636), .A2(n3677), .B1(n7561), .B2(n2472), .ZN(n5844)
         );
  OAI221_X1 U4859 ( .B1(n1537), .B2(n129), .C1(n7371), .C2(N701), .A(n128), 
        .ZN(n7732) );
  XNOR2_X1 U4860 ( .A(HADDR[7]), .B(HADDR[2]), .ZN(n129) );
  OAI22_X1 U4861 ( .A1(n7608), .A2(n4121), .B1(n7674), .B2(n2426), .ZN(n5843)
         );
  OAI221_X1 U4862 ( .B1(n1573), .B2(n1849), .C1(n7432), .C2(n180), .A(n1844), 
        .ZN(n7742) );
  INV_X1 U4863 ( .A(n227), .ZN(n1844) );
  OAI222_X1 U4864 ( .A1(n1847), .A2(n2729), .B1(n2133), .B2(n6727), .C1(n220), 
        .C2(n4761), .ZN(n227) );
  OAI221_X1 U4865 ( .B1(n1529), .B2(n1849), .C1(n7333), .C2(n180), .A(n181), 
        .ZN(n7736) );
  AOI222_X1 U4866 ( .A1(n182), .A2(vis_apsr_o[3]), .B1(n183), .B2(n3879), .C1(
        n1852), .C2(vis_pc_o[30]), .ZN(n181) );
  OAI221_X1 U4867 ( .B1(n1545), .B2(n1849), .C1(n7658), .C2(n180), .A(n1843), 
        .ZN(n7740) );
  INV_X1 U4868 ( .A(n216), .ZN(n1843) );
  OAI222_X1 U4869 ( .A1(n1847), .A2(n2778), .B1(n2133), .B2(n6897), .C1(n220), 
        .C2(n3124), .ZN(n216) );
  OAI22_X1 U4870 ( .A1(n7634), .A2(n3639), .B1(n7639), .B2(n4843), .ZN(n5850)
         );
  OAI21_X1 U4871 ( .B1(n7332), .B2(n4533), .A(n4534), .ZN(n2946) );
  AOI22_X1 U4872 ( .A1(vis_apsr_o[1]), .A2(n3067), .B1(n4536), .B2(n4537), 
        .ZN(n4533) );
  NAND2_X1 U4873 ( .A1(n7332), .A2(Nxkbx6[33]), .ZN(n4534) );
  INV_X1 U4874 ( .A(n4536), .ZN(n3067) );
  INV_X1 U4875 ( .A(n5836), .ZN(n3940) );
  AOI221_X1 U4876 ( .B1(n8255), .B2(n3983), .C1(n8160), .C2(n3955), .A(n5837), 
        .ZN(n5836) );
  OAI22_X1 U4877 ( .A1(n4013), .A2(n7677), .B1(n3644), .B2(n6773), .ZN(n5837)
         );
  OAI22_X1 U4878 ( .A1(n7356), .A2(n5648), .B1(n7527), .B2(n2807), .ZN(n5646)
         );
  OAI211_X1 U4879 ( .C1(n4504), .C2(n5937), .A(n2436), .B(n5700), .ZN(n5697)
         );
  AOI22_X1 U4880 ( .A1(vis_psp_o[25]), .A2(n229), .B1(vis_r12_o[27]), .B2(
        n4290), .ZN(n5700) );
  OAI211_X1 U4881 ( .C1(n4504), .C2(n5948), .A(n2427), .B(n4505), .ZN(n4499)
         );
  AOI22_X1 U4882 ( .A1(vis_psp_o[23]), .A2(n229), .B1(vis_r12_o[25]), .B2(
        n4290), .ZN(n4505) );
  OAI211_X1 U4883 ( .C1(n4504), .C2(n5961), .A(n2432), .B(n4684), .ZN(n4681)
         );
  AOI22_X1 U4884 ( .A1(vis_psp_o[24]), .A2(n229), .B1(vis_r12_o[26]), .B2(
        n4290), .ZN(n4684) );
  OAI22_X1 U4885 ( .A1(n7678), .A2(n3597), .B1(n7616), .B2(n1636), .ZN(n5842)
         );
  OAI221_X1 U4886 ( .B1(n1537), .B2(n130), .C1(n7548), .C2(N701), .A(n128), 
        .ZN(n7733) );
  XNOR2_X1 U4887 ( .A(HADDR[3]), .B(HADDR[5]), .ZN(n130) );
  OAI221_X1 U4888 ( .B1(n1537), .B2(n127), .C1(n7398), .C2(N701), .A(n128), 
        .ZN(n7731) );
  XNOR2_X1 U4889 ( .A(HADDR[3]), .B(HADDR[10]), .ZN(n127) );
  NAND2_X1 U4890 ( .A1(n6411), .A2(n6412), .ZN(n5324) );
  AOI221_X1 U4891 ( .B1(vis_r2_o[16]), .B2(n6003), .C1(vis_r0_o[16]), .C2(n547), .A(n6414), .ZN(n6411) );
  AOI221_X1 U4892 ( .B1(vis_r3_o[16]), .B2(n567), .C1(vis_r7_o[16]), .C2(n5999), .A(n6413), .ZN(n6412) );
  OAI22_X1 U4893 ( .A1(n6006), .A2(n6478), .B1(n6007), .B2(n5386), .ZN(n6414)
         );
  NAND2_X1 U4894 ( .A1(n6073), .A2(n6074), .ZN(n5328) );
  AOI221_X1 U4895 ( .B1(vis_r2_o[24]), .B2(n6003), .C1(vis_r0_o[24]), .C2(n547), .A(n6076), .ZN(n6073) );
  AOI221_X1 U4896 ( .B1(vis_r3_o[24]), .B2(n567), .C1(vis_r7_o[24]), .C2(n5999), .A(n6075), .ZN(n6074) );
  OAI22_X1 U4897 ( .A1(n6006), .A2(n6504), .B1(n6007), .B2(n5419), .ZN(n6076)
         );
  NOR2_X1 U4898 ( .A1(vis_ipsr_o[2]), .A2(vis_ipsr_o[3]), .ZN(n5880) );
  AND3_X1 U4899 ( .A1(vis_ipsr_o[3]), .A2(n5111), .A3(n5888), .ZN(n5878) );
  AND3_X1 U4900 ( .A1(vis_ipsr_o[2]), .A2(vis_ipsr_o[3]), .A3(n5888), .ZN(
        n5869) );
  AND3_X1 U4901 ( .A1(vis_ipsr_o[2]), .A2(n5088), .A3(n5888), .ZN(n5861) );
  OAI211_X1 U4902 ( .C1(n6357), .C2(n6358), .A(n8259), .B(n8257), .ZN(n6126)
         );
  NAND2_X1 U4903 ( .A1(n8240), .A2(n8250), .ZN(n6358) );
  AOI22_X1 U4904 ( .A1(n6359), .A2(n7623), .B1(n7624), .B2(n4467), .ZN(n6357)
         );
  AOI21_X1 U4905 ( .B1(n6777), .B2(n4466), .A(n6735), .ZN(n6359) );
  OAI22_X1 U4906 ( .A1(n3875), .A2(n2297), .B1(n701), .B2(n1529), .ZN(R9ohu6)
         );
  OAI22_X1 U4907 ( .A1(n3875), .A2(n733), .B1(n736), .B2(n1529), .ZN(M9ohu6)
         );
  AND3_X1 U4908 ( .A1(vis_ipsr_o[3]), .A2(n5111), .A3(n5879), .ZN(n5864) );
  OAI21_X1 U4909 ( .B1(n7703), .B2(n5787), .A(n5788), .ZN(n5784) );
  NAND3_X1 U4910 ( .A1(n4350), .A2(n8175), .A3(n7703), .ZN(n5788) );
  AND3_X1 U4911 ( .A1(vis_ipsr_o[2]), .A2(n5088), .A3(n5879), .ZN(n5870) );
  AND3_X1 U4912 ( .A1(vis_ipsr_o[2]), .A2(vis_ipsr_o[3]), .A3(n5879), .ZN(
        n5863) );
  AND2_X1 U4913 ( .A1(Ntkbx6[25]), .A2(n2295), .ZN(Ysihu6) );
  OAI22_X1 U4914 ( .A1(n697), .A2(n1603), .B1(n696), .B2(n4799), .ZN(n2295) );
  AND2_X1 U4915 ( .A1(Ntkbx6[22]), .A2(n5062), .ZN(Apihu6) );
  OAI22_X1 U4916 ( .A1(n697), .A2(n1616), .B1(n696), .B2(n4766), .ZN(n5062) );
  AND2_X1 U4917 ( .A1(Ntkbx6[26]), .A2(n3944), .ZN(Guihu6) );
  OAI22_X1 U4918 ( .A1(n697), .A2(n1596), .B1(n696), .B2(n4797), .ZN(n3944) );
  AND2_X1 U4919 ( .A1(Ntkbx6[24]), .A2(n2775), .ZN(Qrihu6) );
  OAI22_X1 U4920 ( .A1(n701), .A2(n1606), .B1(n696), .B2(n4764), .ZN(n2775) );
  AND2_X1 U4921 ( .A1(Ntkbx6[23]), .A2(n3776), .ZN(Iqihu6) );
  OAI22_X1 U4922 ( .A1(n701), .A2(n1610), .B1(n696), .B2(n4765), .ZN(n3776) );
  NAND2_X1 U4923 ( .A1(n3283), .A2(n5200), .ZN(n2154) );
  OAI211_X1 U4924 ( .C1(n5201), .C2(n4548), .A(n3285), .B(n5202), .ZN(n5200)
         );
  AOI22_X1 U4925 ( .A1(n1978), .A2(n2510), .B1(n7507), .B2(n529), .ZN(n5201)
         );
  NAND3_X1 U4926 ( .A1(n1978), .A2(n4548), .A3(n2511), .ZN(n5202) );
  AOI21_X1 U4927 ( .B1(n7619), .B2(n4470), .A(n7673), .ZN(n6256) );
  NAND2_X1 U4928 ( .A1(n6227), .A2(n6228), .ZN(n6145) );
  OAI21_X1 U4929 ( .B1(n7595), .B2(n7581), .A(n6233), .ZN(n6227) );
  OAI221_X1 U4931 ( .B1(n3119), .B2(n4435), .C1(n6217), .C2(n6216), .A(n6230), 
        .ZN(n6228) );
  INV_X1 U4932 ( .A(n6226), .ZN(n3119) );
  NAND2_X1 U4933 ( .A1(n6044), .A2(n6045), .ZN(n5329) );
  AOI221_X1 U4934 ( .B1(vis_r2_o[23]), .B2(n6003), .C1(vis_r0_o[23]), .C2(n547), .A(n6047), .ZN(n6044) );
  AOI221_X1 U4935 ( .B1(vis_r3_o[23]), .B2(n567), .C1(vis_r7_o[23]), .C2(n5999), .A(n6046), .ZN(n6045) );
  OAI22_X1 U4936 ( .A1(n6006), .A2(n6452), .B1(n6007), .B2(n5394), .ZN(n6047)
         );
  NAND2_X1 U4937 ( .A1(n6061), .A2(n6062), .ZN(n5337) );
  AOI221_X1 U4938 ( .B1(vis_r2_o[27]), .B2(n6003), .C1(vis_r0_o[27]), .C2(n547), .A(n6064), .ZN(n6061) );
  AOI221_X1 U4939 ( .B1(vis_r3_o[27]), .B2(n567), .C1(vis_r7_o[27]), .C2(n5999), .A(n6063), .ZN(n6062) );
  OAI22_X1 U4940 ( .A1(n6006), .A2(n6560), .B1(n6007), .B2(n5451), .ZN(n6064)
         );
  NAND2_X1 U4941 ( .A1(n6415), .A2(n6416), .ZN(n5472) );
  AOI221_X1 U4942 ( .B1(vis_r2_o[17]), .B2(n6003), .C1(vis_r0_o[17]), .C2(n547), .A(n6418), .ZN(n6415) );
  AOI221_X1 U4943 ( .B1(vis_r3_o[17]), .B2(n567), .C1(vis_r7_o[17]), .C2(n5999), .A(n6417), .ZN(n6416) );
  OAI22_X1 U4944 ( .A1(n6006), .A2(n6564), .B1(n6007), .B2(n5460), .ZN(n6418)
         );
  NAND2_X1 U4945 ( .A1(n6407), .A2(n6408), .ZN(n5290) );
  AOI221_X1 U4946 ( .B1(vis_r2_o[19]), .B2(n6003), .C1(vis_r0_o[19]), .C2(n547), .A(n6410), .ZN(n6407) );
  AOI221_X1 U4947 ( .B1(vis_r3_o[19]), .B2(n567), .C1(vis_r7_o[19]), .C2(n5999), .A(n6409), .ZN(n6408) );
  OAI22_X1 U4948 ( .A1(n6006), .A2(n6518), .B1(n6007), .B2(n5427), .ZN(n6410)
         );
  NAND2_X1 U4949 ( .A1(n6069), .A2(n6070), .ZN(n5501) );
  AOI221_X1 U4950 ( .B1(vis_r2_o[25]), .B2(n6003), .C1(vis_r0_o[25]), .C2(n547), .A(n6072), .ZN(n6069) );
  AOI221_X1 U4951 ( .B1(vis_r3_o[25]), .B2(n567), .C1(vis_r7_o[25]), .C2(n5999), .A(n6071), .ZN(n6070) );
  OAI22_X1 U4952 ( .A1(n6006), .A2(n6588), .B1(n6007), .B2(n5326), .ZN(n6072)
         );
  NAND2_X1 U4953 ( .A1(n6065), .A2(n6066), .ZN(n5336) );
  AOI221_X1 U4954 ( .B1(vis_r2_o[26]), .B2(n6003), .C1(vis_r0_o[26]), .C2(n547), .A(n6068), .ZN(n6065) );
  AOI221_X1 U4955 ( .B1(vis_r3_o[26]), .B2(n567), .C1(vis_r7_o[26]), .C2(n5999), .A(n6067), .ZN(n6066) );
  OAI22_X1 U4956 ( .A1(n6006), .A2(n6395), .B1(n6007), .B2(n5369), .ZN(n6068)
         );
  AND2_X1 U4957 ( .A1(Nvkbx6[24]), .A2(n4050), .ZN(Eblhu6) );
  OAI22_X1 U4958 ( .A1(n733), .A2(n4764), .B1(n736), .B2(n1606), .ZN(n4050) );
  AND2_X1 U4959 ( .A1(Nvkbx6[25]), .A2(n3224), .ZN(Lclhu6) );
  OAI22_X1 U4960 ( .A1(n2264), .A2(n4799), .B1(n736), .B2(n1603), .ZN(n3224)
         );
  AND2_X1 U4961 ( .A1(Nvkbx6[26]), .A2(n2687), .ZN(Sdlhu6) );
  OAI22_X1 U4962 ( .A1(n733), .A2(n4797), .B1(n736), .B2(n1596), .ZN(n2687) );
  AND2_X1 U4963 ( .A1(Nvkbx6[22]), .A2(n3011), .ZN(O8lhu6) );
  OAI22_X1 U4964 ( .A1(n733), .A2(n4766), .B1(n736), .B2(n1616), .ZN(n3011) );
  AND2_X1 U4965 ( .A1(Ntkbx6[30]), .A2(n3069), .ZN(Mzihu6) );
  OAI22_X1 U4966 ( .A1(n3124), .A2(n696), .B1(n697), .B2(n1545), .ZN(n3069) );
  AND2_X1 U4967 ( .A1(Nvkbx6[30]), .A2(n2542), .ZN(Uilhu6) );
  OAI22_X1 U4968 ( .A1(n3124), .A2(n733), .B1(n734), .B2(n1545), .ZN(n2542) );
  AOI21_X1 U4969 ( .B1(n7621), .B2(n8244), .A(n7637), .ZN(n6356) );
  OAI211_X1 U4970 ( .C1(n6295), .C2(n6296), .A(n8227), .B(n8225), .ZN(n6135)
         );
  NAND2_X1 U4972 ( .A1(n3669), .A2(n8148), .ZN(n6296) );
  AOI22_X1 U4973 ( .A1(n6297), .A2(n7552), .B1(n7553), .B2(n8232), .ZN(n6295)
         );
  AOI21_X1 U4974 ( .B1(n7551), .B2(n8242), .A(n7636), .ZN(n6297) );
  OAI211_X1 U4975 ( .C1(n6250), .C2(n6251), .A(n8280), .B(n8278), .ZN(n6245)
         );
  NAND2_X1 U4976 ( .A1(n3037), .A2(n8147), .ZN(n6251) );
  AOI22_X1 U4977 ( .A1(n6252), .A2(n7617), .B1(n7618), .B2(n8234), .ZN(n6250)
         );
  AOI21_X1 U4978 ( .B1(n6710), .B2(n8247), .A(n6775), .ZN(n6252) );
  OAI22_X1 U4979 ( .A1(n686), .A2(n8277), .B1(n2321), .B2(n2348), .ZN(Aiphu6)
         );
  OAI22_X1 U4980 ( .A1(n683), .A2(n8275), .B1(n2321), .B2(n2362), .ZN(Ekphu6)
         );
  OAI22_X1 U4981 ( .A1(n683), .A2(n8100), .B1(n2404), .B2(n2362), .ZN(C1thu6)
         );
  OAI22_X1 U4982 ( .A1(n767), .A2(n8069), .B1(n2404), .B2(n2218), .ZN(Gwshu6)
         );
  OAI22_X1 U4983 ( .A1(n686), .A2(n6167), .B1(n2239), .B2(n2348), .ZN(Evshu6)
         );
  OAI22_X1 U4984 ( .A1(n686), .A2(n3031), .B1(n2213), .B2(n2348), .ZN(Aurhu6)
         );
  OAI22_X1 U4985 ( .A1(n682), .A2(n8095), .B1(n2271), .B2(n2362), .ZN(J1thu6)
         );
  OAI22_X1 U4986 ( .A1(n768), .A2(n8063), .B1(n2271), .B2(n764), .ZN(Nwshu6)
         );
  OAI22_X1 U4987 ( .A1(n685), .A2(n5993), .B1(n2271), .B2(n2348), .ZN(Xushu6)
         );
  OAI22_X1 U4988 ( .A1(n775), .A2(n5820), .B1(n2271), .B2(n2214), .ZN(Zashu6)
         );
  OAI22_X1 U4989 ( .A1(n767), .A2(n8273), .B1(n2321), .B2(n764), .ZN(Hiphu6)
         );
  OAI22_X1 U4990 ( .A1(n775), .A2(n8265), .B1(n2321), .B2(n2214), .ZN(Thphu6)
         );
  OAI22_X1 U4991 ( .A1(n683), .A2(n8085), .B1(n2239), .B2(n2362), .ZN(Q1thu6)
         );
  OAI22_X1 U4992 ( .A1(n767), .A2(n8019), .B1(n2239), .B2(n2218), .ZN(Uwshu6)
         );
  OAI22_X1 U4993 ( .A1(n775), .A2(n5814), .B1(n2239), .B2(n2214), .ZN(Zoshu6)
         );
  OAI22_X1 U4994 ( .A1(n683), .A2(n8077), .B1(n2217), .B2(n2362), .ZN(V0thu6)
         );
  OAI22_X1 U4995 ( .A1(n768), .A2(n7824), .B1(n2217), .B2(n2218), .ZN(Zvshu6)
         );
  OAI22_X1 U4996 ( .A1(n685), .A2(n6146), .B1(n2217), .B2(n684), .ZN(Jushu6)
         );
  OAI22_X1 U4997 ( .A1(n772), .A2(n5829), .B1(n2217), .B2(n2214), .ZN(Wrrhu6)
         );
  OAI22_X1 U4998 ( .A1(n686), .A2(n6120), .B1(n2404), .B2(n2348), .ZN(Qushu6)
         );
  OAI22_X1 U4999 ( .A1(n775), .A2(n5849), .B1(n2404), .B2(n2214), .ZN(Rsrhu6)
         );
  OAI22_X1 U5000 ( .A1(n683), .A2(n8098), .B1(n2213), .B2(n681), .ZN(Ewrhu6)
         );
  OAI22_X1 U5001 ( .A1(n767), .A2(n8067), .B1(n2213), .B2(n764), .ZN(Hurhu6)
         );
  OAI22_X1 U5002 ( .A1(n775), .A2(n5811), .B1(n2213), .B2(n2214), .ZN(Zwrhu6)
         );
  OAI22_X1 U5003 ( .A1(n683), .A2(n8083), .B1(n2335), .B2(n2362), .ZN(Q9shu6)
         );
  OAI22_X1 U5004 ( .A1(n768), .A2(n8038), .B1(n2335), .B2(n2218), .ZN(T7shu6)
         );
  OAI22_X1 U5005 ( .A1(n686), .A2(n6129), .B1(n2335), .B2(n684), .ZN(M7shu6)
         );
  OAI22_X1 U5006 ( .A1(n775), .A2(n5848), .B1(n2335), .B2(n2214), .ZN(Sashu6)
         );
  OAI22_X1 U5007 ( .A1(n3294), .A2(n2812), .B1(n3457), .B2(n2609), .ZN(Kgphu6)
         );
  AOI222_X1 U5008 ( .A1(n101), .A2(n3458), .B1(n97), .B2(n2940), .C1(n99), 
        .C2(n211), .ZN(n3457) );
  OAI22_X1 U5009 ( .A1(n7694), .A2(n109), .B1(n110), .B2(n111), .ZN(n7728) );
  NOR2_X1 U5010 ( .A1(n109), .A2(N701), .ZN(n110) );
  NOR2_X1 U5011 ( .A1(n4140), .A2(n113), .ZN(n109) );
  OAI22_X1 U5012 ( .A1(n7291), .A2(n122), .B1(n123), .B2(n124), .ZN(n7730) );
  NOR2_X1 U5013 ( .A1(n122), .A2(N701), .ZN(n123) );
  NOR2_X1 U5014 ( .A1(n125), .A2(n4140), .ZN(n122) );
  OAI22_X1 U5015 ( .A1(n7392), .A2(N701), .B1(n194), .B2(n187), .ZN(n7738) );
  NOR2_X1 U5016 ( .A1(n204), .A2(n205), .ZN(n194) );
  OAI22_X1 U5017 ( .A1(n7380), .A2(N701), .B1(n186), .B2(n187), .ZN(n7737) );
  NOR2_X1 U5018 ( .A1(n188), .A2(n189), .ZN(n186) );
  OAI22_X1 U5019 ( .A1(n6769), .A2(n2152), .B1(n2153), .B2(n1989), .ZN(n7213)
         );
  NAND3_X1 U5020 ( .A1(n952), .A2(n3895), .A3(n7490), .ZN(n3892) );
  NAND2_X1 U5021 ( .A1(n6419), .A2(n6420), .ZN(n5983) );
  AOI221_X1 U5022 ( .B1(vis_r2_o[18]), .B2(n6003), .C1(vis_r0_o[18]), .C2(n547), .A(n6422), .ZN(n6419) );
  AOI221_X1 U5023 ( .B1(vis_r3_o[18]), .B2(n567), .C1(vis_r7_o[18]), .C2(n5999), .A(n6421), .ZN(n6420) );
  OAI22_X1 U5024 ( .A1(n6006), .A2(n8178), .B1(n6007), .B2(n8182), .ZN(n6422)
         );
  OAI222_X1 U5025 ( .A1(n2330), .A2(n3900), .B1(n3907), .B2(n242), .C1(n1804), 
        .C2(n661), .ZN(\eq_3147/A[0] ) );
  NAND2_X1 U5026 ( .A1(n1430), .A2(vis_pc_o[0]), .ZN(n3908) );
  AND2_X1 U5027 ( .A1(n6909), .A2(HMASTER), .ZN(n3923) );
  AND2_X1 U5028 ( .A1(n4915), .A2(n4916), .ZN(n2634) );
  AOI221_X1 U5029 ( .B1(vis_r5_o[18]), .B2(n4867), .C1(vis_r4_o[18]), .C2(
        n4868), .A(n4917), .ZN(n4916) );
  AOI221_X1 U5030 ( .B1(vis_r6_o[18]), .B2(n4872), .C1(vis_r1_o[18]), .C2(
        n4873), .A(n4918), .ZN(n4915) );
  OAI22_X1 U5031 ( .A1(n4870), .A2(n8188), .B1(n4871), .B2(n8185), .ZN(n4917)
         );
  AND2_X1 U5032 ( .A1(n5618), .A2(n5619), .ZN(n2633) );
  AOI221_X1 U5033 ( .B1(vis_r6_o[19]), .B2(n576), .C1(vis_r1_o[19]), .C2(n4873), .A(n5621), .ZN(n5618) );
  AOI221_X1 U5034 ( .B1(vis_r5_o[19]), .B2(n582), .C1(vis_r4_o[19]), .C2(n4868), .A(n5620), .ZN(n5619) );
  OAI22_X1 U5035 ( .A1(n572), .A2(n7821), .B1(n4876), .B2(n5522), .ZN(n5621)
         );
  AND2_X1 U5036 ( .A1(n5007), .A2(n5008), .ZN(n2630) );
  AOI221_X1 U5037 ( .B1(vis_r6_o[21]), .B2(n4872), .C1(vis_r1_o[21]), .C2(
        n4873), .A(n5010), .ZN(n5007) );
  AOI221_X1 U5038 ( .B1(vis_r5_o[21]), .B2(n4867), .C1(vis_r4_o[21]), .C2(
        n4868), .A(n5009), .ZN(n5008) );
  OAI22_X1 U5039 ( .A1(n4875), .A2(n7802), .B1(n4876), .B2(n5485), .ZN(n5010)
         );
  AND2_X1 U5040 ( .A1(n4998), .A2(n4999), .ZN(n2631) );
  AOI221_X1 U5041 ( .B1(vis_r6_o[20]), .B2(n4872), .C1(vis_r1_o[20]), .C2(
        n4873), .A(n5001), .ZN(n4998) );
  AOI221_X1 U5042 ( .B1(vis_r5_o[20]), .B2(n4867), .C1(vis_r4_o[20]), .C2(
        n4868), .A(n5000), .ZN(n4999) );
  OAI22_X1 U5043 ( .A1(n4875), .A2(n8213), .B1(n4876), .B2(n8219), .ZN(n5001)
         );
  AND2_X1 U5044 ( .A1(n4983), .A2(n4984), .ZN(n2635) );
  AOI221_X1 U5045 ( .B1(vis_r6_o[17]), .B2(n4872), .C1(vis_r1_o[17]), .C2(
        n4873), .A(n4986), .ZN(n4983) );
  AOI221_X1 U5046 ( .B1(vis_r5_o[17]), .B2(n4867), .C1(vis_r4_o[17]), .C2(
        n4868), .A(n4985), .ZN(n4984) );
  OAI22_X1 U5047 ( .A1(n4875), .A2(n7745), .B1(n4876), .B2(n5532), .ZN(n4986)
         );
  AND2_X1 U5048 ( .A1(n5083), .A2(n5084), .ZN(n2636) );
  AOI221_X1 U5049 ( .B1(vis_r6_o[16]), .B2(n4872), .C1(vis_r1_o[16]), .C2(
        n4873), .A(n5086), .ZN(n5083) );
  AOI221_X1 U5050 ( .B1(vis_r5_o[16]), .B2(n4867), .C1(vis_r4_o[16]), .C2(
        n4868), .A(n5085), .ZN(n5084) );
  OAI22_X1 U5051 ( .A1(n4875), .A2(n7797), .B1(n4876), .B2(n5465), .ZN(n5086)
         );
  OAI211_X1 U5052 ( .C1(n6161), .C2(n6163), .A(n2227), .B(n3617), .ZN(n5456)
         );
  AOI22_X1 U5053 ( .A1(n6164), .A2(n6157), .B1(n6160), .B2(n4473), .ZN(n6163)
         );
  AOI21_X1 U5054 ( .B1(n7331), .B2(n2781), .A(n7257), .ZN(n6164) );
  INV_X1 U5055 ( .A(n6160), .ZN(n2781) );
  INV_X1 U5056 ( .A(n6232), .ZN(n3118) );
  AOI22_X1 U5057 ( .A1(n6233), .A2(n7605), .B1(n3120), .B2(n6778), .ZN(n6232)
         );
  INV_X1 U5058 ( .A(n5840), .ZN(n3931) );
  OAI222_X1 U5059 ( .A1(n3660), .A2(n6772), .B1(n3558), .B2(n7617), .C1(n2685), 
        .C2(n7673), .ZN(n5840) );
  INV_X1 U5060 ( .A(n5835), .ZN(n3947) );
  OAI22_X1 U5061 ( .A1(n2357), .A2(n6774), .B1(n3649), .B2(n7676), .ZN(n5835)
         );
  INV_X1 U5062 ( .A(n5833), .ZN(n3979) );
  OAI22_X1 U5063 ( .A1(n3778), .A2(n6778), .B1(n3742), .B2(n6702), .ZN(n5833)
         );
  AND2_X1 U5064 ( .A1(Nvkbx6[23]), .A2(n2441), .ZN(W9lhu6) );
  OAI22_X1 U5065 ( .A1(n2264), .A2(n4765), .B1(n734), .B2(n1610), .ZN(n2441)
         );
  OAI22_X1 U5066 ( .A1(n4441), .A2(n4442), .B1(n4453), .B2(n7607), .ZN(n6238)
         );
  INV_X1 U5067 ( .A(n6240), .ZN(n4441) );
  AOI21_X1 U5068 ( .B1(n7607), .B2(n4453), .A(n7674), .ZN(n6240) );
  AOI22_X1 U5069 ( .A1(n4850), .A2(n4649), .B1(n4851), .B2(n102), .ZN(n4849)
         );
  INV_X1 U5070 ( .A(n4909), .ZN(n4002) );
  INV_X1 U5071 ( .A(n4425), .ZN(n4379) );
  AOI22_X1 U5072 ( .A1(n4850), .A2(n4449), .B1(n4851), .B2(n4496), .ZN(n4919)
         );
  INV_X1 U5073 ( .A(n4988), .ZN(n3863) );
  INV_X1 U5074 ( .A(n4666), .ZN(n4378) );
  INV_X1 U5075 ( .A(n4603), .ZN(n3648) );
  INV_X1 U5076 ( .A(n4941), .ZN(n2728) );
  AOI22_X1 U5077 ( .A1(n4851), .A2(n4531), .B1(n4850), .B2(n4878), .ZN(n4877)
         );
  AOI22_X1 U5078 ( .A1(n4850), .A2(n4888), .B1(n4851), .B2(n3297), .ZN(n4887)
         );
  AOI22_X1 U5079 ( .A1(n4850), .A2(n4938), .B1(n4851), .B2(n4939), .ZN(n4937)
         );
  AOI22_X1 U5080 ( .A1(n4850), .A2(n4471), .B1(n4851), .B2(n3458), .ZN(n4889)
         );
  AOI22_X1 U5081 ( .A1(n4850), .A2(n4747), .B1(n4851), .B2(n4678), .ZN(n4957)
         );
  INV_X1 U5082 ( .A(n4471), .ZN(n2478) );
  AOI22_X1 U5083 ( .A1(n4850), .A2(n4955), .B1(n4851), .B2(n4956), .ZN(n4954)
         );
  NAND4_X1 U5084 ( .A1(n6769), .A2(n7354), .A3(n6770), .A4(n4353), .ZN(
        CODENSEQ) );
  AOI221_X1 U5085 ( .B1(n3533), .B2(n2234), .C1(n7532), .C2(n7493), .A(n4354), 
        .ZN(n4353) );
  NAND3_X1 U5086 ( .A1(n4355), .A2(n4356), .A3(n4357), .ZN(CODEHINTDE[2]) );
  NOR4_X1 U5087 ( .A1(n4358), .A2(n4359), .A3(n2894), .A4(n4360), .ZN(n4357)
         );
  AOI21_X1 U5088 ( .B1(n417), .B2(n1945), .A(n2870), .ZN(n4355) );
  AOI22_X1 U5089 ( .A1(n7492), .A2(n4363), .B1(n3123), .B2(n1903), .ZN(n4356)
         );
  AOI22_X1 U5090 ( .A1(n3895), .A2(n7418), .B1(n4118), .B2(n2395), .ZN(n918)
         );
  NAND4_X1 U5091 ( .A1(n4835), .A2(n4753), .A3(vis_pc_o[27]), .A4(n5242), .ZN(
        n1482) );
  NOR3_X1 U5092 ( .A1(n3875), .A2(n4761), .A3(n3124), .ZN(n5242) );
  NOR2_X1 U5093 ( .A1(n7516), .A2(n7514), .ZN(n1612) );
  AOI221_X1 U5094 ( .B1(n3360), .B2(n4717), .C1(n4691), .C2(HRDATA[12]), .A(
        n6083), .ZN(n4638) );
  OAI22_X1 U5095 ( .A1(n2712), .A2(n2176), .B1(n3104), .B2(n2402), .ZN(n6083)
         );
  AOI211_X1 U5096 ( .C1(n2227), .C2(n6681), .A(n2226), .B(n6108), .ZN(n5297)
         );
  NOR3_X1 U5097 ( .A1(n4229), .A2(n7497), .A3(n3766), .ZN(n1660) );
  AOI211_X1 U5098 ( .C1(n1592), .C2(n475), .A(n4572), .B(n1752), .ZN(n4369) );
  AOI22_X1 U5099 ( .A1(n4371), .A2(n2262), .B1(n1908), .B2(n476), .ZN(n4370)
         );
  OAI221_X1 U5100 ( .B1(n7518), .B2(n4372), .C1(n4572), .C2(n4732), .A(n4373), 
        .ZN(n4371) );
  OAI221_X1 U5101 ( .B1(n2396), .B2(n3104), .C1(n817), .C2(n2712), .A(n5443), 
        .ZN(n4527) );
  AOI22_X1 U5102 ( .A1(n4717), .A2(n3322), .B1(HRDATA[14]), .B2(n4691), .ZN(
        n5443) );
  AOI222_X1 U5103 ( .A1(n1110), .A2(n4705), .B1(n3349), .B2(n3725), .C1(n4691), 
        .C2(HRDATA[31]), .ZN(n4488) );
  OAI211_X1 U5104 ( .C1(n6384), .C2(n6363), .A(n3030), .B(n8142), .ZN(n6362)
         );
  AOI22_X1 U5105 ( .A1(n6385), .A2(n6772), .B1(n7565), .B2(n4487), .ZN(n6384)
         );
  AOI21_X1 U5106 ( .B1(n7566), .B2(n4482), .A(n7670), .ZN(n6385) );
  NOR3_X1 U5107 ( .A1(n4674), .A2(n7559), .A3(n4787), .ZN(n2568) );
  NAND4_X1 U5108 ( .A1(n2619), .A2(n4890), .A3(n4891), .A4(n4892), .ZN(n3458)
         );
  NAND2_X1 U5109 ( .A1(n599), .A2(n2814), .ZN(n4890) );
  AOI222_X1 U5110 ( .A1(vis_r10_o[31]), .A2(n4861), .B1(vis_r11_o[31]), .B2(
        n4862), .C1(vis_r9_o[31]), .C2(n602), .ZN(n4891) );
  AOI221_X1 U5111 ( .B1(vis_r14_o[31]), .B2(n5272), .C1(vis_r8_o[31]), .C2(
        n628), .A(n4893), .ZN(n4892) );
  NAND4_X1 U5112 ( .A1(n2620), .A2(n5434), .A3(n5435), .A4(n5436), .ZN(n3297)
         );
  NAND2_X1 U5113 ( .A1(n4864), .A2(n2779), .ZN(n5434) );
  AOI222_X1 U5114 ( .A1(vis_r10_o[30]), .A2(n4861), .B1(vis_r11_o[30]), .B2(
        n615), .C1(vis_r9_o[30]), .C2(n4863), .ZN(n5435) );
  AOI221_X1 U5115 ( .B1(vis_r14_o[30]), .B2(n5272), .C1(vis_r8_o[30]), .C2(
        n4856), .A(n5437), .ZN(n5436) );
  AOI22_X1 U5116 ( .A1(n3895), .A2(n7441), .B1(n4119), .B2(n2395), .ZN(n922)
         );
  NOR3_X1 U5117 ( .A1(n1364), .A2(n7480), .A3(n4116), .ZN(n1366) );
  NOR2_X1 U5118 ( .A1(n2256), .A2(n7399), .ZN(n1613) );
  NOR2_X1 U5119 ( .A1(n3008), .A2(n7414), .ZN(n1144) );
  NOR2_X1 U5120 ( .A1(n2260), .A2(n7510), .ZN(n1684) );
  OAI211_X1 U5121 ( .C1(n6400), .C2(n6401), .A(n8149), .B(n4293), .ZN(n6130)
         );
  NAND2_X1 U5122 ( .A1(n8237), .A2(n8239), .ZN(n6401) );
  AOI22_X1 U5123 ( .A1(n6402), .A2(n6758), .B1(n7558), .B2(n8159), .ZN(n6400)
         );
  AOI21_X1 U5124 ( .B1(n7557), .B2(n8161), .A(n7678), .ZN(n6402) );
  OAI211_X1 U5125 ( .C1(n6298), .C2(n6299), .A(n8203), .B(n8201), .ZN(n6137)
         );
  NAND2_X1 U5126 ( .A1(n8294), .A2(n8292), .ZN(n6299) );
  AOI22_X1 U5127 ( .A1(n6300), .A2(n6759), .B1(n7555), .B2(n8157), .ZN(n6298)
         );
  AOI21_X1 U5128 ( .B1(n7554), .B2(n8158), .A(n7675), .ZN(n6300) );
  OAI211_X1 U5129 ( .C1(n6282), .C2(n6283), .A(n4005), .B(n8139), .ZN(n6275)
         );
  NAND2_X1 U5130 ( .A1(n3310), .A2(n8151), .ZN(n6283) );
  AOI22_X1 U5131 ( .A1(n6284), .A2(n7561), .B1(n7562), .B2(n8231), .ZN(n6282)
         );
  AOI21_X1 U5132 ( .B1(n6712), .B2(n8245), .A(n6773), .ZN(n6284) );
  AOI211_X1 U5133 ( .C1(n8151), .C2(n2852), .A(n4785), .B(n4786), .ZN(n865) );
  OAI222_X1 U5134 ( .A1(n8358), .A2(n4788), .B1(n2202), .B2(n7367), .C1(n1893), 
        .C2(n7368), .ZN(n4786) );
  OAI22_X1 U5135 ( .A1(n756), .A2(n2825), .B1(n4730), .B2(n7588), .ZN(n4785)
         );
  INV_X1 U5136 ( .A(STCALIB[17]), .ZN(n8358) );
  NAND4_X1 U5137 ( .A1(n2623), .A2(n5117), .A3(n5118), .A4(n5119), .ZN(n102)
         );
  NAND2_X1 U5138 ( .A1(n4864), .A2(n8261), .ZN(n5117) );
  AOI222_X1 U5139 ( .A1(vis_r10_o[28]), .A2(n617), .B1(vis_r11_o[28]), .B2(
        n615), .C1(vis_r9_o[28]), .C2(n4863), .ZN(n5118) );
  AOI221_X1 U5140 ( .B1(vis_r14_o[28]), .B2(n5272), .C1(vis_r8_o[28]), .C2(
        n4856), .A(n5120), .ZN(n5119) );
  NAND4_X1 U5141 ( .A1(n2622), .A2(n4879), .A3(n4880), .A4(n4881), .ZN(n4531)
         );
  NAND2_X1 U5142 ( .A1(n599), .A2(n8204), .ZN(n4879) );
  AOI222_X1 U5143 ( .A1(vis_r10_o[29]), .A2(n617), .B1(vis_r11_o[29]), .B2(
        n4862), .C1(vis_r9_o[29]), .C2(n602), .ZN(n4880) );
  AOI221_X1 U5144 ( .B1(vis_r14_o[29]), .B2(n5272), .C1(vis_r8_o[29]), .C2(
        n628), .A(n4882), .ZN(n4881) );
  NOR4_X1 U5145 ( .A1(n7285), .A2(n3998), .A3(n3999), .A4(n4000), .ZN(n3997)
         );
  XNOR2_X1 U5146 ( .A(n7258), .B(n2189), .ZN(n3998) );
  AOI222_X1 U5147 ( .A1(n883), .A2(n853), .B1(n838), .B2(HRDATA[13]), .C1(n839), .C2(vis_pc_o[12]), .ZN(n846) );
  NOR2_X1 U5148 ( .A1(n5063), .A2(n7518), .ZN(n3269) );
  NOR2_X1 U5149 ( .A1(n4123), .A2(n6592), .ZN(n1108) );
  NOR2_X1 U5150 ( .A1(n4123), .A2(n6597), .ZN(n1324) );
  NOR2_X1 U5151 ( .A1(n4123), .A2(n6910), .ZN(n1407) );
  AOI22_X1 U5152 ( .A1(n6245), .A2(n7617), .B1(n3036), .B2(n6775), .ZN(n6204)
         );
  AOI221_X1 U5153 ( .B1(n5345), .B2(n2189), .C1(n2857), .C2(n8291), .A(n5970), 
        .ZN(n5969) );
  OAI22_X1 U5154 ( .A1(n7562), .A2(n2197), .B1(n7611), .B2(n2195), .ZN(n5970)
         );
  AOI22_X1 U5155 ( .A1(n6137), .A2(n7555), .B1(n7554), .B2(n8156), .ZN(n6262)
         );
  AOI22_X1 U5156 ( .A1(n6362), .A2(n7565), .B1(n7566), .B2(n3024), .ZN(n6371)
         );
  OAI221_X1 U5157 ( .B1(n1809), .B2(n2513), .C1(n2569), .C2(n4548), .A(n452), 
        .ZN(n7827) );
  AOI221_X1 U5158 ( .B1(n934), .B2(n453), .C1(Zsfpw6[0]), .C2(n212), .A(n213), 
        .ZN(n452) );
  OAI222_X1 U5159 ( .A1(n2092), .A2(n6850), .B1(n735), .B2(n6830), .C1(n2086), 
        .C2(n7544), .ZN(n852) );
  NAND2_X1 U5160 ( .A1(n6021), .A2(n6022), .ZN(n5499) );
  AOI221_X1 U5161 ( .B1(vis_r2_o[28]), .B2(n561), .C1(vis_r0_o[28]), .C2(n547), 
        .A(n6024), .ZN(n6021) );
  AOI221_X1 U5162 ( .B1(vis_r3_o[28]), .B2(n567), .C1(vis_r7_o[28]), .C2(n5999), .A(n6023), .ZN(n6022) );
  OAI22_X1 U5163 ( .A1(n541), .A2(n8276), .B1(n540), .B2(n8264), .ZN(n6024) );
  OAI211_X1 U5164 ( .C1(n7574), .C2(n4729), .A(n2208), .B(n5292), .ZN(n853) );
  AOI222_X1 U5165 ( .A1(STCALIB[13]), .A2(n2973), .B1(n2975), .B2(n4161), .C1(
        n2976), .C2(Tzfpw6[13]), .ZN(n5292) );
  INV_X1 U5166 ( .A(n5295), .ZN(n2208) );
  AOI221_X1 U5167 ( .B1(n2988), .B2(n4470), .C1(n5345), .C2(n2500), .A(n5962), 
        .ZN(n5952) );
  OAI22_X1 U5168 ( .A1(n4788), .A2(n8356), .B1(n7614), .B2(n2195), .ZN(n5962)
         );
  AOI221_X1 U5169 ( .B1(n1124), .B2(n8224), .C1(n1125), .C2(K7hpw6[19]), .A(
        n1127), .ZN(n1116) );
  OAI22_X1 U5170 ( .A1(n8193), .A2(n2088), .B1(n8311), .B2(n2090), .ZN(n1127)
         );
  AOI221_X1 U5171 ( .B1(n839), .B2(vis_pc_o[30]), .C1(n883), .C2(n1110), .A(
        n1111), .ZN(n1102) );
  OAI22_X1 U5172 ( .A1(n8299), .A2(n2090), .B1(n6844), .B2(n2092), .ZN(n1111)
         );
  AOI221_X1 U5173 ( .B1(n839), .B2(vis_pc_o[29]), .C1(n883), .C2(n888), .A(
        n889), .ZN(n880) );
  OAI22_X1 U5174 ( .A1(n8300), .A2(n2090), .B1(n6855), .B2(n2092), .ZN(n889)
         );
  OAI221_X1 U5175 ( .B1(n2388), .B2(n3104), .C1(n865), .C2(n2712), .A(n4784), 
        .ZN(n4268) );
  AOI22_X1 U5176 ( .A1(n4717), .A2(n3312), .B1(HRDATA[17]), .B2(n4691), .ZN(
        n4784) );
  OAI222_X1 U5177 ( .A1(n2090), .A2(n8319), .B1(n2086), .B2(n7395), .C1(n2092), 
        .C2(n6749), .ZN(n1200) );
  OAI222_X1 U5178 ( .A1(n2090), .A2(n8326), .B1(n2086), .B2(n7547), .C1(n2092), 
        .C2(n6846), .ZN(n1295) );
  OAI222_X1 U5179 ( .A1(n2090), .A2(n8321), .B1(n2086), .B2(n7404), .C1(n2092), 
        .C2(n6699), .ZN(n1215) );
  OAI211_X1 U5180 ( .C1(n6381), .C2(n6382), .A(n8136), .B(n4001), .ZN(n6379)
         );
  NAND2_X1 U5181 ( .A1(n3276), .A2(n8134), .ZN(n6382) );
  AOI22_X1 U5182 ( .A1(n6383), .A2(n7568), .B1(n7567), .B2(n8236), .ZN(n6381)
         );
  AOI21_X1 U5183 ( .B1(n7569), .B2(n8248), .A(n7634), .ZN(n6383) );
  NAND4_X1 U5184 ( .A1(n2624), .A2(n5701), .A3(n5702), .A4(n5703), .ZN(n4939)
         );
  NAND2_X1 U5185 ( .A1(n4864), .A2(n8297), .ZN(n5701) );
  AOI222_X1 U5186 ( .A1(vis_r10_o[27]), .A2(n4861), .B1(vis_r11_o[27]), .B2(
        n615), .C1(vis_r9_o[27]), .C2(n4863), .ZN(n5702) );
  AOI221_X1 U5187 ( .B1(vis_r14_o[27]), .B2(n5272), .C1(vis_r8_o[27]), .C2(
        n4856), .A(n5704), .ZN(n5703) );
  OAI222_X1 U5188 ( .A1(n2088), .A2(n4806), .B1(n2092), .B2(n6757), .C1(n2090), 
        .C2(n8318), .ZN(n1193) );
  OAI222_X1 U5189 ( .A1(n2088), .A2(n4797), .B1(n2092), .B2(n6840), .C1(n2090), 
        .C2(n8304), .ZN(n1027) );
  OAI222_X1 U5190 ( .A1(n2086), .A2(n7333), .B1(n2094), .B2(n6791), .C1(n456), 
        .C2(n7484), .ZN(n1109) );
  OAI222_X1 U5191 ( .A1(n2086), .A2(n7658), .B1(n2094), .B2(n6802), .C1(n456), 
        .C2(n7474), .ZN(n887) );
  OAI222_X1 U5192 ( .A1(n2098), .A2(n7659), .B1(n741), .B2(n742), .C1(n881), 
        .C2(n7681), .ZN(n723) );
  OAI222_X1 U5193 ( .A1(n2098), .A2(n7413), .B1(n2088), .B2(n4799), .C1(n881), 
        .C2(n7693), .ZN(n1172) );
  NOR2_X1 U5194 ( .A1(n7433), .A2(n524), .ZN(n2375) );
  OAI21_X1 U5195 ( .B1(n489), .B2(n4377), .A(n7492), .ZN(n33) );
  NOR3_X1 U5196 ( .A1(n1926), .A2(n3628), .A3(n2251), .ZN(n4377) );
  NOR2_X1 U5197 ( .A1(n4123), .A2(n7479), .ZN(n1136) );
  OAI22_X1 U5198 ( .A1(n7558), .A2(n4285), .B1(n7557), .B2(n6130), .ZN(n6393)
         );
  NOR2_X1 U5199 ( .A1(n4123), .A2(n6572), .ZN(n1135) );
  OAI22_X1 U5200 ( .A1(n7564), .A2(n3869), .B1(n7563), .B2(n6276), .ZN(n6273)
         );
  AOI22_X1 U5201 ( .A1(n2185), .A2(n7626), .B1(n8175), .B2(n2339), .ZN(n5787)
         );
  NOR2_X1 U5202 ( .A1(n7582), .A2(n7598), .ZN(n6217) );
  NOR2_X1 U5203 ( .A1(n4112), .A2(n7481), .ZN(n1365) );
  OAI21_X1 U5204 ( .B1(n492), .B2(n7492), .A(n3760), .ZN(n5233) );
  AOI22_X1 U5205 ( .A1(n6362), .A2(n6772), .B1(n3024), .B2(n7670), .ZN(n6369)
         );
  AOI22_X1 U5206 ( .A1(n6130), .A2(n6758), .B1(n4285), .B2(n7678), .ZN(n6367)
         );
  AOI22_X1 U5207 ( .A1(n6379), .A2(n7568), .B1(n3274), .B2(n7634), .ZN(n6370)
         );
  AOI22_X1 U5208 ( .A1(n6131), .A2(n6700), .B1(n3643), .B2(n7639), .ZN(n6368)
         );
  OAI222_X1 U5209 ( .A1(n2140), .A2(n675), .B1(n7358), .B2(n676), .C1(n677), 
        .C2(n5112), .ZN(n7848) );
  OAI222_X1 U5211 ( .A1(n2139), .A2(n675), .B1(n7324), .B2(n676), .C1(n677), 
        .C2(n3968), .ZN(n7846) );
  AOI22_X1 U5212 ( .A1(n6135), .A2(n7552), .B1(n3668), .B2(n7636), .ZN(n6286)
         );
  AOI22_X1 U5213 ( .A1(n6276), .A2(n6774), .B1(n3869), .B2(n7676), .ZN(n6268)
         );
  OAI222_X1 U5214 ( .A1(n2145), .A2(n675), .B1(n7495), .B2(n676), .C1(n677), 
        .C2(n5126), .ZN(n7849) );
  OAI222_X1 U5215 ( .A1(n2142), .A2(n675), .B1(n7328), .B2(n676), .C1(n677), 
        .C2(n5111), .ZN(n7847) );
  INV_X1 U5216 ( .A(n402), .ZN(n2142) );
  OAI222_X1 U5217 ( .A1(n2146), .A2(n675), .B1(n7494), .B2(n676), .C1(n677), 
        .C2(n5105), .ZN(n7845) );
  INV_X1 U5218 ( .A(n386), .ZN(n2146) );
  OAI222_X1 U5219 ( .A1(n2143), .A2(n675), .B1(n7258), .B2(n676), .C1(n677), 
        .C2(n5088), .ZN(n7844) );
  INV_X1 U5220 ( .A(n393), .ZN(n2143) );
  AOI22_X1 U5221 ( .A1(n6137), .A2(n6759), .B1(n8156), .B2(n7675), .ZN(n6285)
         );
  OAI222_X1 U5222 ( .A1(n8324), .A2(n745), .B1(n7495), .B2(n746), .C1(n756), 
        .C2(n2163), .ZN(n7860) );
  OAI222_X1 U5223 ( .A1(n8325), .A2(n745), .B1(n7494), .B2(n746), .C1(n754), 
        .C2(n2163), .ZN(n7859) );
  OAI222_X1 U5224 ( .A1(n8327), .A2(n745), .B1(n7328), .B2(n746), .C1(n750), 
        .C2(n2163), .ZN(n7857) );
  OAI221_X1 U5225 ( .B1(n728), .B2(n6705), .C1(n2094), .C2(n6707), .A(n2076), 
        .ZN(n814) );
  INV_X1 U5226 ( .A(n816), .ZN(n2076) );
  OAI22_X1 U5227 ( .A1(n6703), .A2(n727), .B1(n6704), .B2(n2082), .ZN(n816) );
  OAI221_X1 U5228 ( .B1(n728), .B2(n6715), .C1(n2094), .C2(n6717), .A(n2037), 
        .ZN(n1045) );
  INV_X1 U5229 ( .A(n1047), .ZN(n2037) );
  OAI22_X1 U5230 ( .A1(n6713), .A2(n727), .B1(n6714), .B2(n2082), .ZN(n1047)
         );
  OAI221_X1 U5231 ( .B1(n728), .B2(n6738), .C1(n2094), .C2(n6740), .A(n2055), 
        .ZN(n896) );
  INV_X1 U5232 ( .A(n898), .ZN(n2055) );
  OAI22_X1 U5233 ( .A1(n6736), .A2(n727), .B1(n6737), .B2(n2082), .ZN(n898) );
  OAI221_X1 U5234 ( .B1(n728), .B2(n6815), .C1(n2094), .C2(n6798), .A(n2062), 
        .ZN(n871) );
  INV_X1 U5235 ( .A(n873), .ZN(n2062) );
  OAI22_X1 U5236 ( .A1(n6868), .A2(n727), .B1(n6892), .B2(n2082), .ZN(n873) );
  OAI221_X1 U5237 ( .B1(n728), .B2(n6805), .C1(n2094), .C2(n6786), .A(n2041), 
        .ZN(n1037) );
  INV_X1 U5238 ( .A(n1039), .ZN(n2041) );
  OAI22_X1 U5239 ( .A1(n6858), .A2(n727), .B1(n6878), .B2(n2082), .ZN(n1039)
         );
  OAI221_X1 U5240 ( .B1(n728), .B2(n6807), .C1(n2094), .C2(n6788), .A(n2069), 
        .ZN(n862) );
  INV_X1 U5241 ( .A(n864), .ZN(n2069) );
  OAI22_X1 U5242 ( .A1(n6860), .A2(n727), .B1(n6880), .B2(n2082), .ZN(n864) );
  OAI222_X1 U5243 ( .A1(n8328), .A2(n745), .B1(n7324), .B2(n746), .C1(n2211), 
        .C2(n2163), .ZN(n7856) );
  INV_X1 U5244 ( .A(HRDATA[1]), .ZN(n8328) );
  OAI222_X1 U5245 ( .A1(n8326), .A2(n745), .B1(n7258), .B2(n746), .C1(n752), 
        .C2(n2163), .ZN(n7858) );
  OAI222_X1 U5246 ( .A1(n8329), .A2(n745), .B1(n7358), .B2(n746), .C1(n795), 
        .C2(n2163), .ZN(n7869) );
  NAND2_X1 U5247 ( .A1(n6269), .A2(n6270), .ZN(n5306) );
  OAI21_X1 U5248 ( .B1(n7588), .B2(n7576), .A(n6275), .ZN(n6269) );
  OAI221_X1 U5249 ( .B1(n3296), .B2(n3868), .C1(n3866), .C2(n3869), .A(n6272), 
        .ZN(n6270) );
  INV_X1 U5250 ( .A(n6265), .ZN(n3296) );
  NAND4_X1 U5251 ( .A1(n5966), .A2(n5967), .A3(n5968), .A4(n5969), .ZN(n837)
         );
  AOI221_X1 U5252 ( .B1(n2985), .B2(n8242), .C1(n2884), .C2(n8244), .A(n5975), 
        .ZN(n5968) );
  AOI221_X1 U5253 ( .B1(n2866), .B2(n8250), .C1(n2852), .C2(n8240), .A(n5977), 
        .ZN(n5967) );
  AOI211_X1 U5254 ( .C1(STCALIB[15]), .C2(n2973), .A(n5979), .B(n4714), .ZN(
        n5966) );
  OAI22_X1 U5255 ( .A1(n683), .A2(n8079), .B1(n2269), .B2(n2362), .ZN(Ucrhu6)
         );
  OAI22_X1 U5256 ( .A1(n768), .A2(n8008), .B1(n2269), .B2(n2218), .ZN(Xarhu6)
         );
  OAI22_X1 U5257 ( .A1(n685), .A2(n6122), .B1(n2269), .B2(n2348), .ZN(Qarhu6)
         );
  OAI22_X1 U5258 ( .A1(n775), .A2(n5877), .B1(n2269), .B2(n771), .ZN(Jarhu6)
         );
  OAI22_X1 U5259 ( .A1(n686), .A2(n8222), .B1(n2276), .B2(n2348), .ZN(B6rhu6)
         );
  OAI22_X1 U5260 ( .A1(n683), .A2(n8220), .B1(n2276), .B2(n2362), .ZN(F8rhu6)
         );
  OAI22_X1 U5261 ( .A1(n767), .A2(n8218), .B1(n2276), .B2(n764), .ZN(I6rhu6)
         );
  OAI22_X1 U5262 ( .A1(n775), .A2(n8210), .B1(n2276), .B2(n2214), .ZN(U5rhu6)
         );
  OAI22_X1 U5263 ( .A1(n683), .A2(n8089), .B1(n2230), .B2(n681), .ZN(Muqhu6)
         );
  OAI22_X1 U5264 ( .A1(n683), .A2(n8084), .B1(n2343), .B2(n2362), .ZN(Q3rhu6)
         );
  OAI22_X1 U5265 ( .A1(n683), .A2(n8075), .B1(n2314), .B2(n2362), .ZN(Xpqhu6)
         );
  OAI22_X1 U5266 ( .A1(n768), .A2(n8059), .B1(n2230), .B2(n764), .ZN(Psqhu6)
         );
  OAI22_X1 U5267 ( .A1(n768), .A2(n8040), .B1(n2343), .B2(n2218), .ZN(T1rhu6)
         );
  OAI22_X1 U5268 ( .A1(n685), .A2(n6150), .B1(n2230), .B2(n684), .ZN(Isqhu6)
         );
  OAI22_X1 U5269 ( .A1(n686), .A2(n6136), .B1(n2343), .B2(n684), .ZN(M1rhu6)
         );
  OAI22_X1 U5270 ( .A1(n685), .A2(n6119), .B1(n2314), .B2(n2348), .ZN(Tnqhu6)
         );
  OAI22_X1 U5271 ( .A1(n775), .A2(n5897), .B1(n2230), .B2(n2214), .ZN(Bsqhu6)
         );
  OAI22_X1 U5272 ( .A1(n775), .A2(n5887), .B1(n2343), .B2(n2214), .ZN(F1rhu6)
         );
  OAI22_X1 U5273 ( .A1(n775), .A2(n5875), .B1(n2314), .B2(n771), .ZN(Mnqhu6)
         );
  OAI22_X1 U5274 ( .A1(n768), .A2(n4004), .B1(n2314), .B2(n2218), .ZN(Aoqhu6)
         );
  NOR3_X1 U5275 ( .A1(n3709), .A2(n7497), .A3(n4203), .ZN(n5234) );
  OAI221_X1 U5276 ( .B1(n6692), .B2(n2133), .C1(n220), .C2(n3871), .A(n240), 
        .ZN(n7747) );
  AOI22_X1 U5277 ( .A1(n241), .A2(\eq_3147/A[25] ), .B1(n1851), .B2(n8297), 
        .ZN(n240) );
  OAI221_X1 U5278 ( .B1(n7653), .B2(n2133), .C1(n220), .C2(n4797), .A(n248), 
        .ZN(n7750) );
  AOI22_X1 U5279 ( .A1(n241), .A2(\eq_3147/A[24] ), .B1(n1851), .B2(n8283), 
        .ZN(n248) );
  OAI221_X1 U5280 ( .B1(n6741), .B2(n2133), .C1(n220), .C2(n4766), .A(n278), 
        .ZN(n7762) );
  AOI22_X1 U5281 ( .A1(n241), .A2(\eq_3147/A[20] ), .B1(n1851), .B2(n8196), 
        .ZN(n278) );
  OAI221_X1 U5282 ( .B1(n6912), .B2(n2133), .C1(n220), .C2(n4765), .A(n271), 
        .ZN(n7759) );
  AOI22_X1 U5283 ( .A1(n241), .A2(\eq_3147/A[21] ), .B1(n1851), .B2(n8195), 
        .ZN(n271) );
  OAI221_X1 U5284 ( .B1(n6903), .B2(n2133), .C1(n220), .C2(n8174), .A(n299), 
        .ZN(n7774) );
  AOI22_X1 U5285 ( .A1(n241), .A2(\eq_3147/A[16] ), .B1(n1851), .B2(n8177), 
        .ZN(n299) );
  OAI221_X1 U5286 ( .B1(n6907), .B2(n2133), .C1(n220), .C2(n4772), .A(n284), 
        .ZN(n7765) );
  AOI22_X1 U5287 ( .A1(n241), .A2(\eq_3147/A[19] ), .B1(n1851), .B2(n3672), 
        .ZN(n284) );
  OAI221_X1 U5288 ( .B1(n6905), .B2(n2133), .C1(n220), .C2(n4773), .A(n304), 
        .ZN(n7777) );
  AOI22_X1 U5289 ( .A1(n241), .A2(\eq_3147/A[15] ), .B1(n1851), .B2(n3280), 
        .ZN(n304) );
  OAI22_X1 U5290 ( .A1(n2825), .A2(n2211), .B1(n4730), .B2(n7586), .ZN(n5295)
         );
  OAI22_X1 U5291 ( .A1(n3335), .A2(n2086), .B1(n6834), .B2(n735), .ZN(n1171)
         );
  OAI221_X1 U5292 ( .B1(n6904), .B2(n2133), .C1(n220), .C2(n8193), .A(n294), 
        .ZN(n7771) );
  AOI22_X1 U5293 ( .A1(n241), .A2(\eq_3147/A[17] ), .B1(n1851), .B2(n8224), 
        .ZN(n294) );
  OAI221_X1 U5294 ( .B1(n6718), .B2(n2133), .C1(n220), .C2(n4184), .A(n289), 
        .ZN(n7768) );
  AOI22_X1 U5295 ( .A1(n241), .A2(\eq_3147/A[18] ), .B1(n1851), .B2(n8223), 
        .ZN(n289) );
  OAI21_X1 U5296 ( .B1(n6106), .B2(n4673), .A(n7550), .ZN(n795) );
  AOI211_X1 U5297 ( .C1(n4789), .C2(n6107), .A(n5453), .B(n5297), .ZN(n6106)
         );
  OAI22_X1 U5298 ( .A1(n6109), .A2(n6110), .B1(n6111), .B2(n4790), .ZN(n6107)
         );
  AOI21_X1 U5299 ( .B1(n5314), .B2(n6112), .A(n6113), .ZN(n6111) );
  NAND3_X1 U5300 ( .A1(n808), .A2(n1663), .A3(n7497), .ZN(n4080) );
  OAI221_X1 U5301 ( .B1(n1580), .B2(n1849), .C1(n7344), .C2(n180), .A(n1846), 
        .ZN(n7744) );
  INV_X1 U5302 ( .A(n235), .ZN(n1846) );
  OAI222_X1 U5303 ( .A1(n1847), .A2(n8260), .B1(n2133), .B2(n6882), .C1(n220), 
        .C2(n4110), .ZN(n235) );
  OAI221_X1 U5304 ( .B1(n1606), .B2(n1849), .C1(n7706), .C2(n180), .A(n264), 
        .ZN(n7756) );
  AOI222_X1 U5305 ( .A1(vis_tbit_o), .A2(n182), .B1(n183), .B2(n3388), .C1(
        vis_pc_o[23]), .C2(n1852), .ZN(n264) );
  OAI221_X1 U5306 ( .B1(n1603), .B2(n1849), .C1(n3335), .C2(n180), .A(n255), 
        .ZN(n7753) );
  AOI221_X1 U5307 ( .B1(vis_pc_o[24]), .B2(n1852), .C1(n183), .C2(n3618), .A(
        n257), .ZN(n255) );
  AND4_X1 U5308 ( .A1(n180), .A2(n258), .A3(n259), .A4(vis_control_o), .ZN(
        n257) );
  OAI221_X1 U5309 ( .B1(n3503), .B2(n2167), .C1(n7531), .C2(n798), .A(n792), 
        .ZN(Wfphu6) );
  NOR3_X1 U5310 ( .A1(n5401), .A2(n5402), .A3(n2869), .ZN(n874) );
  OAI21_X1 U5311 ( .B1(n1894), .B2(n7702), .A(n903), .ZN(n5402) );
  INV_X1 U5312 ( .A(n5404), .ZN(n2869) );
  OAI22_X1 U5313 ( .A1(n754), .A2(n2825), .B1(n4723), .B2(n6634), .ZN(n5401)
         );
  OAI22_X1 U5314 ( .A1(n7628), .A2(n2706), .B1(n2707), .B2(n3733), .ZN(Ruphu6)
         );
  INV_X1 U5315 ( .A(n2706), .ZN(n3733) );
  AOI211_X1 U5316 ( .C1(n504), .C2(n3805), .A(n3749), .B(n961), .ZN(n2706) );
  AOI22_X1 U5317 ( .A1(n358), .A2(n810), .B1(n3765), .B2(n2709), .ZN(n2707) );
  AND2_X1 U5318 ( .A1(Ntkbx6[19]), .A2(n4277), .ZN(Clihu6) );
  OAI22_X1 U5319 ( .A1(n701), .A2(n1639), .B1(n2297), .B2(n8193), .ZN(n4277)
         );
  AND2_X1 U5320 ( .A1(Ntkbx6[13]), .A2(n3969), .ZN(Gdihu6) );
  OAI22_X1 U5321 ( .A1(n697), .A2(n1709), .B1(n2297), .B2(n4802), .ZN(n3969)
         );
  AND2_X1 U5322 ( .A1(Ntkbx6[12]), .A2(n2329), .ZN(Ybihu6) );
  OAI22_X1 U5323 ( .A1(n701), .A2(n1718), .B1(n2297), .B2(n4805), .ZN(n2329)
         );
  AND2_X1 U5324 ( .A1(Ntkbx6[20]), .A2(n3452), .ZN(Kmihu6) );
  OAI22_X1 U5325 ( .A1(n697), .A2(n1633), .B1(n696), .B2(n4184), .ZN(n3452) );
  AND2_X1 U5326 ( .A1(Ntkbx6[17]), .A2(n3100), .ZN(Miihu6) );
  OAI22_X1 U5327 ( .A1(n697), .A2(n1656), .B1(n696), .B2(n4773), .ZN(n3100) );
  AND2_X1 U5328 ( .A1(Ntkbx6[14]), .A2(n3005), .ZN(Oeihu6) );
  OAI22_X1 U5329 ( .A1(n701), .A2(n1693), .B1(n696), .B2(n4801), .ZN(n3005) );
  AND2_X1 U5330 ( .A1(Ntkbx6[11]), .A2(n2791), .ZN(Qaihu6) );
  OAI22_X1 U5331 ( .A1(n701), .A2(n1738), .B1(n696), .B2(n4806), .ZN(n2791) );
  AND2_X1 U5332 ( .A1(Ntkbx6[10]), .A2(n3834), .ZN(I9ihu6) );
  OAI22_X1 U5333 ( .A1(n701), .A2(n1766), .B1(n696), .B2(n4807), .ZN(n3834) );
  AND2_X1 U5334 ( .A1(Ntkbx6[9]), .A2(n5412), .ZN(A8ihu6) );
  OAI22_X1 U5335 ( .A1(n701), .A2(n1769), .B1(n696), .B2(n4777), .ZN(n5412) );
  AND2_X1 U5336 ( .A1(Ntkbx6[15]), .A2(n2431), .ZN(Wfihu6) );
  OAI22_X1 U5337 ( .A1(n701), .A2(n1681), .B1(n2297), .B2(n4776), .ZN(n2431)
         );
  NAND4_X1 U5338 ( .A1(n3522), .A2(n3729), .A3(n4366), .A4(n4367), .ZN(n4363)
         );
  NAND4_X1 U5339 ( .A1(n4374), .A2(n476), .A3(n7399), .A4(n4375), .ZN(n4366)
         );
  AOI21_X1 U5340 ( .B1(n1749), .B2(n228), .A(n4368), .ZN(n4367) );
  OAI21_X1 U5341 ( .B1(n7514), .B2(n1493), .A(n4587), .ZN(n4374) );
  AND2_X1 U5342 ( .A1(Ntkbx6[21]), .A2(n2673), .ZN(Snihu6) );
  OAI22_X1 U5343 ( .A1(n697), .A2(n1631), .B1(n696), .B2(n4772), .ZN(n2673) );
  AND2_X1 U5344 ( .A1(Ntkbx6[18]), .A2(n2540), .ZN(Ujihu6) );
  OAI22_X1 U5345 ( .A1(n697), .A2(n1652), .B1(n696), .B2(n8174), .ZN(n2540) );
  AND2_X1 U5346 ( .A1(Nvkbx6[10]), .A2(n2417), .ZN(Wskhu6) );
  OAI22_X1 U5347 ( .A1(n733), .A2(n4807), .B1(n736), .B2(n1766), .ZN(n2417) );
  NAND2_X1 U5348 ( .A1(n6034), .A2(n6035), .ZN(n5286) );
  AOI221_X1 U5349 ( .B1(vis_r2_o[31]), .B2(n6003), .C1(vis_r0_o[31]), .C2(n547), .A(n6037), .ZN(n6034) );
  AOI221_X1 U5350 ( .B1(vis_r3_o[31]), .B2(n567), .C1(vis_r7_o[31]), .C2(n5999), .A(n6036), .ZN(n6035) );
  OAI22_X1 U5351 ( .A1(n6006), .A2(n6577), .B1(n6007), .B2(n5319), .ZN(n6037)
         );
  NAND2_X1 U5352 ( .A1(n6025), .A2(n6026), .ZN(n5498) );
  AOI221_X1 U5353 ( .B1(vis_r2_o[29]), .B2(n561), .C1(vis_r0_o[29]), .C2(n547), 
        .A(n6028), .ZN(n6025) );
  AOI221_X1 U5354 ( .B1(vis_r3_o[29]), .B2(n5998), .C1(vis_r7_o[29]), .C2(
        n5999), .A(n6027), .ZN(n6026) );
  OAI22_X1 U5355 ( .A1(n6006), .A2(n6590), .B1(n6007), .B2(n5333), .ZN(n6028)
         );
  NAND2_X1 U5356 ( .A1(n6029), .A2(n6030), .ZN(n5489) );
  AOI221_X1 U5357 ( .B1(vis_r2_o[30]), .B2(n561), .C1(vis_r0_o[30]), .C2(n547), 
        .A(n6032), .ZN(n6029) );
  AOI221_X1 U5358 ( .B1(vis_r3_o[30]), .B2(n5998), .C1(vis_r7_o[30]), .C2(
        n5999), .A(n6031), .ZN(n6030) );
  OAI22_X1 U5359 ( .A1(n6006), .A2(n6486), .B1(n6007), .B2(n5433), .ZN(n6032)
         );
  XNOR2_X1 U5360 ( .A(n7324), .B(n2211), .ZN(n3996) );
  AND2_X1 U5361 ( .A1(Nvkbx6[18]), .A2(n3839), .ZN(I3lhu6) );
  OAI22_X1 U5362 ( .A1(n733), .A2(n8174), .B1(n736), .B2(n1652), .ZN(n3839) );
  AND2_X1 U5363 ( .A1(Nvkbx6[17]), .A2(n5623), .ZN(A2lhu6) );
  OAI22_X1 U5364 ( .A1(n733), .A2(n4773), .B1(n736), .B2(n1656), .ZN(n5623) );
  AND2_X1 U5365 ( .A1(Nvkbx6[16]), .A2(n2701), .ZN(S0lhu6) );
  OAI22_X1 U5366 ( .A1(n2264), .A2(n4774), .B1(n736), .B2(n1671), .ZN(n2701)
         );
  AND2_X1 U5367 ( .A1(Nvkbx6[14]), .A2(n4200), .ZN(Cykhu6) );
  OAI22_X1 U5368 ( .A1(n733), .A2(n4801), .B1(n734), .B2(n1693), .ZN(n4200) );
  AND2_X1 U5369 ( .A1(Nvkbx6[12]), .A2(n3079), .ZN(Mvkhu6) );
  OAI22_X1 U5370 ( .A1(n2264), .A2(n4805), .B1(n736), .B2(n1718), .ZN(n3079)
         );
  AND2_X1 U5371 ( .A1(Nvkbx6[19]), .A2(n2810), .ZN(Q4lhu6) );
  OAI22_X1 U5372 ( .A1(n2264), .A2(n8193), .B1(n736), .B2(n1639), .ZN(n2810)
         );
  AND2_X1 U5373 ( .A1(Nvkbx6[13]), .A2(n2518), .ZN(Uwkhu6) );
  OAI22_X1 U5375 ( .A1(n2264), .A2(n4802), .B1(n734), .B2(n1709), .ZN(n2518)
         );
  AND2_X1 U5376 ( .A1(Nvkbx6[15]), .A2(n3291), .ZN(Kzkhu6) );
  OAI22_X1 U5377 ( .A1(n2264), .A2(n4776), .B1(n736), .B2(n1681), .ZN(n3291)
         );
  AND2_X1 U5378 ( .A1(Nvkbx6[9]), .A2(n2971), .ZN(Orkhu6) );
  OAI22_X1 U5379 ( .A1(n2264), .A2(n4777), .B1(n736), .B2(n1769), .ZN(n2971)
         );
  OAI211_X1 U5380 ( .C1(n6278), .C2(n6277), .A(n4061), .B(n8141), .ZN(n6276)
         );
  AOI22_X1 U5381 ( .A1(n6279), .A2(n6774), .B1(n7564), .B2(n4474), .ZN(n6278)
         );
  AOI21_X1 U5382 ( .B1(n7563), .B2(n4478), .A(n7676), .ZN(n6279) );
  OAI22_X1 U5383 ( .A1(n682), .A2(n8194), .B1(n2209), .B2(n681), .ZN(Bzqhu6)
         );
  OAI22_X1 U5384 ( .A1(n767), .A2(n8191), .B1(n2209), .B2(n2218), .ZN(Exqhu6)
         );
  OAI22_X1 U5385 ( .A1(n686), .A2(n6175), .B1(n2288), .B2(n684), .ZN(Cushu6)
         );
  OAI22_X1 U5386 ( .A1(n686), .A2(n6168), .B1(n2248), .B2(n2348), .ZN(Ejqhu6)
         );
  OAI22_X1 U5387 ( .A1(n775), .A2(n8183), .B1(n2209), .B2(n771), .ZN(Qwqhu6)
         );
  OAI22_X1 U5388 ( .A1(n686), .A2(n8179), .B1(n2209), .B2(n2348), .ZN(Xwqhu6)
         );
  OAI22_X1 U5389 ( .A1(n683), .A2(n8090), .B1(n2299), .B2(n681), .ZN(Msshu6)
         );
  OAI22_X1 U5390 ( .A1(n768), .A2(n8060), .B1(n2299), .B2(n764), .ZN(Pqshu6)
         );
  OAI22_X1 U5391 ( .A1(n686), .A2(n6151), .B1(n2299), .B2(n684), .ZN(Iqshu6)
         );
  OAI22_X1 U5392 ( .A1(n772), .A2(n5865), .B1(n2299), .B2(n771), .ZN(Otshu6)
         );
  OAI22_X1 U5393 ( .A1(n683), .A2(n8096), .B1(n2248), .B2(n681), .ZN(Ilqhu6)
         );
  OAI22_X1 U5394 ( .A1(n768), .A2(n8065), .B1(n2248), .B2(n764), .ZN(Ljqhu6)
         );
  OAI22_X1 U5395 ( .A1(n772), .A2(n5825), .B1(n2248), .B2(n2214), .ZN(Xiqhu6)
         );
  OAI22_X1 U5396 ( .A1(n682), .A2(n8094), .B1(n2325), .B2(n681), .ZN(Jhrhu6)
         );
  OAI22_X1 U5397 ( .A1(n682), .A2(n8081), .B1(n2318), .B2(n2362), .ZN(Qnshu6)
         );
  OAI22_X1 U5398 ( .A1(n767), .A2(n8064), .B1(n2325), .B2(n764), .ZN(Mfrhu6)
         );
  OAI22_X1 U5399 ( .A1(n767), .A2(n8036), .B1(n2318), .B2(n764), .ZN(Tlshu6)
         );
  OAI22_X1 U5400 ( .A1(n685), .A2(n6156), .B1(n2325), .B2(n684), .ZN(Ffrhu6)
         );
  OAI22_X1 U5401 ( .A1(n685), .A2(n6128), .B1(n2318), .B2(n684), .ZN(Mlshu6)
         );
  OAI22_X1 U5402 ( .A1(n685), .A2(n6121), .B1(n2236), .B2(n684), .ZN(Qorhu6)
         );
  OAI22_X1 U5403 ( .A1(n772), .A2(n5876), .B1(n2236), .B2(n2214), .ZN(Jorhu6)
         );
  OAI22_X1 U5404 ( .A1(n775), .A2(n5851), .B1(n2288), .B2(n2214), .ZN(Prrhu6)
         );
  OAI22_X1 U5405 ( .A1(n775), .A2(n5846), .B1(n2318), .B2(n771), .ZN(Soshu6)
         );
  OAI22_X1 U5406 ( .A1(n775), .A2(n5822), .B1(n2325), .B2(n2214), .ZN(Yerhu6)
         );
  NAND4_X1 U5407 ( .A1(n1101), .A2(n1102), .A3(n2022), .A4(n1104), .ZN(n7898)
         );
  AOI221_X1 U5408 ( .B1(n239), .B2(n3880), .C1(n856), .C2(n3877), .A(n858), 
        .ZN(n1101) );
  AOI221_X1 U5409 ( .B1(ECOREVNUM[23]), .B2(n2002), .C1(n884), .C2(n4336), .A(
        n1106), .ZN(n1104) );
  INV_X1 U5410 ( .A(n1109), .ZN(n2022) );
  NAND4_X1 U5411 ( .A1(n879), .A2(n880), .A3(n2024), .A4(n882), .ZN(n7878) );
  AOI221_X1 U5412 ( .B1(n239), .B2(n4151), .C1(n856), .C2(n3125), .A(n858), 
        .ZN(n879) );
  AOI221_X1 U5413 ( .B1(ECOREVNUM[22]), .B2(n2002), .C1(n884), .C2(n4335), .A(
        n886), .ZN(n882) );
  INV_X1 U5414 ( .A(n887), .ZN(n2024) );
  NAND4_X1 U5415 ( .A1(n1076), .A2(n1077), .A3(n2084), .A4(n1079), .ZN(n7896)
         );
  AOI21_X1 U5416 ( .B1(n856), .B2(n8205), .A(n858), .ZN(n1076) );
  AOI222_X1 U5417 ( .A1(n1080), .A2(E1hpw6[29]), .B1(n883), .B2(n1082), .C1(
        ECOREVNUM[21]), .C2(n2002), .ZN(n1079) );
  AOI222_X1 U5418 ( .A1(n239), .A2(n8206), .B1(n838), .B2(HRDATA[29]), .C1(
        n839), .C2(vis_pc_o[28]), .ZN(n1077) );
  OAI21_X1 U5419 ( .B1(n6685), .B2(N701), .A(n2064), .ZN(n6917) );
  NAND3_X1 U5420 ( .A1(n2065), .A2(N701), .A3(n2066), .ZN(n2064) );
  AOI221_X1 U5421 ( .B1(n2067), .B2(n2068), .C1(n1957), .C2(n4674), .A(n1144), 
        .ZN(n2066) );
  OR2_X1 U5422 ( .A1(n2073), .A2(n1960), .ZN(n2068) );
  INV_X1 U5423 ( .A(n5296), .ZN(n2211) );
  OAI211_X1 U5424 ( .C1(n5297), .C2(n5298), .A(n7705), .B(n7550), .ZN(n5296)
         );
  AOI221_X1 U5425 ( .B1(n2783), .B2(n5300), .C1(n5301), .C2(n4790), .A(n2212), 
        .ZN(n5298) );
  OAI22_X1 U5426 ( .A1(n3638), .A2(n3014), .B1(n5314), .B2(n5315), .ZN(n5300)
         );
  NAND4_X1 U5427 ( .A1(n2003), .A2(n1160), .A3(n2028), .A4(n1162), .ZN(n7902)
         );
  AOI221_X1 U5428 ( .B1(n876), .B2(n8176), .C1(n883), .C2(n1164), .A(n1165), 
        .ZN(n1162) );
  INV_X1 U5429 ( .A(n1172), .ZN(n2003) );
  AOI221_X1 U5430 ( .B1(n1125), .B2(K7hpw6[25]), .C1(n838), .C2(HRDATA[25]), 
        .A(n1171), .ZN(n1160) );
  OAI21_X1 U5431 ( .B1(n6682), .B2(N701), .A(n2169), .ZN(n7256) );
  OAI21_X1 U5432 ( .B1(n2170), .B2(n2171), .A(N701), .ZN(n2169) );
  NAND2_X1 U5433 ( .A1(n806), .A2(n3993), .ZN(n793) );
  NAND4_X1 U5434 ( .A1(n3994), .A2(n3995), .A3(n3996), .A4(n3997), .ZN(n3993)
         );
  XNOR2_X1 U5435 ( .A(n7328), .B(n750), .ZN(n3994) );
  XNOR2_X1 U5436 ( .A(n2232), .B(n2181), .ZN(n3995) );
  OAI211_X1 U5437 ( .C1(n7682), .C2(n798), .A(n2319), .B(n792), .ZN(Yhvhu6) );
  NAND3_X1 U5438 ( .A1(HRDATA[15]), .A2(n798), .A3(n3503), .ZN(n2319) );
  OAI211_X1 U5439 ( .C1(n8317), .C2(n745), .A(n785), .B(n786), .ZN(n7867) );
  NAND2_X1 U5440 ( .A1(Xlfpw6[7]), .A2(n763), .ZN(n785) );
  AOI22_X1 U5441 ( .A1(n2167), .A2(n3546), .B1(IRQLATENCY[6]), .B2(n2164), 
        .ZN(n786) );
  OAI211_X1 U5442 ( .C1(n8318), .C2(n745), .A(n781), .B(n782), .ZN(n7866) );
  NAND2_X1 U5443 ( .A1(Xlfpw6[6]), .A2(n763), .ZN(n781) );
  AOI22_X1 U5444 ( .A1(n2167), .A2(n3545), .B1(IRQLATENCY[5]), .B2(n2164), 
        .ZN(n782) );
  OAI211_X1 U5445 ( .C1(n8319), .C2(n745), .A(n777), .B(n778), .ZN(n7865) );
  NAND2_X1 U5446 ( .A1(Xlfpw6[5]), .A2(n763), .ZN(n777) );
  AOI22_X1 U5447 ( .A1(n2167), .A2(n3544), .B1(IRQLATENCY[4]), .B2(n2164), 
        .ZN(n778) );
  OAI211_X1 U5448 ( .C1(n8320), .C2(n745), .A(n773), .B(n774), .ZN(n7864) );
  NAND2_X1 U5449 ( .A1(Xlfpw6[4]), .A2(n763), .ZN(n773) );
  AOI22_X1 U5450 ( .A1(n2167), .A2(n3543), .B1(IRQLATENCY[3]), .B2(n2164), 
        .ZN(n774) );
  OAI211_X1 U5451 ( .C1(n8321), .C2(n745), .A(n769), .B(n770), .ZN(n7863) );
  NAND2_X1 U5452 ( .A1(Xlfpw6[3]), .A2(n763), .ZN(n769) );
  AOI22_X1 U5453 ( .A1(n2167), .A2(n3540), .B1(IRQLATENCY[2]), .B2(n2164), 
        .ZN(n770) );
  OAI211_X1 U5454 ( .C1(n8322), .C2(n745), .A(n765), .B(n766), .ZN(n7862) );
  INV_X1 U5455 ( .A(HRDATA[7]), .ZN(n8322) );
  NAND2_X1 U5456 ( .A1(Xlfpw6[2]), .A2(n763), .ZN(n765) );
  AOI22_X1 U5457 ( .A1(n2167), .A2(n3538), .B1(IRQLATENCY[1]), .B2(n2164), 
        .ZN(n766) );
  OAI211_X1 U5458 ( .C1(n8323), .C2(n745), .A(n758), .B(n759), .ZN(n7861) );
  INV_X1 U5459 ( .A(HRDATA[6]), .ZN(n8323) );
  NAND2_X1 U5460 ( .A1(Xlfpw6[1]), .A2(n763), .ZN(n758) );
  AOI22_X1 U5461 ( .A1(n2167), .A2(n3535), .B1(IRQLATENCY[0]), .B2(n2164), 
        .ZN(n759) );
  OAI211_X1 U5462 ( .C1(n8316), .C2(n745), .A(n789), .B(n790), .ZN(n7868) );
  NAND2_X1 U5463 ( .A1(Xlfpw6[8]), .A2(n763), .ZN(n789) );
  AOI22_X1 U5464 ( .A1(n2167), .A2(n3534), .B1(IRQLATENCY[7]), .B2(n2164), 
        .ZN(n790) );
  INV_X1 U5465 ( .A(STCALIB[25]), .ZN(n8356) );
  OR4_X1 U5466 ( .A1(n811), .A2(n812), .A3(n813), .A4(n814), .ZN(n7872) );
  OAI221_X1 U5467 ( .B1(n881), .B2(n7641), .C1(n2098), .C2(n6667), .A(n819), 
        .ZN(n811) );
  OAI222_X1 U5468 ( .A1(n2092), .A2(n6709), .B1(n735), .B2(n6706), .C1(n2086), 
        .C2(n7446), .ZN(n813) );
  OAI222_X1 U5469 ( .A1(n741), .A2(n817), .B1(n2090), .B2(n8315), .C1(n2088), 
        .C2(n4801), .ZN(n812) );
  OR4_X1 U5471 ( .A1(n1042), .A2(n1043), .A3(n1044), .A4(n1045), .ZN(n7894) );
  OAI221_X1 U5472 ( .B1(n881), .B2(n7661), .C1(n2098), .C2(n7662), .A(n901), 
        .ZN(n1042) );
  OAI222_X1 U5473 ( .A1(n741), .A2(n2840), .B1(n2090), .B2(n8310), .C1(n2088), 
        .C2(n4184), .ZN(n1043) );
  OAI222_X1 U5474 ( .A1(n2092), .A2(n6719), .B1(n456), .B2(n6716), .C1(n2086), 
        .C2(n7660), .ZN(n1044) );
  OR4_X1 U5475 ( .A1(n893), .A2(n2012), .A3(n895), .A4(n896), .ZN(n7879) );
  OAI221_X1 U5476 ( .B1(n881), .B2(n7667), .C1(n2098), .C2(n6662), .A(n901), 
        .ZN(n893) );
  INV_X1 U5477 ( .A(n899), .ZN(n2012) );
  OAI222_X1 U5478 ( .A1(n2092), .A2(n6742), .B1(n456), .B2(n6739), .C1(n2086), 
        .C2(n7666), .ZN(n895) );
  OR4_X1 U5479 ( .A1(n829), .A2(n2009), .A3(n831), .A4(n832), .ZN(n7874) );
  OAI221_X1 U5480 ( .B1(n881), .B2(n7437), .C1(n2098), .C2(n6666), .A(n819), 
        .ZN(n829) );
  OAI222_X1 U5481 ( .A1(n2092), .A2(n6767), .B1(n456), .B2(n6764), .C1(n2086), 
        .C2(n7436), .ZN(n831) );
  OAI221_X1 U5482 ( .B1(n728), .B2(n6763), .C1(n2094), .C2(n6765), .A(n2075), 
        .ZN(n832) );
  OR4_X1 U5483 ( .A1(n868), .A2(n869), .A3(n870), .A4(n871), .ZN(n7877) );
  OAI221_X1 U5484 ( .B1(n881), .B2(n7387), .C1(n2098), .C2(n7386), .A(n867), 
        .ZN(n868) );
  OAI222_X1 U5485 ( .A1(n741), .A2(n874), .B1(n2090), .B2(n8314), .C1(n2088), 
        .C2(n4774), .ZN(n869) );
  OAI222_X1 U5486 ( .A1(n2092), .A2(n6851), .B1(n735), .B2(n6831), .C1(n2086), 
        .C2(n7385), .ZN(n870) );
  OR4_X1 U5487 ( .A1(n1034), .A2(n1035), .A3(n1036), .A4(n1037), .ZN(n7893) );
  OAI221_X1 U5488 ( .B1(n881), .B2(n7664), .C1(n2098), .C2(n7665), .A(n901), 
        .ZN(n1034) );
  OAI222_X1 U5489 ( .A1(n741), .A2(n2833), .B1(n2090), .B2(n8309), .C1(n2088), 
        .C2(n4772), .ZN(n1035) );
  OAI222_X1 U5490 ( .A1(n2092), .A2(n6839), .B1(n735), .B2(n6821), .C1(n2086), 
        .C2(n7663), .ZN(n1036) );
  OR4_X1 U5491 ( .A1(n859), .A2(n860), .A3(n861), .A4(n862), .ZN(n7876) );
  OAI221_X1 U5492 ( .B1(n881), .B2(n7648), .C1(n2098), .C2(n6664), .A(n867), 
        .ZN(n859) );
  OAI222_X1 U5493 ( .A1(n2092), .A2(n6841), .B1(n456), .B2(n6823), .C1(n2086), 
        .C2(n7647), .ZN(n861) );
  OAI222_X1 U5494 ( .A1(n741), .A2(n865), .B1(n2090), .B2(n8313), .C1(n2088), 
        .C2(n4773), .ZN(n860) );
  OR4_X1 U5495 ( .A1(n1151), .A2(n1152), .A3(n1153), .A4(n1154), .ZN(n7901) );
  OAI222_X1 U5496 ( .A1(n2098), .A2(n7650), .B1(n741), .B2(n1158), .C1(n881), 
        .C2(n7657), .ZN(n1151) );
  OAI222_X1 U5497 ( .A1(n2086), .A2(n7649), .B1(n2094), .B2(n6691), .C1(n735), 
        .C2(n6690), .ZN(n1153) );
  OAI222_X1 U5498 ( .A1(n2088), .A2(n3871), .B1(n2092), .B2(n6693), .C1(n2090), 
        .C2(n8303), .ZN(n1152) );
  OR4_X1 U5499 ( .A1(n723), .A2(n724), .A3(n725), .A4(n726), .ZN(n7855) );
  OAI222_X1 U5500 ( .A1(n2086), .A2(n7680), .B1(n2094), .B2(n6733), .C1(n456), 
        .C2(n6732), .ZN(n725) );
  OAI222_X1 U5501 ( .A1(n2088), .A2(n4765), .B1(n2092), .B2(n6734), .C1(n2090), 
        .C2(n8307), .ZN(n724) );
  OAI221_X1 U5502 ( .B1(n727), .B2(n6729), .C1(n728), .C2(n6731), .A(n2018), 
        .ZN(n726) );
  OR4_X1 U5503 ( .A1(n1199), .A2(n1200), .A3(n1201), .A4(n1202), .ZN(n7905) );
  OAI222_X1 U5504 ( .A1(n456), .A2(n6747), .B1(n728), .B2(n6746), .C1(n2094), 
        .C2(n6748), .ZN(n1201) );
  OAI222_X1 U5505 ( .A1(n2098), .A2(n7396), .B1(n2088), .B2(n4807), .C1(n881), 
        .C2(n7397), .ZN(n1199) );
  OAI221_X1 U5506 ( .B1(n2082), .B2(n6745), .C1(n727), .C2(n6744), .A(n1203), 
        .ZN(n1202) );
  OR4_X1 U5507 ( .A1(n1192), .A2(n1193), .A3(n1194), .A4(n1195), .ZN(n7904) );
  OAI222_X1 U5508 ( .A1(n2098), .A2(n6652), .B1(n741), .B2(n2835), .C1(n881), 
        .C2(n7631), .ZN(n1192) );
  OAI221_X1 U5509 ( .B1(n727), .B2(n6751), .C1(n728), .C2(n6753), .A(n1196), 
        .ZN(n1195) );
  OAI222_X1 U5510 ( .A1(n2086), .A2(n7630), .B1(n2094), .B2(n6755), .C1(n456), 
        .C2(n6754), .ZN(n1194) );
  OR4_X1 U5511 ( .A1(n820), .A2(n821), .A3(n822), .A4(n823), .ZN(n7873) );
  OAI221_X1 U5512 ( .B1(n881), .B2(n7450), .C1(n2098), .C2(n7449), .A(n819), 
        .ZN(n820) );
  OAI222_X1 U5513 ( .A1(n2086), .A2(n7629), .B1(n2094), .B2(n6796), .C1(n735), 
        .C2(n6829), .ZN(n822) );
  OAI222_X1 U5515 ( .A1(n2088), .A2(n4805), .B1(n2092), .B2(n6849), .C1(n2090), 
        .C2(n8317), .ZN(n821) );
  OR4_X1 U5516 ( .A1(n1294), .A2(n1295), .A3(n1296), .A4(n1297), .ZN(n7911) );
  OAI222_X1 U5517 ( .A1(n456), .A2(n1397), .B1(n728), .B2(n1515), .C1(n2094), 
        .C2(n6793), .ZN(n1296) );
  OAI222_X1 U5518 ( .A1(n4048), .A2(n2098), .B1(n2088), .B2(n4787), .C1(n881), 
        .C2(n7418), .ZN(n1294) );
  OAI221_X1 U5519 ( .B1(n2082), .B2(n1256), .C1(n727), .C2(n1119), .A(n1298), 
        .ZN(n1297) );
  OR4_X1 U5520 ( .A1(n1214), .A2(n1215), .A3(n1216), .A4(n1217), .ZN(n7907) );
  OAI222_X1 U5521 ( .A1(n735), .A2(n6697), .B1(n728), .B2(n6696), .C1(n2094), 
        .C2(n6698), .ZN(n1216) );
  OAI222_X1 U5522 ( .A1(n2098), .A2(n7405), .B1(n2088), .B2(n4810), .C1(n881), 
        .C2(n7406), .ZN(n1214) );
  OAI221_X1 U5523 ( .B1(n2082), .B2(n6695), .C1(n727), .C2(n6694), .A(n1218), 
        .ZN(n1217) );
  OR4_X1 U5524 ( .A1(n1206), .A2(n1207), .A3(n1208), .A4(n1209), .ZN(n7906) );
  OAI222_X1 U5525 ( .A1(n2098), .A2(n6651), .B1(n741), .B2(n2828), .C1(n881), 
        .C2(n7407), .ZN(n1206) );
  OAI222_X1 U5526 ( .A1(n2086), .A2(n7408), .B1(n2094), .B2(n6785), .C1(n735), 
        .C2(n6820), .ZN(n1208) );
  OAI222_X1 U5527 ( .A1(n2088), .A2(n4777), .B1(n2092), .B2(n6838), .C1(n2090), 
        .C2(n8320), .ZN(n1207) );
  OR4_X1 U5528 ( .A1(n1026), .A2(n1027), .A3(n1028), .A4(n1029), .ZN(n7892) );
  OAI221_X1 U5529 ( .B1(n881), .B2(n7655), .C1(n2098), .C2(n6658), .A(n901), 
        .ZN(n1026) );
  OAI221_X1 U5530 ( .B1(n727), .B2(n6859), .C1(n728), .C2(n6806), .A(n1030), 
        .ZN(n1029) );
  OAI222_X1 U5531 ( .A1(n2086), .A2(n7654), .B1(n2094), .B2(n6787), .C1(n735), 
        .C2(n6822), .ZN(n1028) );
  INV_X1 U5532 ( .A(n6101), .ZN(n2176) );
  OAI211_X1 U5533 ( .C1(n6629), .C2(n4729), .A(n6102), .B(n6103), .ZN(n6101)
         );
  AOI222_X1 U5534 ( .A1(STCALIB[12]), .A2(n2973), .B1(n2975), .B2(n8104), .C1(
        n2976), .C2(Tzfpw6[12]), .ZN(n6103) );
  AOI22_X1 U5535 ( .A1(n2181), .A2(n5345), .B1(n2866), .B2(n8106), .ZN(n6102)
         );
  AND4_X1 U5536 ( .A1(n5446), .A2(n5447), .A3(n5448), .A4(n2191), .ZN(n817) );
  AOI221_X1 U5537 ( .B1(n2886), .B2(n8254), .C1(n2882), .C2(n8256), .A(n5466), 
        .ZN(n5448) );
  AOI221_X1 U5538 ( .B1(n2978), .B2(n8255), .C1(n2866), .C2(n8259), .A(n5469), 
        .ZN(n5447) );
  AOI221_X1 U5539 ( .B1(n2976), .B2(Tzfpw6[14]), .C1(STCALIB[14]), .C2(n2973), 
        .A(n4714), .ZN(n5446) );
  INV_X1 U5540 ( .A(n6274), .ZN(n3293) );
  AOI22_X1 U5541 ( .A1(n6275), .A2(n7561), .B1(n3300), .B2(n6773), .ZN(n6274)
         );
  INV_X1 U5542 ( .A(n835), .ZN(n2009) );
  AOI222_X1 U5543 ( .A1(n883), .A2(n837), .B1(n838), .B2(HRDATA[15]), .C1(n839), .C2(vis_pc_o[14]), .ZN(n835) );
  OR3_X1 U5544 ( .A1(n1318), .A2(n1319), .A3(n1320), .ZN(n7912) );
  OAI22_X1 U5545 ( .A1(n728), .A2(n1516), .B1(n735), .B2(n1399), .ZN(n1318) );
  OAI221_X1 U5546 ( .B1(n2086), .B2(n7545), .C1(n2088), .C2(n4795), .A(n1321), 
        .ZN(n1320) );
  OAI222_X1 U5547 ( .A1(n727), .A2(n1122), .B1(n741), .B2(n1327), .C1(n2082), 
        .C2(n1257), .ZN(n1319) );
  INV_X1 U5548 ( .A(n1087), .ZN(n2084) );
  OAI22_X1 U5549 ( .A1(n2086), .A2(n7432), .B1(n2092), .B2(n6728), .ZN(n1087)
         );
  INV_X1 U5550 ( .A(n5450), .ZN(n2191) );
  OAI221_X1 U5551 ( .B1(n750), .B2(n2825), .C1(n2195), .C2(n6701), .A(n2986), 
        .ZN(n5450) );
  INV_X1 U5552 ( .A(n5452), .ZN(n2986) );
  OAI22_X1 U5553 ( .A1(n7552), .A2(n2194), .B1(n7561), .B2(n2197), .ZN(n5452)
         );
  OAI221_X1 U5554 ( .B1(n727), .B2(n6866), .C1(n728), .C2(n6813), .A(n2078), 
        .ZN(n823) );
  INV_X1 U5555 ( .A(n825), .ZN(n2078) );
  OAI22_X1 U5556 ( .A1(n6876), .A2(n2082), .B1(n826), .B2(n741), .ZN(n825) );
  AND2_X1 U5557 ( .A1(n827), .A2(n2176), .ZN(n826) );
  INV_X1 U5558 ( .A(n730), .ZN(n2018) );
  OAI21_X1 U5559 ( .B1(n6730), .B2(n2082), .A(n732), .ZN(n730) );
  OAI221_X1 U5560 ( .B1(n727), .B2(n6687), .C1(n728), .C2(n6689), .A(n2016), 
        .ZN(n1154) );
  INV_X1 U5561 ( .A(n1156), .ZN(n2016) );
  OAI21_X1 U5562 ( .B1(n6688), .B2(n2082), .A(n732), .ZN(n1156) );
  OAI221_X1 U5563 ( .B1(n727), .B2(n6857), .C1(n728), .C2(n6804), .A(n2080), 
        .ZN(n1209) );
  INV_X1 U5564 ( .A(n1211), .ZN(n2080) );
  OAI21_X1 U5565 ( .B1(n6877), .B2(n2082), .A(n2096), .ZN(n1211) );
  INV_X1 U5566 ( .A(n1167), .ZN(n2028) );
  OAI221_X1 U5567 ( .B1(n728), .B2(n6818), .C1(n2094), .C2(n6801), .A(n2035), 
        .ZN(n1167) );
  INV_X1 U5568 ( .A(n1169), .ZN(n2035) );
  OAI22_X1 U5569 ( .A1(n6916), .A2(n727), .B1(n6896), .B2(n2082), .ZN(n1169)
         );
  INV_X1 U5570 ( .A(n834), .ZN(n2075) );
  OAI22_X1 U5571 ( .A1(n6761), .A2(n727), .B1(n6762), .B2(n2082), .ZN(n834) );
  OAI221_X1 U5572 ( .B1(n728), .B2(n6814), .C1(n2094), .C2(n6797), .A(n2070), 
        .ZN(n849) );
  INV_X1 U5573 ( .A(n851), .ZN(n2070) );
  OAI22_X1 U5574 ( .A1(n6867), .A2(n727), .B1(n6891), .B2(n2082), .ZN(n851) );
  AND2_X1 U5575 ( .A1(Ntkbx6[16]), .A2(n4043), .ZN(Ehihu6) );
  OAI22_X1 U5576 ( .A1(n701), .A2(n1671), .B1(n2297), .B2(n4774), .ZN(n4043)
         );
  AND2_X1 U5577 ( .A1(Nvkbx6[21]), .A2(n3974), .ZN(G7lhu6) );
  OAI22_X1 U5578 ( .A1(n733), .A2(n4772), .B1(n736), .B2(n1631), .ZN(n3974) );
  AND2_X1 U5579 ( .A1(Nvkbx6[20]), .A2(n2337), .ZN(Y5lhu6) );
  OAI22_X1 U5580 ( .A1(n2264), .A2(n4184), .B1(n736), .B2(n1633), .ZN(n2337)
         );
  AND2_X1 U5581 ( .A1(Nvkbx6[11]), .A2(n4030), .ZN(Eukhu6) );
  OAI22_X1 U5582 ( .A1(n733), .A2(n4806), .B1(n736), .B2(n1738), .ZN(n4030) );
  OAI221_X1 U5583 ( .B1(n2094), .B2(n6724), .C1(n456), .C2(n6723), .A(n2031), 
        .ZN(n1121) );
  INV_X1 U5584 ( .A(n1123), .ZN(n2031) );
  OAI22_X1 U5585 ( .A1(n6722), .A2(n728), .B1(n6720), .B2(n727), .ZN(n1123) );
  NOR3_X1 U5586 ( .A1(n2118), .A2(n6637), .A3(n354), .ZN(n711) );
  NOR4_X1 U5587 ( .A1(n7519), .A2(n7359), .A3(n7329), .A4(n7325), .ZN(n1589)
         );
  OAI21_X2 U5588 ( .B1(n484), .B2(n963), .A(n397), .ZN(n180) );
  NOR4_X1 U5589 ( .A1(n487), .A2(n488), .A3(n489), .A4(n490), .ZN(n484) );
  OAI21_X1 U5590 ( .B1(n493), .B2(n494), .A(n495), .ZN(n488) );
  NOR3_X1 U5591 ( .A1(n1925), .A2(n7510), .A3(n3628), .ZN(n490) );
  OAI22_X1 U5592 ( .A1(n3104), .A2(n2358), .B1(n2712), .B2(n1251), .ZN(n5527)
         );
  OAI21_X1 U5593 ( .B1(n924), .B2(n925), .A(n2102), .ZN(n910) );
  NAND4_X1 U5594 ( .A1(n7429), .A2(n7655), .A3(n926), .A4(n7657), .ZN(n925) );
  NAND4_X1 U5595 ( .A1(n7681), .A2(n7693), .A3(n7667), .A4(n927), .ZN(n924) );
  AND2_X1 U5596 ( .A1(n7664), .A2(n7661), .ZN(n926) );
  NOR4_X1 U5597 ( .A1(n354), .A2(n1431), .A3(n2118), .A4(n7507), .ZN(n1412) );
  AOI222_X1 U5598 ( .A1(n3333), .A2(n3725), .B1(n4691), .B2(HRDATA[28]), .C1(
        n2822), .C2(n4705), .ZN(n4632) );
  INV_X1 U5599 ( .A(n1091), .ZN(n2822) );
  AOI222_X1 U5600 ( .A1(n2364), .A2(n3725), .B1(n4691), .B2(HRDATA[7]), .C1(
        n1228), .C2(n4705), .ZN(n4143) );
  NOR2_X1 U5601 ( .A1(n963), .A2(n7507), .ZN(n1996) );
  NOR2_X1 U5602 ( .A1(n7399), .A2(n225), .ZN(n1576) );
  NOR2_X1 U5603 ( .A1(n961), .A2(n7507), .ZN(n451) );
  NOR2_X1 U5604 ( .A1(n7510), .A2(n7399), .ZN(n2893) );
  NOR2_X1 U5605 ( .A1(n963), .A2(n7507), .ZN(n450) );
  AOI221_X1 U5606 ( .B1(n1302), .B2(n4705), .C1(n4691), .C2(HRDATA[3]), .A(
        n2342), .ZN(n4836) );
  INV_X1 U5607 ( .A(n5664), .ZN(n2342) );
  AOI22_X1 U5608 ( .A1(n4717), .A2(n3382), .B1(n4690), .B2(n3380), .ZN(n5664)
         );
  AOI221_X1 U5609 ( .B1(n3365), .B2(n4690), .C1(n4691), .C2(HRDATA[10]), .A(
        n4692), .ZN(n4411) );
  OAI22_X1 U5610 ( .A1(n2712), .A2(n2832), .B1(n3106), .B2(n2396), .ZN(n4692)
         );
  OAI22_X1 U5611 ( .A1(n7529), .A2(n3860), .B1(n2643), .B2(n3804), .ZN(n6503)
         );
  OAI21_X1 U5612 ( .B1(n5571), .B2(n5564), .A(n5572), .ZN(n4636) );
  AOI21_X1 U5613 ( .B1(n7626), .B2(n5573), .A(n429), .ZN(n5571) );
  OAI21_X1 U5614 ( .B1(n266), .B2(n3730), .A(n3768), .ZN(n5573) );
  NOR4_X1 U5615 ( .A1(Affpw6[1]), .A2(n4247), .A3(n4248), .A4(n4249), .ZN(
        n3434) );
  NOR4_X1 U5616 ( .A1(n7400), .A2(n7530), .A3(n4261), .A4(n4364), .ZN(n4247)
         );
  OAI21_X1 U5617 ( .B1(n4251), .B2(n3811), .A(n4252), .ZN(n4248) );
  NOR2_X1 U5618 ( .A1(n4993), .A2(n7519), .ZN(n1592) );
  NOR4_X1 U5619 ( .A1(n5528), .A2(n5529), .A3(n5530), .A4(n5531), .ZN(n1251)
         );
  OAI222_X1 U5620 ( .A1(n2193), .A2(n7639), .B1(n2199), .B2(n6775), .C1(n2200), 
        .C2(n7634), .ZN(n5530) );
  OAI222_X1 U5621 ( .A1(n4729), .A2(n7633), .B1(n2198), .B2(n6778), .C1(n4730), 
        .C2(n6578), .ZN(n5529) );
  OAI221_X1 U5622 ( .B1(n2194), .B2(n7636), .C1(n2196), .C2(n7637), .A(n2901), 
        .ZN(n5531) );
  AOI222_X1 U5624 ( .A1(n438), .A2(Nxkbx6[6]), .B1(n4834), .B2(vis_ipsr_o[5]), 
        .C1(n5101), .C2(n2551), .ZN(n3396) );
  AOI21_X1 U5625 ( .B1(n5030), .B2(n5031), .A(n961), .ZN(n3022) );
  AOI221_X1 U5626 ( .B1(n7283), .B2(n1938), .C1(n1642), .C2(n1902), .A(n4304), 
        .ZN(n5031) );
  AOI221_X1 U5627 ( .B1(n1584), .B2(n2921), .C1(n1672), .C2(n5034), .A(n5035), 
        .ZN(n5030) );
  OAI211_X1 U5628 ( .C1(n1612), .C2(n2260), .A(n5038), .B(n5039), .ZN(n5034)
         );
  NOR2_X1 U5629 ( .A1(n4123), .A2(n6569), .ZN(n911) );
  NAND4_X1 U5630 ( .A1(n7507), .A2(n3712), .A3(n1428), .A4(n1376), .ZN(n705)
         );
  OAI21_X1 U5631 ( .B1(n4548), .B2(n2234), .A(n1430), .ZN(n1428) );
  AOI221_X1 U5632 ( .B1(n1149), .B2(n4705), .C1(n3378), .C2(n4690), .A(n2353), 
        .ZN(n4262) );
  INV_X1 U5633 ( .A(n4767), .ZN(n2353) );
  AOI22_X1 U5634 ( .A1(n4717), .A2(n3371), .B1(HRDATA[1]), .B2(n4691), .ZN(
        n4767) );
  OR2_X1 U5635 ( .A1(n4152), .A2(n7533), .ZN(n3878) );
  OAI21_X1 U5636 ( .B1(n4296), .B2(n1699), .A(n1837), .ZN(n1917) );
  NOR3_X1 U5637 ( .A1(n2251), .A2(n7519), .A3(n3628), .ZN(n4296) );
  OAI211_X1 U5638 ( .C1(n5473), .C2(n4726), .A(n5474), .B(n5475), .ZN(n4525)
         );
  NAND3_X1 U5639 ( .A1(n3346), .A2(n2349), .A3(n3725), .ZN(n5474) );
  AOI22_X1 U5640 ( .A1(HRDATA[30]), .A2(n4691), .B1(n4705), .B2(n888), .ZN(
        n5475) );
  OAI222_X1 U5641 ( .A1(n8359), .A2(n4788), .B1(n2202), .B2(n7635), .C1(n1893), 
        .C2(n7445), .ZN(n5528) );
  INV_X1 U5642 ( .A(STCALIB[6]), .ZN(n8359) );
  NAND4_X1 U5643 ( .A1(n1166), .A2(n2096), .A3(n1234), .A4(n1235), .ZN(n7909)
         );
  AOI22_X1 U5644 ( .A1(n883), .A2(n1237), .B1(n1124), .B2(n6679), .ZN(n1234)
         );
  AOI222_X1 U5645 ( .A1(n856), .A2(n4297), .B1(n838), .B2(HRDATA[6]), .C1(n239), .C2(Jshpw6[6]), .ZN(n1235) );
  NAND4_X1 U5646 ( .A1(n1238), .A2(n1239), .A3(n1240), .A4(n1241), .ZN(n1237)
         );
  OAI221_X1 U5647 ( .B1(n7501), .B2(n2111), .C1(n7514), .C2(n1376), .A(n1394), 
        .ZN(n7931) );
  AOI222_X1 U5648 ( .A1(n2119), .A2(n4721), .B1(n715), .B2(HRDATA[26]), .C1(
        n716), .C2(HRDATA[10]), .ZN(n1394) );
  OAI221_X1 U5649 ( .B1(n7495), .B2(n2111), .C1(n7523), .C2(n1376), .A(n1385), 
        .ZN(n7927) );
  AOI222_X1 U5650 ( .A1(n2119), .A2(n4704), .B1(n715), .B2(HRDATA[21]), .C1(
        n716), .C2(HRDATA[5]), .ZN(n1385) );
  OAI221_X1 U5651 ( .B1(n7502), .B2(n2111), .C1(n270), .C2(n1376), .A(n1396), 
        .ZN(n7932) );
  AOI222_X1 U5652 ( .A1(n2119), .A2(n4724), .B1(n715), .B2(HRDATA[27]), .C1(
        n716), .C2(HRDATA[11]), .ZN(n1396) );
  OAI221_X1 U5653 ( .B1(n7545), .B2(n180), .C1(n3012), .C2(n397), .A(n404), 
        .ZN(n7823) );
  AOI222_X1 U5654 ( .A1(n241), .A2(\eq_3147/A[0] ), .B1(n1852), .B2(
        vis_pc_o[1]), .C1(n182), .C2(vis_ipsr_o[2]), .ZN(n404) );
  OAI221_X1 U5655 ( .B1(n7334), .B2(n928), .C1(n7313), .C2(n913), .A(n2034), 
        .ZN(n8050) );
  AOI222_X1 U5656 ( .A1(n236), .A2(n3877), .B1(ECOREVNUM[27]), .B2(n542), .C1(
        n544), .C2(n4038), .ZN(n2034) );
  OAI221_X1 U5657 ( .B1(n7409), .B2(n928), .C1(n7334), .C2(n913), .A(n2032), 
        .ZN(n8049) );
  AOI222_X1 U5658 ( .A1(n236), .A2(n3125), .B1(ECOREVNUM[26]), .B2(n542), .C1(
        n544), .C2(n4038), .ZN(n2032) );
  OAI221_X1 U5659 ( .B1(n7346), .B2(n928), .C1(n7431), .C2(n913), .A(n2030), 
        .ZN(n8048) );
  AOI222_X1 U5660 ( .A1(n236), .A2(n3004), .B1(ECOREVNUM[24]), .B2(n542), .C1(
        n544), .C2(n4040), .ZN(n2030) );
  AOI222_X1 U5661 ( .A1(n3481), .A2(vis_pc_o[27]), .B1(n2961), .B2(n8261), 
        .C1(n1064), .C2(HRDATA[28]), .ZN(n1093) );
  AOI222_X1 U5662 ( .A1(n3476), .A2(E1hpw6[4]), .B1(ECOREVNUM[8]), .B2(n1075), 
        .C1(ECOREVNUM[4]), .C2(n1066), .ZN(n1262) );
  NOR4_X1 U5663 ( .A1(n2955), .A2(n1058), .A3(n1059), .A4(n2826), .ZN(n1056)
         );
  OAI21_X1 U5664 ( .B1(n4782), .B2(n1020), .A(n3443), .ZN(n1058) );
  INV_X1 U5665 ( .A(n1062), .ZN(n2955) );
  AOI221_X1 U5666 ( .B1(n8082), .B2(n2961), .C1(HRDATA[5]), .C2(n1064), .A(
        n1065), .ZN(n1062) );
  NOR4_X1 U5667 ( .A1(n1265), .A2(n1266), .A3(n1059), .A4(n1267), .ZN(n1264)
         );
  OAI221_X1 U5668 ( .B1(n6827), .B2(n1004), .C1(n7546), .C2(n1009), .A(n3446), 
        .ZN(n1265) );
  OAI222_X1 U5669 ( .A1(n4783), .A2(n1020), .B1(n8325), .B2(n2965), .C1(n6647), 
        .C2(n1008), .ZN(n1266) );
  INV_X1 U5670 ( .A(n1280), .ZN(n3446) );
  NOR3_X1 U5671 ( .A1(n3634), .A2(n1894), .A3(n914), .ZN(n1892) );
  AOI222_X1 U5672 ( .A1(n883), .A2(n900), .B1(n838), .B2(HRDATA[22]), .C1(n839), .C2(vis_pc_o[21]), .ZN(n899) );
  OAI211_X1 U5673 ( .C1(n7259), .C2(n1376), .A(n1377), .B(n1378), .ZN(n7925)
         );
  AOI22_X1 U5674 ( .A1(n6641), .A2(n2119), .B1(n711), .B2(n4855), .ZN(n1377)
         );
  AOI222_X1 U5675 ( .A1(n716), .A2(HRDATA[3]), .B1(n1379), .B2(n2131), .C1(
        n715), .C2(HRDATA[19]), .ZN(n1378) );
  OAI211_X1 U5676 ( .C1(n7519), .C2(n1376), .A(n1389), .B(n1390), .ZN(n7929)
         );
  AOI22_X1 U5677 ( .A1(n6640), .A2(n2119), .B1(n711), .B2(n3538), .ZN(n1389)
         );
  AOI222_X1 U5678 ( .A1(n716), .A2(HRDATA[7]), .B1(n1391), .B2(n2131), .C1(
        n715), .C2(HRDATA[23]), .ZN(n1390) );
  OAI22_X1 U5679 ( .A1(n7286), .A2(n3860), .B1(n2618), .B2(n3804), .ZN(n6445)
         );
  NOR4_X1 U5680 ( .A1(n2960), .A2(n1227), .A3(n1059), .A4(n1228), .ZN(n1225)
         );
  OAI21_X1 U5681 ( .B1(n4811), .B2(n1020), .A(n3443), .ZN(n1227) );
  INV_X1 U5682 ( .A(n1229), .ZN(n2960) );
  AOI221_X1 U5683 ( .B1(n4940), .B2(n2961), .C1(HRDATA[7]), .C2(n1064), .A(
        n1230), .ZN(n1229) );
  AOI222_X1 U5684 ( .A1(STCALIB[7]), .A2(n2973), .B1(n2975), .B2(n8235), .C1(
        n2976), .C2(Tzfpw6[7]), .ZN(n5931) );
  AOI222_X1 U5685 ( .A1(STCALIB[22]), .A2(n2973), .B1(n2975), .B2(n8197), .C1(
        n2976), .C2(Tzfpw6[22]), .ZN(n5502) );
  NOR2_X1 U5686 ( .A1(n7433), .A2(n7381), .ZN(n1755) );
  NOR4_X1 U5687 ( .A1(n996), .A2(n997), .A3(n998), .A4(n999), .ZN(n978) );
  OAI221_X1 U5688 ( .B1(n7452), .B2(n125), .C1(n7414), .C2(n1000), .A(n3404), 
        .ZN(n996) );
  INV_X1 U5689 ( .A(n1002), .ZN(n3404) );
  NOR2_X1 U5690 ( .A1(n4123), .A2(n6898), .ZN(n119) );
  NOR2_X1 U5691 ( .A1(n475), .A2(n7516), .ZN(n472) );
  AOI21_X1 U5692 ( .B1(HWDATA[26]), .B2(n3687), .A(n3691), .ZN(n1777) );
  NOR4_X1 U5693 ( .A1(n1891), .A2(n1890), .A3(n7570), .A4(n7352), .ZN(n3691)
         );
  NOR4_X1 U5694 ( .A1(n1328), .A2(n1329), .A3(n1330), .A4(n1841), .ZN(n1327)
         );
  OAI222_X1 U5695 ( .A1(n113), .A2(n7456), .B1(n988), .B2(n6792), .C1(n984), 
        .C2(n7463), .ZN(n1330) );
  INV_X1 U5696 ( .A(n1332), .ZN(n1841) );
  OAI221_X1 U5697 ( .B1(n1005), .B2(n7459), .C1(n2965), .C2(n8327), .A(n3472), 
        .ZN(n1329) );
  NOR3_X1 U5698 ( .A1(n3763), .A2(n7530), .A3(n3712), .ZN(n4464) );
  OAI221_X1 U5699 ( .B1(n7431), .B2(n928), .C1(n7409), .C2(n913), .A(n539), 
        .ZN(n7833) );
  AOI221_X1 U5700 ( .B1(n236), .B2(n8205), .C1(ECOREVNUM[25]), .C2(n542), .A(
        n543), .ZN(n539) );
  AND3_X1 U5701 ( .A1(n544), .A2(n1817), .A3(n545), .ZN(n543) );
  OAI21_X1 U5702 ( .B1(n7349), .B2(n7348), .A(n4040), .ZN(n545) );
  OAI221_X1 U5703 ( .B1(n7426), .B2(n881), .C1(n7646), .C2(n2098), .A(n1131), 
        .ZN(n7900) );
  AOI221_X1 U5704 ( .B1(n2004), .B2(\Aphpw6[2] ), .C1(n883), .C2(n1133), .A(
        n2001), .ZN(n1131) );
  NAND4_X1 U5705 ( .A1(n1139), .A2(n1140), .A3(n2963), .A4(n1142), .ZN(n1133)
         );
  INV_X1 U5706 ( .A(n1147), .ZN(n2963) );
  OAI221_X1 U5707 ( .B1(n1769), .B2(n1849), .C1(n7408), .C2(n180), .A(n351), 
        .ZN(n7801) );
  AOI221_X1 U5708 ( .B1(vis_pc_o[8]), .B2(n1852), .C1(n183), .C2(n3922), .A(
        n353), .ZN(n351) );
  NOR3_X1 U5709 ( .A1(n1847), .A2(n7628), .A3(n354), .ZN(n353) );
  OAI221_X1 U5710 ( .B1(n7627), .B2(n180), .C1(n397), .C2(n3259), .A(n440), 
        .ZN(n7826) );
  AOI221_X1 U5711 ( .B1(n182), .B2(vis_ipsr_o[1]), .C1(n1852), .C2(vis_pc_o[0]), .A(n441), .ZN(n440) );
  AND4_X1 U5712 ( .A1(n2614), .A2(n443), .A3(n444), .A4(n241), .ZN(n441) );
  AOI221_X1 U5713 ( .B1(ECOREVNUM[5]), .B2(n1066), .C1(n3476), .C2(E1hpw6[5]), 
        .A(n1069), .ZN(n1055) );
  OAI22_X1 U5714 ( .A1(n6779), .A2(n985), .B1(n6781), .B2(n989), .ZN(n1069) );
  AOI221_X1 U5715 ( .B1(n3474), .B2(K7hpw6[6]), .C1(ECOREVNUM[18]), .C2(n1070), 
        .A(n1255), .ZN(n1240) );
  NAND2_X1 U5716 ( .A1(n3480), .A2(n992), .ZN(n1255) );
  AOI221_X1 U5717 ( .B1(ECOREVNUM[16]), .B2(n1070), .C1(ECOREVNUM[12]), .C2(
        n1074), .A(n1281), .ZN(n1263) );
  OAI211_X1 U5718 ( .C1(n6847), .C2(n990), .A(n3480), .B(n1282), .ZN(n1281) );
  AOI221_X1 U5719 ( .B1(Ezohu6), .B2(n7598), .C1(F3phu6), .C2(n7584), .A(n2481), .ZN(n3680) );
  INV_X1 U5720 ( .A(n3731), .ZN(n2481) );
  AOI222_X1 U5721 ( .A1(n7602), .A2(Cyohu6), .B1(n3645), .B2(A4phu6), .C1(
        n7587), .C2(D2phu6), .ZN(n3731) );
  AOI221_X1 U5722 ( .B1(ECOREVNUM[7]), .B2(n1066), .C1(n3476), .C2(E1hpw6[7]), 
        .A(n1232), .ZN(n1224) );
  OAI22_X1 U5723 ( .A1(n6865), .A2(n985), .B1(n6812), .B2(n989), .ZN(n1232) );
  AOI221_X1 U5724 ( .B1(ECOREVNUM[17]), .B2(n1070), .C1(n3474), .C2(K7hpw6[5]), 
        .A(n1073), .ZN(n1054) );
  AOI221_X1 U5725 ( .B1(n1064), .B2(HRDATA[1]), .C1(n3481), .C2(vis_pc_o[0]), 
        .A(n1148), .ZN(n1140) );
  OAI22_X1 U5726 ( .A1(n7453), .A2(n125), .B1(n7467), .B2(n1008), .ZN(n1148)
         );
  OAI211_X1 U5727 ( .C1(n7330), .C2(n2714), .A(n6527), .B(n6535), .ZN(n5194)
         );
  AOI22_X1 U5728 ( .A1(n6529), .A2(n3576), .B1(n6530), .B2(n2466), .ZN(n6535)
         );
  NOR2_X1 U5729 ( .A1(n3759), .A2(n2306), .ZN(Npghu6) );
  AOI221_X1 U5730 ( .B1(n2500), .B2(n906), .C1(n7549), .C2(NMI), .A(n2305), 
        .ZN(n3759) );
  AOI221_X1 U5731 ( .B1(n2976), .B2(Tzfpw6[16]), .C1(STCALIB[16]), .C2(n2973), 
        .A(n5405), .ZN(n5404) );
  OAI22_X1 U5732 ( .A1(n7361), .A2(n2202), .B1(n7589), .B2(n4730), .ZN(n5405)
         );
  OAI221_X1 U5733 ( .B1(n4755), .B2(n3344), .C1(n3101), .C2(n4726), .A(n4757), 
        .ZN(n4270) );
  AOI21_X1 U5734 ( .B1(n3725), .B2(n3318), .A(n4717), .ZN(n4755) );
  AOI22_X1 U5735 ( .A1(n4705), .A2(n1164), .B1(HRDATA[25]), .B2(n4691), .ZN(
        n4757) );
  OAI221_X1 U5736 ( .B1(n3102), .B2(n4726), .C1(n4727), .C2(n3342), .A(n4728), 
        .ZN(n4414) );
  AOI21_X1 U5737 ( .B1(n3725), .B2(n3319), .A(n4717), .ZN(n4727) );
  AOI22_X1 U5738 ( .A1(n4705), .A2(n1032), .B1(HRDATA[26]), .B2(n4691), .ZN(
        n4728) );
  OAI211_X1 U5739 ( .C1(n439), .C2(n1801), .A(n4819), .B(n4820), .ZN(n3432) );
  AOI22_X1 U5740 ( .A1(n635), .A2(n3981), .B1(vis_ipsr_o[3]), .B2(n4834), .ZN(
        n4819) );
  AOI221_X1 U5742 ( .B1(n2551), .B2(n4821), .C1(n4822), .C2(n4823), .A(
        Affpw6[3]), .ZN(n4820) );
  OAI22_X1 U5743 ( .A1(n2732), .A2(n4824), .B1(n4825), .B2(n3796), .ZN(n4822)
         );
  OAI222_X1 U5744 ( .A1(n2098), .A2(n6656), .B1(n741), .B2(n2827), .C1(n881), 
        .C2(n7428), .ZN(n1129) );
  OAI221_X1 U5745 ( .B1(n5671), .B2(n3336), .C1(n4735), .C2(n4726), .A(n5672), 
        .ZN(n4840) );
  AOI21_X1 U5746 ( .B1(n3725), .B2(n3340), .A(n4717), .ZN(n5671) );
  AOI22_X1 U5747 ( .A1(HRDATA[27]), .A2(n4691), .B1(n4705), .B2(n2834), .ZN(
        n5672) );
  INV_X1 U5748 ( .A(n1158), .ZN(n2834) );
  OAI21_X1 U5749 ( .B1(n3253), .B2(n4818), .A(n3254), .ZN(n2480) );
  AOI21_X1 U5750 ( .B1(n1620), .B2(n1571), .A(n3277), .ZN(n3253) );
  OAI21_X1 U5751 ( .B1(n3255), .B2(n3256), .A(N701), .ZN(n3254) );
  NOR3_X1 U5752 ( .A1(n3766), .A2(n7497), .A3(n266), .ZN(n3277) );
  OAI211_X1 U5753 ( .C1(n7274), .C2(n2714), .A(n6527), .B(n6528), .ZN(n5173)
         );
  AOI22_X1 U5754 ( .A1(n6529), .A2(n4506), .B1(n6530), .B2(n5307), .ZN(n6528)
         );
  NOR2_X1 U5756 ( .A1(n4123), .A2(n6872), .ZN(n710) );
  OAI22_X1 U5757 ( .A1(n7530), .A2(n3860), .B1(n2621), .B2(n3804), .ZN(n6481)
         );
  OAI21_X1 U5758 ( .B1(n7476), .B2(N701), .A(n1968), .ZN(n8011) );
  NAND4_X1 U5759 ( .A1(n1969), .A2(n3439), .A3(n1971), .A4(HALTED), .ZN(n1968)
         );
  NOR2_X1 U5760 ( .A1(n7412), .A2(n963), .ZN(n1971) );
  OAI22_X1 U5761 ( .A1(n3449), .A2(n3851), .B1(n3688), .B2(n3689), .ZN(n2172)
         );
  AOI21_X1 U5762 ( .B1(n226), .B2(HWDATA[28]), .A(n7599), .ZN(n3688) );
  OAI21_X1 U5763 ( .B1(n8333), .B2(n8279), .A(n3448), .ZN(n3689) );
  OAI21_X1 U5764 ( .B1(n7283), .B2(n4361), .A(n4362), .ZN(n4358) );
  OAI21_X1 U5765 ( .B1(n1902), .B2(n875), .A(n521), .ZN(n4362) );
  AOI22_X1 U5766 ( .A1(n1624), .A2(n7373), .B1(n1620), .B2(n479), .ZN(n4361)
         );
  AND2_X1 U5767 ( .A1(n4718), .A2(n4719), .ZN(n1021) );
  AOI221_X1 U5768 ( .B1(n2866), .B2(n4061), .C1(n2975), .C2(n4163), .A(n4722), 
        .ZN(n4719) );
  AOI221_X1 U5769 ( .B1(n2976), .B2(Tzfpw6[18]), .C1(STCALIB[18]), .C2(n2973), 
        .A(n4714), .ZN(n4718) );
  NAND2_X1 U5770 ( .A1(n1589), .A2(n7518), .ZN(n1493) );
  NOR2_X1 U5771 ( .A1(n7414), .A2(n7415), .ZN(n6162) );
  NAND2_X1 U5772 ( .A1(n7491), .A2(HRESP), .ZN(n2430) );
  AOI221_X1 U5773 ( .B1(n7435), .B2(n2475), .C1(n7705), .C2(n699), .A(n3683), 
        .ZN(n3681) );
  INV_X1 U5774 ( .A(n1634), .ZN(n2475) );
  OAI221_X1 U5775 ( .B1(n1777), .B2(n3617), .C1(n8280), .C2(n2172), .A(n3685), 
        .ZN(n3683) );
  NAND3_X1 U5776 ( .A1(HWDATA[28]), .A2(n3775), .A3(n3687), .ZN(n3685) );
  OAI222_X1 U5777 ( .A1(n7422), .A2(n881), .B1(n1220), .B2(n741), .C1(n2098), 
        .C2(n8284), .ZN(n7908) );
  AND4_X1 U5778 ( .A1(n1222), .A2(n1223), .A3(n1224), .A4(n1225), .ZN(n1220)
         );
  AOI22_X1 U5779 ( .A1(ECOREVNUM[15]), .A2(n1074), .B1(ECOREVNUM[11]), .B2(
        n1075), .ZN(n1222) );
  AOI22_X1 U5780 ( .A1(n3474), .A2(K7hpw6[7]), .B1(ECOREVNUM[19]), .B2(n1070), 
        .ZN(n1223) );
  OAI21_X1 U5781 ( .B1(n1982), .B2(n5256), .A(n1987), .ZN(n8016) );
  NAND4_X1 U5782 ( .A1(n1643), .A2(n7533), .A3(n1988), .A4(n4512), .ZN(n1987)
         );
  OAI22_X1 U5783 ( .A1(vis_pc_o[1]), .A2(n3765), .B1(n457), .B2(n810), .ZN(
        n1988) );
  OAI221_X1 U5784 ( .B1(n7499), .B2(n2111), .C1(n7518), .C2(n1376), .A(n1400), 
        .ZN(n7934) );
  AOI222_X1 U5785 ( .A1(n2119), .A2(n4713), .B1(n715), .B2(HRDATA[24]), .C1(
        n716), .C2(HRDATA[8]), .ZN(n1400) );
  OAI221_X1 U5786 ( .B1(n909), .B2(n916), .C1(n7419), .C2(N701), .A(n910), 
        .ZN(n7886) );
  XNOR2_X1 U5787 ( .A(n4402), .B(n918), .ZN(n916) );
  OAI221_X1 U5788 ( .B1(n909), .B2(n921), .C1(n7448), .C2(N701), .A(n910), 
        .ZN(n7888) );
  XNOR2_X1 U5789 ( .A(n4145), .B(n922), .ZN(n921) );
  OAI221_X1 U5790 ( .B1(n909), .B2(n923), .C1(n7388), .C2(N701), .A(n910), 
        .ZN(n7889) );
  AOI22_X1 U5791 ( .A1(n856), .A2(n6644), .B1(Tnhpw6[2]), .B2(n239), .ZN(n1321) );
  OAI221_X1 U5792 ( .B1(n7503), .B2(n2111), .C1(n7510), .C2(n1376), .A(n1398), 
        .ZN(n7933) );
  AOI222_X1 U5793 ( .A1(n2119), .A2(n5258), .B1(n715), .B2(HRDATA[28]), .C1(
        n716), .C2(HRDATA[12]), .ZN(n1398) );
  AOI221_X1 U5794 ( .B1(n4691), .B2(HRDATA[21]), .C1(n3318), .C2(n4717), .A(
        n5325), .ZN(n4594) );
  OAI22_X1 U5795 ( .A1(n2712), .A2(n2833), .B1(n3104), .B2(n2423), .ZN(n5325)
         );
  INV_X1 U5796 ( .A(n3312), .ZN(n2423) );
  OAI221_X1 U5797 ( .B1(n6750), .B2(n2133), .C1(n220), .C2(n4807), .A(n348), 
        .ZN(n7799) );
  AOI22_X1 U5798 ( .A1(n241), .A2(\eq_3147/A[8] ), .B1(n1851), .B2(n8171), 
        .ZN(n348) );
  OAI221_X1 U5799 ( .B1(n6900), .B2(n2133), .C1(n220), .C2(n4816), .A(n372), 
        .ZN(n7810) );
  AOI22_X1 U5800 ( .A1(n241), .A2(\eq_3147/A[4] ), .B1(n1851), .B2(n6679), 
        .ZN(n372) );
  OAI221_X1 U5801 ( .B1(n6756), .B2(n2133), .C1(n220), .C2(n4806), .A(n342), 
        .ZN(n7796) );
  AOI22_X1 U5802 ( .A1(n241), .A2(\eq_3147/A[9] ), .B1(n1851), .B2(n8163), 
        .ZN(n342) );
  OAI221_X1 U5803 ( .B1(n6875), .B2(n2133), .C1(n220), .C2(n4805), .A(n333), 
        .ZN(n7792) );
  AOI22_X1 U5804 ( .A1(n241), .A2(\eq_3147/A[10] ), .B1(n1851), .B2(n8103), 
        .ZN(n333) );
  OAI221_X1 U5805 ( .B1(n6889), .B2(n2133), .C1(n220), .C2(n4811), .A(n369), 
        .ZN(n7808) );
  AOI22_X1 U5806 ( .A1(n241), .A2(\eq_3147/A[5] ), .B1(n1851), .B2(n4940), 
        .ZN(n369) );
  OAI221_X1 U5807 ( .B1(n6906), .B2(n2133), .C1(n220), .C2(n4774), .A(n309), 
        .ZN(n7780) );
  AOI22_X1 U5808 ( .A1(n241), .A2(\eq_3147/A[14] ), .B1(n1851), .B2(n4185), 
        .ZN(n309) );
  OAI221_X1 U5809 ( .B1(n6902), .B2(n2133), .C1(n220), .C2(n4810), .A(n363), 
        .ZN(n7805) );
  AOI22_X1 U5810 ( .A1(n241), .A2(\eq_3147/A[6] ), .B1(n1851), .B2(n4009), 
        .ZN(n363) );
  OAI221_X1 U5811 ( .B1(n6908), .B2(n2133), .C1(n220), .C2(n4802), .A(n327), 
        .ZN(n7789) );
  AOI22_X1 U5812 ( .A1(n241), .A2(\eq_3147/A[11] ), .B1(n1851), .B2(n3041), 
        .ZN(n327) );
  NAND2_X1 U5813 ( .A1(n445), .A2(n180), .ZN(n220) );
  OAI21_X1 U5814 ( .B1(n446), .B2(n4738), .A(n447), .ZN(n445) );
  AOI21_X1 U5815 ( .B1(n7259), .B2(n4341), .A(n449), .ZN(n446) );
  NOR3_X1 U5816 ( .A1(n2430), .A2(n7332), .A3(n5786), .ZN(n5785) );
  OAI221_X1 U5817 ( .B1(n5268), .B2(n3338), .C1(n1085), .C2(n2712), .A(n5269), 
        .ZN(n4590) );
  AOI21_X1 U5818 ( .B1(n3725), .B2(n3339), .A(n4717), .ZN(n5268) );
  AOI22_X1 U5819 ( .A1(n2445), .A2(n5271), .B1(HRDATA[29]), .B2(n4691), .ZN(
        n5269) );
  INV_X1 U5820 ( .A(n4726), .ZN(n2445) );
  AOI211_X1 U5821 ( .C1(n3980), .C2(n762), .A(n3445), .B(n8333), .ZN(Kqthu6)
         );
  INV_X1 U5822 ( .A(n3449), .ZN(n3980) );
  NAND3_X1 U5823 ( .A1(n897), .A2(n3447), .A3(n3448), .ZN(n3445) );
  OAI21_X1 U5824 ( .B1(n3449), .B2(n3851), .A(n6584), .ZN(n3447) );
  AOI211_X1 U5825 ( .C1(n3971), .C2(n762), .A(n3953), .B(n8345), .ZN(Gothu6)
         );
  OAI211_X1 U5826 ( .C1(n3751), .C2(n8105), .A(n897), .B(n3753), .ZN(n3953) );
  INV_X1 U5827 ( .A(IRQ[12]), .ZN(n8345) );
  OAI21_X1 U5828 ( .B1(n4628), .B2(n2607), .A(n4365), .ZN(n1903) );
  NAND3_X1 U5830 ( .A1(n267), .A2(n7283), .A3(n1567), .ZN(n4365) );
  OAI221_X1 U5831 ( .B1(n7500), .B2(n2111), .C1(n7516), .C2(n1376), .A(n1392), 
        .ZN(n7930) );
  AOI222_X1 U5832 ( .A1(n2119), .A2(n4720), .B1(n715), .B2(HRDATA[25]), .C1(
        n716), .C2(HRDATA[9]), .ZN(n1392) );
  NAND3_X1 U5833 ( .A1(vis_tbit_o), .A2(n2430), .A3(n6769), .ZN(n1413) );
  NAND3_X1 U5834 ( .A1(N701), .A2(n4107), .A3(n4108), .ZN(n2851) );
  NOR3_X1 U5835 ( .A1(n7440), .A2(n6683), .A3(n7414), .ZN(n4108) );
  NAND4_X1 U5836 ( .A1(n524), .A2(n3568), .A3(n3851), .A4(n2548), .ZN(n4107)
         );
  OAI211_X1 U5837 ( .C1(n7399), .C2(n1376), .A(n2110), .B(n1417), .ZN(n7938)
         );
  AOI221_X1 U5838 ( .B1(n716), .B2(HRDATA[15]), .C1(n715), .C2(HRDATA[31]), 
        .A(n1418), .ZN(n1417) );
  INV_X1 U5839 ( .A(n1422), .ZN(n2110) );
  NOR3_X1 U5840 ( .A1(n1419), .A2(n6906), .A3(n4123), .ZN(n1418) );
  OAI211_X1 U5841 ( .C1(n7402), .C2(n2202), .A(n5407), .B(n5408), .ZN(n1219)
         );
  AOI22_X1 U5842 ( .A1(n2866), .A2(n4010), .B1(n2852), .B2(n8138), .ZN(n5407)
         );
  AOI22_X1 U5843 ( .A1(n2976), .A2(Tzfpw6[8]), .B1(STCALIB[8]), .B2(n2973), 
        .ZN(n5408) );
  OAI221_X1 U5844 ( .B1(n7450), .B2(n909), .C1(n7451), .C2(N701), .A(n910), 
        .ZN(n7882) );
  OAI221_X1 U5845 ( .B1(n915), .B2(n909), .C1(n7438), .C2(N701), .A(n910), 
        .ZN(n7885) );
  XNOR2_X1 U5846 ( .A(n7632), .B(n7437), .ZN(n915) );
  OAI221_X1 U5847 ( .B1(n919), .B2(n909), .C1(n7425), .C2(N701), .A(n910), 
        .ZN(n7887) );
  AOI21_X1 U5848 ( .B1(n7424), .B2(n918), .A(n920), .ZN(n919) );
  OAI221_X1 U5849 ( .B1(n7407), .B2(n909), .C1(n7411), .C2(N701), .A(n910), 
        .ZN(n7884) );
  OAI21_X1 U5850 ( .B1(n8315), .B2(n1413), .A(n7380), .ZN(n801) );
  OAI221_X1 U5851 ( .B1(n7504), .B2(n2111), .C1(n7433), .C2(n1376), .A(n1414), 
        .ZN(n7937) );
  AOI222_X1 U5852 ( .A1(n2119), .A2(n5266), .B1(n715), .B2(HRDATA[29]), .C1(
        n716), .C2(HRDATA[13]), .ZN(n1414) );
  OAI221_X1 U5853 ( .B1(n6708), .B2(n2133), .C1(n220), .C2(n4801), .A(n321), 
        .ZN(n7786) );
  AOI22_X1 U5854 ( .A1(n241), .A2(\eq_3147/A[12] ), .B1(n1851), .B2(n8252), 
        .ZN(n321) );
  OAI221_X1 U5855 ( .B1(n6766), .B2(n2133), .C1(n220), .C2(n4776), .A(n315), 
        .ZN(n7783) );
  AOI22_X1 U5856 ( .A1(n241), .A2(\eq_3147/A[13] ), .B1(n1851), .B2(n8116), 
        .ZN(n315) );
  OAI21_X1 U5857 ( .B1(n8300), .B2(n1413), .A(n7392), .ZN(n1411) );
  OAI221_X1 U5858 ( .B1(n1793), .B2(n1849), .C1(n7546), .C2(n180), .A(n388), 
        .ZN(n7817) );
  AOI222_X1 U5859 ( .A1(n182), .A2(vis_ipsr_o[4]), .B1(n183), .B2(n4139), .C1(
        vis_pc_o[3]), .C2(n1852), .ZN(n388) );
  OAI221_X1 U5860 ( .B1(n1798), .B2(n1849), .C1(n7547), .C2(n180), .A(n395), 
        .ZN(n7820) );
  AOI222_X1 U5861 ( .A1(n182), .A2(vis_ipsr_o[3]), .B1(n183), .B2(n4049), .C1(
        n1852), .C2(vis_pc_o[2]), .ZN(n395) );
  OAI221_X1 U5862 ( .B1(n1788), .B2(n1849), .C1(n7625), .C2(n180), .A(n381), 
        .ZN(n7814) );
  AOI222_X1 U5863 ( .A1(n182), .A2(vis_ipsr_o[5]), .B1(n183), .B2(n4409), .C1(
        vis_pc_o[4]), .C2(n1852), .ZN(n381) );
  OAI22_X1 U5864 ( .A1(n5270), .A2(n705), .B1(n2111), .B2(n7682), .ZN(n1422)
         );
  OAI221_X1 U5865 ( .B1(n1832), .B2(n719), .C1(n7683), .C2(n720), .A(n1360), 
        .ZN(n7921) );
  NAND2_X1 U5866 ( .A1(n277), .A2(n1998), .ZN(n1360) );
  OAI221_X1 U5867 ( .B1(n6911), .B2(n719), .C1(n7423), .C2(n720), .A(n1356), 
        .ZN(n7917) );
  NAND2_X1 U5868 ( .A1(n283), .A2(n1998), .ZN(n1356) );
  OAI221_X1 U5869 ( .B1(n6887), .B2(n719), .C1(n7424), .C2(n720), .A(n1357), 
        .ZN(n7918) );
  NAND2_X1 U5870 ( .A1(n279), .A2(n1998), .ZN(n1357) );
  OAI221_X1 U5871 ( .B1(n6885), .B2(n719), .C1(n7418), .C2(n720), .A(n1358), 
        .ZN(n7919) );
  NAND2_X1 U5872 ( .A1(n287), .A2(n1998), .ZN(n1358) );
  OAI221_X1 U5873 ( .B1(n7424), .B2(n881), .C1(n2098), .C2(n3883), .A(n1258), 
        .ZN(n7910) );
  AOI22_X1 U5874 ( .A1(n2004), .A2(n4144), .B1(n883), .B2(n1260), .ZN(n1258)
         );
  NAND4_X1 U5875 ( .A1(n3467), .A2(n1262), .A3(n1263), .A4(n1264), .ZN(n1260)
         );
  OAI221_X1 U5876 ( .B1(n7525), .B2(n1914), .C1(n1915), .C2(n1916), .A(n1917), 
        .ZN(n8005) );
  AOI222_X1 U5877 ( .A1(n1918), .A2(n4572), .B1(n1919), .B2(n5042), .C1(n1920), 
        .C2(n4908), .ZN(n1915) );
  OAI221_X1 U5878 ( .B1(n1011), .B2(n741), .C1(n7427), .C2(n881), .A(n1012), 
        .ZN(n7891) );
  NOR4_X1 U5879 ( .A1(n1015), .A2(n1016), .A3(n1017), .A4(n1018), .ZN(n1011)
         );
  AOI21_X1 U5880 ( .B1(n856), .B2(n4055), .A(n2000), .ZN(n1012) );
  OAI222_X1 U5881 ( .A1(n6832), .A2(n1004), .B1(n6893), .B2(n1006), .C1(n7700), 
        .C2(n1009), .ZN(n1017) );
  OAI221_X1 U5882 ( .B1(n3012), .B2(n719), .C1(n7441), .C2(n720), .A(n1359), 
        .ZN(n7920) );
  NAND2_X1 U5883 ( .A1(Vrkbx6[3]), .A2(n1998), .ZN(n1359) );
  OAI221_X1 U5884 ( .B1(n6902), .B2(n719), .C1(n7406), .C2(n720), .A(n1353), 
        .ZN(n7914) );
  NAND2_X1 U5885 ( .A1(n285), .A2(n1998), .ZN(n1353) );
  OAI221_X1 U5886 ( .B1(n6900), .B2(n719), .C1(n7632), .C2(n720), .A(n1355), 
        .ZN(n7916) );
  NAND2_X1 U5887 ( .A1(n281), .A2(n1998), .ZN(n1355) );
  OAI221_X1 U5888 ( .B1(n6889), .B2(n719), .C1(n7422), .C2(n720), .A(n1354), 
        .ZN(n7915) );
  NAND2_X1 U5889 ( .A1(n288), .A2(n1998), .ZN(n1354) );
  OAI221_X1 U5890 ( .B1(n6901), .B2(n719), .C1(n7407), .C2(n720), .A(n1352), 
        .ZN(n7913) );
  NAND2_X1 U5891 ( .A1(n290), .A2(n1998), .ZN(n1352) );
  OAI221_X1 U5892 ( .B1(n7494), .B2(n2111), .C1(n7393), .C2(n1376), .A(n1383), 
        .ZN(n7926) );
  AOI222_X1 U5893 ( .A1(n2119), .A2(n4703), .B1(n715), .B2(HRDATA[20]), .C1(
        n716), .C2(HRDATA[4]), .ZN(n1383) );
  OAI221_X1 U5894 ( .B1(n3259), .B2(n719), .C1(n7426), .C2(n720), .A(n721), 
        .ZN(n7854) );
  NAND2_X1 U5895 ( .A1(Vrkbx6[2]), .A2(n1998), .ZN(n721) );
  OAI221_X1 U5896 ( .B1(n7496), .B2(n2111), .C1(n7505), .C2(n1376), .A(n1387), 
        .ZN(n7928) );
  AOI222_X1 U5897 ( .A1(n2119), .A2(n4707), .B1(n715), .B2(HRDATA[22]), .C1(
        n716), .C2(HRDATA[6]), .ZN(n1387) );
  OAI22_X1 U5898 ( .A1(n7468), .A2(n728), .B1(n7470), .B2(n727), .ZN(n886) );
  OAI22_X1 U5899 ( .A1(n7483), .A2(n728), .B1(n7486), .B2(n727), .ZN(n1106) );
  OAI221_X1 U5900 ( .B1(n4294), .B2(n1916), .C1(n6601), .C2(n4295), .A(n1917), 
        .ZN(Cfthu6) );
  AOI221_X1 U5901 ( .B1(n1918), .B2(n470), .C1(n2374), .C2(n4932), .A(n4320), 
        .ZN(n4294) );
  AOI21_X1 U5902 ( .B1(n1924), .B2(n3551), .A(n1916), .ZN(n4295) );
  OAI21_X1 U5903 ( .B1(n7510), .B2(n2377), .A(n4321), .ZN(n4320) );
  OAI221_X1 U5904 ( .B1(n2369), .B2(n1916), .C1(n7524), .C2(n1837), .A(n1917), 
        .ZN(Xfthu6) );
  AOI222_X1 U5905 ( .A1(n1918), .A2(n4670), .B1(n1919), .B2(n464), .C1(n1920), 
        .C2(n3690), .ZN(n2369) );
  OAI221_X1 U5906 ( .B1(n7535), .B2(n1858), .C1(n7369), .C2(n872), .A(n1862), 
        .ZN(n7980) );
  NAND2_X1 U5907 ( .A1(L6gpw6[23]), .A2(n866), .ZN(n1862) );
  AOI21_X1 U5908 ( .B1(n4191), .B2(n4192), .A(n2534), .ZN(D2phu6) );
  OAI22_X1 U5909 ( .A1(n8259), .A2(n2532), .B1(n672), .B2(n332), .ZN(n4192) );
  NAND2_X1 U5910 ( .A1(n6598), .A2(IRQ[14]), .ZN(n4191) );
  AOI21_X1 U5911 ( .B1(n3735), .B2(n3736), .A(n2683), .ZN(Jyohu6) );
  OAI22_X1 U5912 ( .A1(n2811), .A2(n2681), .B1(n672), .B2(n349), .ZN(n3736) );
  NAND2_X1 U5913 ( .A1(n6593), .A2(IRQ[30]), .ZN(n3735) );
  NAND3_X1 U5914 ( .A1(n3711), .A2(n8154), .A3(n3712), .ZN(n1891) );
  NAND3_X1 U5915 ( .A1(n8361), .A2(n8356), .A3(n7442), .ZN(n3711) );
  INV_X1 U5916 ( .A(STCLKEN), .ZN(n8361) );
  AOI21_X1 U5917 ( .B1(n4019), .B2(n4020), .A(n4021), .ZN(Ezohu6) );
  OAI22_X1 U5918 ( .A1(n8296), .A2(n4023), .B1(n672), .B2(n352), .ZN(n4020) );
  NAND2_X1 U5919 ( .A1(IRQ[27]), .A2(n6573), .ZN(n4019) );
  AOI22_X1 U5920 ( .A1(Gqgpw6[26]), .A2(n884), .B1(n1032), .B2(n883), .ZN(
        n1030) );
  OAI221_X1 U5921 ( .B1(n7488), .B2(n881), .C1(n7345), .C2(n2098), .A(n1089), 
        .ZN(n7897) );
  AOI22_X1 U5922 ( .A1(n883), .A2(n1090), .B1(ECOREVNUM[20]), .B2(n2002), .ZN(
        n1089) );
  NAND4_X1 U5923 ( .A1(n1091), .A2(n2136), .A3(n1093), .A4(n1094), .ZN(n1090)
         );
  AOI211_X1 U5924 ( .C1(n3475), .C2(Trgpw6[28]), .A(n1097), .B(n1098), .ZN(
        n1094) );
  AOI21_X1 U5925 ( .B1(n4197), .B2(n4198), .A(n2798), .ZN(Cyohu6) );
  OAI22_X1 U5926 ( .A1(n5192), .A2(n2796), .B1(n672), .B2(n356), .ZN(n4198) );
  NAND2_X1 U5927 ( .A1(n6591), .A2(IRQ[31]), .ZN(n4197) );
  OAI221_X1 U5928 ( .B1(n4764), .B2(n1020), .C1(n7291), .C2(n125), .A(n1186), 
        .ZN(n1178) );
  AOI22_X1 U5929 ( .A1(n2961), .A2(n3484), .B1(n1064), .B2(HRDATA[24]), .ZN(
        n1186) );
  AOI21_X1 U5930 ( .B1(n3738), .B2(n3739), .A(n2424), .ZN(Lzohu6) );
  OAI22_X1 U5931 ( .A1(n5154), .A2(n2422), .B1(n672), .B2(n344), .ZN(n3739) );
  NAND2_X1 U5932 ( .A1(n6602), .A2(IRQ[26]), .ZN(n3738) );
  AOI21_X1 U5933 ( .B1(n3754), .B2(n3755), .A(n3756), .ZN(Nwdpw6) );
  OAI22_X1 U5934 ( .A1(n3121), .A2(n3758), .B1(n672), .B2(n2632), .ZN(n3755)
         );
  NAND2_X1 U5935 ( .A1(IRQ[24]), .A2(n6580), .ZN(n3754) );
  OAI22_X1 U5936 ( .A1(n7533), .A2(N701), .B1(n2617), .B2(n963), .ZN(n7032) );
  OAI22_X1 U5937 ( .A1(n1889), .A2(n2979), .B1(n7530), .B2(n2980), .ZN(Oethu6)
         );
  NOR4_X1 U5938 ( .A1(n2981), .A2(n2982), .A3(n3707), .A4(n2984), .ZN(n2979)
         );
  AOI21_X1 U5939 ( .B1(n2501), .B2(n2495), .A(n1889), .ZN(n2980) );
  NOR3_X1 U5940 ( .A1(n2501), .A2(n2527), .A3(n3083), .ZN(n2984) );
  OAI22_X1 U5941 ( .A1(n7508), .A2(n451), .B1(n8301), .B2(n1997), .ZN(n8033)
         );
  INV_X1 U5942 ( .A(HRDATA[29]), .ZN(n8301) );
  OAI22_X1 U5943 ( .A1(n7509), .A2(n450), .B1(n8302), .B2(n1997), .ZN(n8032)
         );
  INV_X1 U5944 ( .A(HRDATA[28]), .ZN(n8302) );
  OAI22_X1 U5945 ( .A1(n7511), .A2(n1996), .B1(n8303), .B2(n1997), .ZN(n8031)
         );
  OAI22_X1 U5946 ( .A1(n7513), .A2(n451), .B1(n8304), .B2(n1997), .ZN(n8030)
         );
  OAI22_X1 U5947 ( .A1(n7515), .A2(n450), .B1(n8305), .B2(n1997), .ZN(n8029)
         );
  INV_X1 U5948 ( .A(HRDATA[25]), .ZN(n8305) );
  OAI22_X1 U5949 ( .A1(n7517), .A2(n1996), .B1(n8306), .B2(n1997), .ZN(n8028)
         );
  OAI22_X1 U5950 ( .A1(n1996), .A2(n4708), .B1(n8307), .B2(n1997), .ZN(n8027)
         );
  OAI22_X1 U5951 ( .A1(n7521), .A2(n451), .B1(n8308), .B2(n1997), .ZN(n8026)
         );
  OAI22_X1 U5952 ( .A1(n7522), .A2(n450), .B1(n8309), .B2(n1997), .ZN(n8025)
         );
  OAI22_X1 U5953 ( .A1(n7528), .A2(n1996), .B1(n8310), .B2(n1997), .ZN(n8024)
         );
  OAI22_X1 U5954 ( .A1(n451), .A2(n4702), .B1(n8311), .B2(n1997), .ZN(n8023)
         );
  AOI22_X1 U5955 ( .A1(ECOREVNUM[14]), .A2(n1074), .B1(ECOREVNUM[10]), .B2(
        n1075), .ZN(n1239) );
  NAND3_X1 U5956 ( .A1(n5476), .A2(n5477), .A3(n5478), .ZN(n888) );
  AOI221_X1 U5957 ( .B1(n2882), .B2(n8160), .C1(n2978), .C2(n4442), .A(n5486), 
        .ZN(n5477) );
  NOR4_X1 U5958 ( .A1(n5479), .A2(n5480), .A3(n5481), .A4(n5482), .ZN(n5478)
         );
  AOI221_X1 U5959 ( .B1(n2866), .B2(n2811), .C1(STCALIB[24]), .C2(n2973), .A(
        n4714), .ZN(n5476) );
  OAI22_X1 U5960 ( .A1(n7378), .A2(n1643), .B1(n2113), .B2(n4818), .ZN(n7023)
         );
  OAI211_X1 U5961 ( .C1(n705), .C2(n4700), .A(n707), .B(n708), .ZN(n7852) );
  AOI222_X1 U5962 ( .A1(n2131), .A2(n710), .B1(n711), .B2(n4841), .C1(n2118), 
        .C2(n4908), .ZN(n708) );
  AOI22_X1 U5963 ( .A1(n715), .A2(HRDATA[17]), .B1(n716), .B2(HRDATA[1]), .ZN(
        n707) );
  OAI211_X1 U5964 ( .C1(n705), .C2(n3673), .A(n1403), .B(n1404), .ZN(n7935) );
  AOI222_X1 U5965 ( .A1(n2118), .A2(n3690), .B1(n711), .B2(n2232), .C1(n2131), 
        .C2(n1407), .ZN(n1404) );
  AOI22_X1 U5966 ( .A1(n715), .A2(HRDATA[16]), .B1(n716), .B2(HRDATA[0]), .ZN(
        n1403) );
  OAI211_X1 U5967 ( .C1(n705), .C2(n4701), .A(n1373), .B(n1374), .ZN(n7924) );
  AOI222_X1 U5968 ( .A1(n2131), .A2(n119), .B1(n711), .B2(n3065), .C1(n2118), 
        .C2(n4910), .ZN(n1374) );
  AOI22_X1 U5969 ( .A1(n715), .A2(HRDATA[18]), .B1(n716), .B2(HRDATA[2]), .ZN(
        n1373) );
  OAI22_X1 U5970 ( .A1(n7491), .A2(N701), .B1(n961), .B2(n946), .ZN(n7207) );
  OAI22_X1 U5971 ( .A1(\sub_3151/A[0] ), .A2(n4818), .B1(n7497), .B2(n1643), 
        .ZN(n8017) );
  OAI22_X1 U5972 ( .A1(n7250), .A2(n2098), .B1(n856), .B2(n2393), .ZN(X3yhu6)
         );
  OAI22_X1 U5973 ( .A1(n7274), .A2(n1927), .B1(n2448), .B2(n2408), .ZN(Vxohu6)
         );
  AOI211_X1 U5974 ( .C1(n82), .C2(n4506), .A(n2450), .B(n2599), .ZN(n2448) );
  INV_X1 U5975 ( .A(n2414), .ZN(n2599) );
  OAI211_X1 U5976 ( .C1(n7259), .C2(n2275), .A(n2452), .B(n2453), .ZN(n2450)
         );
  AND2_X1 U5977 ( .A1(Ntkbx6[8]), .A2(n2695), .ZN(S6ihu6) );
  OAI22_X1 U5978 ( .A1(n697), .A2(n1774), .B1(n696), .B2(n4810), .ZN(n2695) );
  AOI22_X1 U5979 ( .A1(ECOREVNUM[6]), .A2(n1066), .B1(n3476), .B2(E1hpw6[6]), 
        .ZN(n1238) );
  OAI22_X1 U5980 ( .A1(n1808), .A2(n1979), .B1(n7626), .B2(n409), .ZN(Lirhu6)
         );
  OAI22_X1 U5981 ( .A1(n7387), .A2(n890), .B1(n6906), .B2(n719), .ZN(Zcxhu6)
         );
  OAI22_X1 U5982 ( .A1(n7437), .A2(n890), .B1(n6766), .B2(n885), .ZN(Gdxhu6)
         );
  OAI22_X1 U5983 ( .A1(n7430), .A2(n890), .B1(n6727), .B2(n885), .ZN(M9xhu6)
         );
  NAND2_X1 U5984 ( .A1(n8291), .A2(n6403), .ZN(n6154) );
  NAND3_X1 U5985 ( .A1(n6404), .A2(n2227), .A3(n6681), .ZN(n6403) );
  OAI21_X1 U5986 ( .B1(n7615), .B2(n3785), .A(n6405), .ZN(n6404) );
  OAI211_X1 U5987 ( .C1(n7434), .C2(n4454), .A(n4459), .B(n7679), .ZN(n6405)
         );
  OAI22_X1 U5988 ( .A1(n7657), .A2(n890), .B1(n6692), .B2(n885), .ZN(Aaxhu6)
         );
  OAI22_X1 U5989 ( .A1(n7667), .A2(n890), .B1(n6741), .B2(n885), .ZN(Jbxhu6)
         );
  OAI22_X1 U5990 ( .A1(n7428), .A2(n890), .B1(n6904), .B2(n885), .ZN(Ecxhu6)
         );
  OAI22_X1 U5991 ( .A1(n7397), .A2(n890), .B1(n6750), .B2(n719), .ZN(Pexhu6)
         );
  OAI22_X1 U5992 ( .A1(n7661), .A2(n890), .B1(n6718), .B2(n719), .ZN(Xbxhu6)
         );
  OAI22_X1 U5993 ( .A1(n7648), .A2(n890), .B1(n6905), .B2(n719), .ZN(Scxhu6)
         );
  AOI21_X1 U5994 ( .B1(n7283), .B2(n961), .A(n2554), .ZN(Twohu6) );
  AND4_X1 U5995 ( .A1(n2555), .A2(n2556), .A3(n2557), .A4(n2558), .ZN(n2554)
         );
  AOI221_X1 U5996 ( .B1(n1945), .B2(n529), .C1(n1761), .C2(n1482), .A(n2573), 
        .ZN(n2556) );
  NOR4_X1 U5997 ( .A1(n2559), .A2(n1737), .A3(n2560), .A4(n1653), .ZN(n2558)
         );
  OAI22_X1 U5998 ( .A1(n7488), .A2(n890), .B1(n6882), .B2(n719), .ZN(T9xhu6)
         );
  OAI22_X1 U5999 ( .A1(n7429), .A2(n890), .B1(n6894), .B2(n719), .ZN(Vaxhu6)
         );
  OAI22_X1 U6000 ( .A1(n7410), .A2(n890), .B1(n6897), .B2(n885), .ZN(F9xhu6)
         );
  OAI22_X1 U6001 ( .A1(n7664), .A2(n890), .B1(n6907), .B2(n719), .ZN(Qbxhu6)
         );
  OAI22_X1 U6002 ( .A1(n7681), .A2(n890), .B1(n6912), .B2(n885), .ZN(Cbxhu6)
         );
  OAI22_X1 U6003 ( .A1(n7427), .A2(n890), .B1(n6903), .B2(n885), .ZN(Lcxhu6)
         );
  OAI22_X1 U6004 ( .A1(n7655), .A2(n890), .B1(n7653), .B2(n885), .ZN(Haxhu6)
         );
  NAND3_X1 U6005 ( .A1(n4768), .A2(n4769), .A3(n4770), .ZN(n1149) );
  AOI22_X1 U6006 ( .A1(n2866), .A2(n3276), .B1(n2852), .B2(n8134), .ZN(n4768)
         );
  AOI221_X1 U6007 ( .B1(n2976), .B2(Tzfpw6[1]), .C1(STCALIB[1]), .C2(n2973), 
        .A(n4771), .ZN(n4770) );
  AOI222_X1 U6008 ( .A1(n2201), .A2(n4491), .B1(n2998), .B2(n8155), .C1(
        ECOREVNUM[1]), .C2(n4714), .ZN(n4769) );
  OAI22_X1 U6009 ( .A1(n7693), .A2(n890), .B1(n6915), .B2(n719), .ZN(Oaxhu6)
         );
  OAI22_X1 U6010 ( .A1(n7487), .A2(n890), .B1(n6884), .B2(n719), .ZN(O2yhu6)
         );
  OAI22_X1 U6011 ( .A1(n7641), .A2(n890), .B1(n6708), .B2(n885), .ZN(Ndxhu6)
         );
  OAI22_X1 U6012 ( .A1(n7631), .A2(n890), .B1(n6756), .B2(n885), .ZN(Iexhu6)
         );
  OAI22_X1 U6013 ( .A1(n7447), .A2(n890), .B1(n6908), .B2(n719), .ZN(Udxhu6)
         );
  OAI211_X1 U6014 ( .C1(n7354), .C2(n1376), .A(n1424), .B(n1425), .ZN(n7939)
         );
  AOI22_X1 U6015 ( .A1(n711), .A2(n3533), .B1(n1412), .B2(n797), .ZN(n1424) );
  AOI221_X1 U6016 ( .B1(n1410), .B2(n1426), .C1(n2119), .C2(n4699), .A(n2131), 
        .ZN(n1425) );
  OAI22_X1 U6017 ( .A1(n7450), .A2(n890), .B1(n6875), .B2(n885), .ZN(Bexhu6)
         );
  OAI22_X1 U6018 ( .A1(n1811), .A2(n1979), .B1(n7703), .B2(n409), .ZN(Levhu6)
         );
  AOI21_X1 U6019 ( .B1(Gqgpw6[11]), .B2(n884), .A(n877), .ZN(n1196) );
  OAI22_X1 U6020 ( .A1(n7375), .A2(N701), .B1(n1437), .B2(n961), .ZN(n7941) );
  AND4_X1 U6021 ( .A1(n1438), .A2(n1439), .A3(n1440), .A4(n1441), .ZN(n1437)
         );
  AOI221_X1 U6022 ( .B1(n474), .B2(n1539), .C1(n1540), .C2(n7283), .A(n1541), 
        .ZN(n1438) );
  AOI211_X1 U6023 ( .C1(n1442), .C2(n1443), .A(n1444), .B(n1445), .ZN(n1441)
         );
  NAND3_X1 U6024 ( .A1(n4709), .A2(n4710), .A3(n4711), .ZN(n1343) );
  AOI22_X1 U6025 ( .A1(n2866), .A2(n3030), .B1(n2852), .B2(n8142), .ZN(n4709)
         );
  AOI221_X1 U6026 ( .B1(n2976), .B2(Tzfpw6[2]), .C1(STCALIB[2]), .C2(n2973), 
        .A(n4712), .ZN(n4711) );
  AOI221_X1 U6027 ( .B1(n2201), .B2(n8133), .C1(ECOREVNUM[2]), .C2(n4714), .A(
        n4715), .ZN(n4710) );
  AOI21_X1 U6028 ( .B1(n7442), .B2(n8356), .A(n1894), .ZN(n4715) );
  AOI21_X1 U6029 ( .B1(n1204), .B2(n883), .A(n877), .ZN(n1203) );
  OAI21_X1 U6030 ( .B1(n991), .B2(n6743), .A(n2832), .ZN(n1204) );
  AOI21_X1 U6031 ( .B1(n1299), .B2(n883), .A(n877), .ZN(n1298) );
  OR4_X1 U6032 ( .A1(n1300), .A2(n1301), .A3(n3397), .A4(n1302), .ZN(n1299) );
  OAI21_X1 U6033 ( .B1(n1000), .B2(n2227), .A(n1313), .ZN(n1301) );
  OAI221_X1 U6034 ( .B1(n7460), .B2(n1005), .C1(n6645), .C2(n1008), .A(n3456), 
        .ZN(n1300) );
  OAI22_X1 U6035 ( .A1(n7284), .A2(n3022), .B1(n3070), .B2(n1913), .ZN(Mwohu6)
         );
  NOR2_X1 U6036 ( .A1(n3071), .A2(n2270), .ZN(n3070) );
  OAI221_X1 U6037 ( .B1(n7393), .B2(n3029), .C1(n7516), .C2(n3028), .A(n3076), 
        .ZN(n3071) );
  INV_X1 U6038 ( .A(n3073), .ZN(n2270) );
  OAI221_X1 U6039 ( .B1(n7423), .B2(n881), .C1(n7640), .C2(n2098), .A(n1051), 
        .ZN(n7895) );
  AOI21_X1 U6040 ( .B1(n883), .B2(n1052), .A(n2002), .ZN(n1051) );
  NAND4_X1 U6041 ( .A1(n1053), .A2(n1054), .A3(n1055), .A4(n1056), .ZN(n1052)
         );
  AOI22_X1 U6042 ( .A1(ECOREVNUM[13]), .A2(n1074), .B1(ECOREVNUM[9]), .B2(
        n1075), .ZN(n1053) );
  NOR2_X1 U6043 ( .A1(n4012), .A2(n2672), .ZN(F3phu6) );
  AOI21_X1 U6044 ( .B1(n6594), .B2(IRQ[10]), .A(n4014), .ZN(n4012) );
  AOI22_X1 U6045 ( .A1(HWDATA[10]), .A2(n226), .B1(n2669), .B2(n7584), .ZN(
        n4014) );
  OAI22_X1 U6046 ( .A1(n7343), .A2(n3022), .B1(n3023), .B2(n1913), .ZN(Ntohu6)
         );
  AOI211_X1 U6047 ( .C1(n3025), .C2(n3690), .A(n3026), .B(n3027), .ZN(n3023)
         );
  OAI22_X1 U6048 ( .A1(n7518), .A2(n3028), .B1(n7259), .B2(n3029), .ZN(n3026)
         );
  INV_X1 U6049 ( .A(n1953), .ZN(n1855) );
  AOI22_X1 U6050 ( .A1(n1954), .A2(SLEEPHOLDACKn), .B1(SLEEPHOLDREQn), .B2(
        N701), .ZN(n1953) );
  OAI211_X1 U6051 ( .C1(n2519), .C2(n3786), .A(n1955), .B(n1956), .ZN(n1954)
         );
  NOR2_X1 U6052 ( .A1(n878), .A2(n1960), .ZN(n1955) );
  OAI22_X1 U6053 ( .A1(n7332), .A2(N701), .B1(n1928), .B2(n961), .ZN(n8007) );
  NOR4_X1 U6054 ( .A1(n1929), .A2(n1930), .A3(n1931), .A4(n1932), .ZN(n1928)
         );
  OAI221_X1 U6055 ( .B1(n1933), .B2(n3860), .C1(n2529), .C2(n3737), .A(n1935), 
        .ZN(n1930) );
  OAI221_X1 U6056 ( .B1(n1940), .B2(n4265), .C1(n1941), .C2(n1518), .A(n1942), 
        .ZN(n1929) );
  OAI21_X1 U6057 ( .B1(n7532), .B2(N701), .A(n2120), .ZN(n7027) );
  OAI211_X1 U6058 ( .C1(n2511), .C2(n5284), .A(n1978), .B(N701), .ZN(n2120) );
  OAI21_X1 U6059 ( .B1(n1982), .B2(n4546), .A(n1983), .ZN(n8015) );
  OAI211_X1 U6060 ( .C1(n1984), .C2(n1985), .A(n4512), .B(n1643), .ZN(n1983)
         );
  NOR2_X1 U6061 ( .A1(n7378), .A2(n7533), .ZN(n1985) );
  AND3_X1 U6062 ( .A1(n7533), .A2(n3952), .A3(n3765), .ZN(n1984) );
  AND2_X1 U6063 ( .A1(Nvkbx6[8]), .A2(n3949), .ZN(Gqkhu6) );
  OAI22_X1 U6064 ( .A1(n2264), .A2(n4810), .B1(n736), .B2(n1774), .ZN(n3949)
         );
  NAND3_X1 U6065 ( .A1(n1966), .A2(n1840), .A3(EDBGRQ), .ZN(n1961) );
  OAI22_X1 U6066 ( .A1(n1889), .A2(n3227), .B1(n7326), .B2(n3228), .ZN(L7vhu6)
         );
  NOR4_X1 U6067 ( .A1(n3229), .A2(n3230), .A3(n3707), .A4(n3231), .ZN(n3227)
         );
  AOI21_X1 U6068 ( .B1(n7529), .B2(n2495), .A(n1889), .ZN(n3228) );
  NOR3_X1 U6069 ( .A1(n5294), .A2(n7529), .A3(n2527), .ZN(n3231) );
  OAI22_X1 U6070 ( .A1(n2658), .A2(n1694), .B1(n7356), .B2(n2659), .ZN(Ssohu6)
         );
  AOI221_X1 U6071 ( .B1(n1697), .B2(n4987), .C1(n1698), .C2(n470), .A(n2661), 
        .ZN(n2658) );
  AOI21_X1 U6072 ( .B1(n1705), .B2(n3566), .A(n1694), .ZN(n2659) );
  OAI22_X1 U6073 ( .A1(n7393), .A2(n1701), .B1(n7495), .B2(n1700), .ZN(n2661)
         );
  OAI22_X1 U6074 ( .A1(n7506), .A2(n3093), .B1(n3094), .B2(n1694), .ZN(Miohu6)
         );
  AOI22_X1 U6075 ( .A1(n3095), .A2(n4670), .B1(n2258), .B2(n4993), .ZN(n3094)
         );
  AOI21_X1 U6076 ( .B1(n1705), .B2(n3099), .A(n1694), .ZN(n3093) );
  NAND2_X1 U6077 ( .A1(n3097), .A2(n3098), .ZN(n3095) );
  OAI22_X1 U6078 ( .A1(n7527), .A2(n3206), .B1(n3207), .B2(n1694), .ZN(Leohu6)
         );
  AOI22_X1 U6079 ( .A1(n2258), .A2(n4987), .B1(n1697), .B2(n4993), .ZN(n3207)
         );
  AOI21_X1 U6080 ( .B1(n1705), .B2(n3554), .A(n1694), .ZN(n3206) );
  INV_X1 U6081 ( .A(n2807), .ZN(n3554) );
  OAI211_X1 U6082 ( .C1(n1173), .C2(n741), .A(n1166), .B(n1174), .ZN(n7903) );
  NOR4_X1 U6083 ( .A1(n1176), .A2(n1177), .A3(n1178), .A4(n1179), .ZN(n1173)
         );
  AOI22_X1 U6084 ( .A1(n239), .A2(n3389), .B1(n6654), .B2(n856), .ZN(n1174) );
  OAI221_X1 U6085 ( .B1(n6836), .B2(n991), .C1(n6853), .C2(n990), .A(n3468), 
        .ZN(n1176) );
  OAI221_X1 U6086 ( .B1(n3115), .B2(n180), .C1(n397), .C2(n1832), .A(n465), 
        .ZN(n7828) );
  AOI222_X1 U6087 ( .A1(n241), .A2(n466), .B1(n467), .B2(n258), .C1(n182), 
        .C2(vis_ipsr_o[0]), .ZN(n465) );
  OAI21_X1 U6088 ( .B1(n1849), .B2(n3486), .A(n478), .ZN(n467) );
  NAND3_X1 U6089 ( .A1(n259), .A2(n180), .A3(vis_primask_o), .ZN(n478) );
  OAI22_X1 U6090 ( .A1(n7529), .A2(n2480), .B1(n1889), .B2(n2837), .ZN(Pgvhu6)
         );
  NOR2_X1 U6091 ( .A1(n2838), .A2(n2839), .ZN(n2837) );
  OAI221_X1 U6092 ( .B1(n7359), .B2(n2254), .C1(n485), .C2(n2524), .A(n2841), 
        .ZN(n2839) );
  NAND4_X1 U6093 ( .A1(n2603), .A2(n3805), .A3(n2843), .A4(n2844), .ZN(n2838)
         );
  OAI22_X1 U6094 ( .A1(n7520), .A2(n3022), .B1(n3964), .B2(n1913), .ZN(Gfohu6)
         );
  AOI21_X1 U6095 ( .B1(n3965), .B2(n4670), .A(n3027), .ZN(n3964) );
  OAI21_X1 U6096 ( .B1(n7514), .B2(n3966), .A(n3761), .ZN(n3965) );
  NAND3_X1 U6097 ( .A1(n3085), .A2(n5916), .A3(n5917), .ZN(n5903) );
  NAND4_X1 U6098 ( .A1(n3712), .A2(n7530), .A3(n4458), .A4(n5070), .ZN(n5917)
         );
  NAND4_X1 U6099 ( .A1(n52), .A2(n80), .A3(n5918), .A4(n272), .ZN(n5916) );
  INV_X1 U6100 ( .A(n4464), .ZN(n3085) );
  OAI22_X1 U6101 ( .A1(n7360), .A2(n1927), .B1(n3160), .B2(n2408), .ZN(Lsohu6)
         );
  AOI211_X1 U6102 ( .C1(n1751), .C2(n3690), .A(n3161), .B(n3162), .ZN(n3160)
         );
  OAI221_X1 U6103 ( .B1(n7505), .B2(n2256), .C1(n7524), .C2(n2572), .A(n2414), 
        .ZN(n3161) );
  OAI22_X1 U6104 ( .A1(n7259), .A2(n2412), .B1(n3163), .B2(n2515), .ZN(n3162)
         );
  OAI22_X1 U6105 ( .A1(n7394), .A2(n1927), .B1(n2801), .B2(n2408), .ZN(Q4xhu6)
         );
  NOR4_X1 U6106 ( .A1(n2802), .A2(n2803), .A3(n1563), .A4(n2804), .ZN(n2801)
         );
  OAI22_X1 U6107 ( .A1(n7325), .A2(n2275), .B1(n7393), .B2(n2412), .ZN(n2803)
         );
  NOR2_X1 U6108 ( .A1(n2805), .A2(n2515), .ZN(n2804) );
  OAI22_X1 U6109 ( .A1(n7330), .A2(n1927), .B1(n2407), .B2(n2408), .ZN(Wuohu6)
         );
  AOI211_X1 U6110 ( .C1(n1684), .C2(n464), .A(n2409), .B(n2410), .ZN(n2407) );
  OAI22_X1 U6112 ( .A1(n7329), .A2(n2275), .B1(n7523), .B2(n2412), .ZN(n2410)
         );
  OAI221_X1 U6113 ( .B1(n1706), .B2(n2515), .C1(n7526), .C2(n2572), .A(n2414), 
        .ZN(n2409) );
  OAI21_X1 U6114 ( .B1(n7507), .B2(N701), .A(n1989), .ZN(n7026) );
  NAND2_X1 U6115 ( .A1(n7380), .A2(n3505), .ZN(n797) );
  OAI22_X1 U6116 ( .A1(n7493), .A2(N701), .B1(n2553), .B2(n1976), .ZN(n8013)
         );
  INV_X1 U6117 ( .A(n1978), .ZN(n2553) );
  AOI21_X1 U6118 ( .B1(n1430), .B2(N701), .A(n1977), .ZN(n1976) );
  OAI22_X1 U6119 ( .A1(n6770), .A2(n1996), .B1(n3488), .B2(n4695), .ZN(n7025)
         );
  NOR3_X1 U6120 ( .A1(n2531), .A2(n2532), .A3(n8344), .ZN(Uothu6) );
  OAI221_X1 U6121 ( .B1(n2534), .B2(n8258), .C1(n234), .C2(n2536), .A(n897), 
        .ZN(n2531) );
  INV_X1 U6122 ( .A(IRQ[14]), .ZN(n8344) );
  NOR3_X1 U6123 ( .A1(n2795), .A2(n2796), .A3(n8330), .ZN(Q6vhu6) );
  OAI221_X1 U6124 ( .B1(n2798), .B2(n5180), .C1(n234), .C2(n2800), .A(n897), 
        .ZN(n2795) );
  INV_X1 U6125 ( .A(IRQ[31]), .ZN(n8330) );
  NOR3_X1 U6126 ( .A1(n2680), .A2(n2681), .A3(n8331), .ZN(Sgthu6) );
  OAI221_X1 U6127 ( .B1(n2683), .B2(n5175), .C1(n234), .C2(n2685), .A(n897), 
        .ZN(n2680) );
  INV_X1 U6128 ( .A(IRQ[30]), .ZN(n8331) );
  NOR3_X1 U6129 ( .A1(n2421), .A2(n2422), .A3(n8334), .ZN(Wpthu6) );
  OAI221_X1 U6130 ( .B1(n2424), .B2(n5148), .C1(n234), .C2(n2426), .A(n897), 
        .ZN(n2421) );
  INV_X1 U6131 ( .A(IRQ[26]), .ZN(n8334) );
  OAI22_X1 U6132 ( .A1(n7286), .A2(n2480), .B1(n1889), .B2(n2482), .ZN(Vethu6)
         );
  NOR2_X1 U6133 ( .A1(n2483), .A2(n2484), .ZN(n2482) );
  OAI221_X1 U6134 ( .B1(n4725), .B2(n2250), .C1(n265), .C2(n4633), .A(n2487), 
        .ZN(n2484) );
  OAI221_X1 U6135 ( .B1(n2272), .B2(n2491), .C1(n7329), .C2(n2492), .A(n2493), 
        .ZN(n2483) );
  OAI22_X1 U6136 ( .A1(n7382), .A2(n3022), .B1(n5020), .B2(n1913), .ZN(Aqohu6)
         );
  AOI211_X1 U6137 ( .C1(n3025), .C2(n4910), .A(n5021), .B(n3027), .ZN(n5020)
         );
  OAI22_X1 U6138 ( .A1(n7514), .A2(n3028), .B1(n7523), .B2(n3029), .ZN(n5021)
         );
  OAI22_X1 U6139 ( .A1(n6768), .A2(N701), .B1(n2114), .B2(n2115), .ZN(n7024)
         );
  OAI221_X1 U6140 ( .B1(n2117), .B2(n254), .C1(n7355), .C2(n508), .A(n272), 
        .ZN(n2114) );
  NAND2_X1 U6141 ( .A1(n2116), .A2(N701), .ZN(n2115) );
  NOR3_X1 U6142 ( .A1(n503), .A2(n4512), .A3(n2572), .ZN(n2117) );
  OAI22_X1 U6143 ( .A1(n3084), .A2(n4364), .B1(n4455), .B2(n4456), .ZN(Brrhu6)
         );
  AOI22_X1 U6144 ( .A1(n4457), .A2(n4458), .B1(vis_pc_o[1]), .B2(n4753), .ZN(
        n4455) );
  INV_X1 U6145 ( .A(n4456), .ZN(n3084) );
  NAND2_X1 U6146 ( .A1(N701), .A2(n4461), .ZN(n4456) );
  NOR2_X1 U6147 ( .A1(n3750), .A2(n3751), .ZN(R2phu6) );
  AOI21_X1 U6148 ( .B1(IRQ[12]), .B2(n6579), .A(n3752), .ZN(n3750) );
  AOI22_X1 U6149 ( .A1(HWDATA[12]), .A2(n226), .B1(n3753), .B2(n7583), .ZN(
        n3752) );
  NOR2_X1 U6150 ( .A1(n3578), .A2(n2245), .ZN(Y2phu6) );
  AOI21_X1 U6151 ( .B1(n6606), .B2(IRQ[11]), .A(n3580), .ZN(n3578) );
  AOI22_X1 U6152 ( .A1(HWDATA[11]), .A2(n226), .B1(n2241), .B2(n7585), .ZN(
        n3580) );
  AND2_X1 U6153 ( .A1(Ntkbx6[6]), .A2(n4403), .ZN(C4ihu6) );
  OAI22_X1 U6154 ( .A1(n701), .A2(n1785), .B1(n2297), .B2(n4816), .ZN(n4403)
         );
  AND2_X1 U6155 ( .A1(Nvkbx6[6]), .A2(n2780), .ZN(Qnkhu6) );
  OAI22_X1 U6156 ( .A1(n2264), .A2(n4816), .B1(n734), .B2(n1785), .ZN(n2780)
         );
  NOR2_X1 U6157 ( .A1(n3741), .A2(n3038), .ZN(K2phu6) );
  AOI21_X1 U6158 ( .B1(n6587), .B2(IRQ[13]), .A(n3743), .ZN(n3741) );
  AOI22_X1 U6159 ( .A1(HWDATA[13]), .A2(n226), .B1(n3035), .B2(n7586), .ZN(
        n3743) );
  NOR2_X1 U6160 ( .A1(n3613), .A2(n2476), .ZN(n7271) );
  INV_X1 U6161 ( .A(n3615), .ZN(n2476) );
  OAI221_X1 U6162 ( .B1(n7357), .B2(n3616), .C1(n8343), .C2(n8249), .A(n3619), 
        .ZN(n3615) );
  NOR2_X1 U6163 ( .A1(n1835), .A2(n672), .ZN(n3616) );
  OAI21_X1 U6164 ( .B1(DBGRESTART), .B2(n963), .A(n1965), .ZN(n8010) );
  OAI21_X1 U6165 ( .B1(n963), .B2(n1966), .A(DBGRESTARTED), .ZN(n1965) );
  NAND2_X1 U6166 ( .A1(n6475), .A2(n6476), .ZN(n1267) );
  AOI221_X1 U6167 ( .B1(n2201), .B2(n4535), .C1(n2866), .C2(n5197), .A(n6477), 
        .ZN(n6476) );
  AOI222_X1 U6168 ( .A1(STCALIB[4]), .A2(n2973), .B1(n2975), .B2(n4545), .C1(
        n2976), .C2(Tzfpw6[4]), .ZN(n6475) );
  OAI22_X1 U6169 ( .A1(n5105), .A2(n2825), .B1(n7685), .B2(n4729), .ZN(n6477)
         );
  OAI21_X1 U6170 ( .B1(n7400), .B2(n1689), .A(n1690), .ZN(n7945) );
  AOI21_X1 U6171 ( .B1(n1705), .B2(n1706), .A(n1694), .ZN(n1689) );
  OAI21_X1 U6172 ( .B1(n1691), .B2(n2238), .A(n1885), .ZN(n1690) );
  OAI221_X1 U6173 ( .B1(n7494), .B2(n1700), .C1(n7259), .C2(n1701), .A(n1702), 
        .ZN(n1691) );
  OAI21_X1 U6174 ( .B1(n3569), .B2(n3570), .A(n4535), .ZN(n3567) );
  NAND4_X1 U6175 ( .A1(n3572), .A2(n3573), .A3(n3574), .A4(n3575), .ZN(n3570)
         );
  NAND4_X1 U6176 ( .A1(n3678), .A2(n3679), .A3(n3680), .A4(n3681), .ZN(n3569)
         );
  AOI221_X1 U6177 ( .B1(n7260), .B2(n7593), .C1(n7254), .C2(n7592), .A(n2682), 
        .ZN(n3572) );
  NAND2_X1 U6178 ( .A1(n5665), .A2(n5666), .ZN(n1302) );
  AOI211_X1 U6179 ( .C1(ECOREVNUM[3]), .C2(n4714), .A(n5667), .B(n4781), .ZN(
        n5666) );
  AOI221_X1 U6180 ( .B1(n2976), .B2(Tzfpw6[3]), .C1(STCALIB[3]), .C2(n2973), 
        .A(n5670), .ZN(n5665) );
  OAI22_X1 U6181 ( .A1(n7690), .A2(n4729), .B1(n7689), .B2(n4730), .ZN(n5667)
         );
  OAI21_X1 U6182 ( .B1(n3559), .B2(n2502), .A(n3560), .ZN(J4xhu6) );
  OAI21_X1 U6183 ( .B1(n2519), .B2(n1959), .A(n2502), .ZN(n3560) );
  NOR4_X1 U6184 ( .A1(n3564), .A2(n3565), .A3(RXEV), .A4(TXEV), .ZN(n3559) );
  NAND3_X1 U6185 ( .A1(n3567), .A2(n3568), .A3(n3712), .ZN(n3564) );
  NAND2_X1 U6186 ( .A1(n5396), .A2(n5397), .ZN(n997) );
  AOI221_X1 U6187 ( .B1(n2976), .B2(Tzfpw6[0]), .C1(STCALIB[0]), .C2(n2973), 
        .A(n5399), .ZN(n5396) );
  AOI221_X1 U6188 ( .B1(n2998), .B2(n8154), .C1(ECOREVNUM[0]), .C2(n4714), .A(
        n5398), .ZN(n5397) );
  OAI22_X1 U6189 ( .A1(n7351), .A2(n2202), .B1(n5112), .B2(n2825), .ZN(n5399)
         );
  NAND2_X1 U6190 ( .A1(n4778), .A2(n4779), .ZN(n1213) );
  AOI211_X1 U6191 ( .C1(n2866), .C2(n3930), .A(n4780), .B(n4781), .ZN(n4779)
         );
  AOI221_X1 U6192 ( .B1(n2976), .B2(Tzfpw6[9]), .C1(STCALIB[9]), .C2(n2973), 
        .A(n4714), .ZN(n4778) );
  OAI22_X1 U6193 ( .A1(n7698), .A2(n2202), .B1(n7697), .B2(n4729), .ZN(n4780)
         );
  OAI211_X1 U6194 ( .C1(n7292), .C2(n2098), .A(n970), .B(n971), .ZN(n7890) );
  AOI222_X1 U6195 ( .A1(n239), .A2(Tnhpw6[0]), .B1(n883), .B2(n973), .C1(n2004), .C2(n4142), .ZN(n971) );
  NAND4_X1 U6196 ( .A1(n1822), .A2(n3453), .A3(n978), .A4(n979), .ZN(n973) );
  INV_X1 U6197 ( .A(n1003), .ZN(n3453) );
  INV_X1 U6198 ( .A(HRDATA[18]), .ZN(n8312) );
  NAND2_X1 U6199 ( .A1(n7392), .A2(n3505), .ZN(n1426) );
  INV_X1 U6200 ( .A(HRDATA[4]), .ZN(n8325) );
  INV_X1 U6201 ( .A(HRDATA[2]), .ZN(n8327) );
  INV_X1 U6202 ( .A(HRDATA[20]), .ZN(n8310) );
  INV_X1 U6203 ( .A(HRDATA[0]), .ZN(n8329) );
  INV_X1 U6204 ( .A(HRDATA[19]), .ZN(n8311) );
  INV_X1 U6205 ( .A(HRDATA[23]), .ZN(n8307) );
  INV_X1 U6206 ( .A(HRDATA[16]), .ZN(n8314) );
  INV_X1 U6207 ( .A(HRDATA[11]), .ZN(n8318) );
  INV_X1 U6208 ( .A(HRDATA[9]), .ZN(n8320) );
  INV_X1 U6209 ( .A(n4696), .ZN(n2832) );
  OAI211_X1 U6210 ( .C1(n7365), .C2(n2202), .A(n4697), .B(n4698), .ZN(n4696)
         );
  AOI22_X1 U6211 ( .A1(n2866), .A2(n8170), .B1(n2852), .B2(n8169), .ZN(n4697)
         );
  AOI22_X1 U6212 ( .A1(n2976), .A2(Tzfpw6[10]), .B1(STCALIB[10]), .B2(n2973), 
        .ZN(n4698) );
  INV_X1 U6213 ( .A(n5686), .ZN(n2827) );
  OAI211_X1 U6214 ( .C1(n7379), .C2(n2202), .A(n5687), .B(n5688), .ZN(n5686)
         );
  AOI22_X1 U6215 ( .A1(n2866), .A2(n3870), .B1(n2852), .B2(n8143), .ZN(n5687)
         );
  AOI221_X1 U6216 ( .B1(n2976), .B2(Tzfpw6[19]), .C1(STCALIB[19]), .C2(n2973), 
        .A(n4714), .ZN(n5688) );
  INV_X1 U6217 ( .A(n5679), .ZN(n2835) );
  OAI211_X1 U6218 ( .C1(n7327), .C2(n2202), .A(n5680), .B(n5681), .ZN(n5679)
         );
  AOI22_X1 U6219 ( .A1(n2866), .A2(n8166), .B1(n2852), .B2(n8165), .ZN(n5680)
         );
  AOI22_X1 U6220 ( .A1(n2976), .A2(Tzfpw6[11]), .B1(STCALIB[11]), .B2(n2973), 
        .ZN(n5681) );
  INV_X1 U6221 ( .A(n6077), .ZN(n2840) );
  OAI211_X1 U6222 ( .C1(n7277), .C2(n2202), .A(n6078), .B(n6079), .ZN(n6077)
         );
  AOI22_X1 U6223 ( .A1(n2866), .A2(n8227), .B1(n2852), .B2(n8225), .ZN(n6078)
         );
  AOI22_X1 U6224 ( .A1(n2976), .A2(Tzfpw6[20]), .B1(STCALIB[20]), .B2(n2973), 
        .ZN(n6079) );
  NOR3_X1 U6225 ( .A1(n1242), .A2(n2855), .A3(n1244), .ZN(n1241) );
  OAI21_X1 U6226 ( .B1(n4816), .B2(n1020), .A(n3443), .ZN(n1244) );
  OAI221_X1 U6227 ( .B1(n6808), .B2(n989), .C1(n6861), .C2(n985), .A(n3450), 
        .ZN(n1242) );
  INV_X1 U6228 ( .A(n1251), .ZN(n2855) );
  INV_X1 U6229 ( .A(n5330), .ZN(n2833) );
  OAI211_X1 U6230 ( .C1(n7289), .C2(n2202), .A(n5331), .B(n5332), .ZN(n5330)
         );
  AOI22_X1 U6231 ( .A1(n2866), .A2(n3669), .B1(n2852), .B2(n8148), .ZN(n5331)
         );
  AOI22_X1 U6232 ( .A1(n2976), .A2(Tzfpw6[21]), .B1(STCALIB[21]), .B2(n2973), 
        .ZN(n5332) );
  AND4_X1 U6233 ( .A1(n7488), .A2(n3880), .A3(n8206), .A4(n4151), .ZN(n3850)
         );
  NAND2_X1 U6234 ( .A1(HRESP), .A2(n4152), .ZN(n2393) );
  INV_X1 U6235 ( .A(n5344), .ZN(n2826) );
  AOI211_X1 U6236 ( .C1(vis_ipsr_o[5]), .C2(n5345), .A(n5346), .B(n5347), .ZN(
        n5344) );
  OAI22_X1 U6237 ( .A1(n4730), .A2(n3645), .B1(n4729), .B2(n7572), .ZN(n5346)
         );
  OAI222_X1 U6238 ( .A1(n8360), .A2(n4788), .B1(n2202), .B2(n7338), .C1(n1893), 
        .C2(n7339), .ZN(n5347) );
  AND3_X1 U6239 ( .A1(n4401), .A2(n7401), .A3(n4748), .ZN(n403) );
  OAI21_X1 U6240 ( .B1(n911), .B2(n909), .A(n912), .ZN(n7883) );
  OR3_X1 U6241 ( .A1(n2102), .A2(n7412), .A3(n914), .ZN(n912) );
  NAND3_X1 U6242 ( .A1(n1895), .A2(n1896), .A3(n1897), .ZN(n8004) );
  OAI21_X1 U6243 ( .B1(n1505), .B2(n963), .A(n479), .ZN(n1895) );
  OAI21_X1 U6244 ( .B1(n1898), .B2(n1899), .A(N701), .ZN(n1897) );
  NAND3_X1 U6245 ( .A1(n7375), .A2(n7492), .A3(n1643), .ZN(n1896) );
  AOI221_X1 U6246 ( .B1(K2phu6), .B2(n7586), .C1(Lzohu6), .C2(n6581), .A(n2645), .ZN(n3679) );
  INV_X1 U6247 ( .A(n3734), .ZN(n2645) );
  AOI222_X1 U6248 ( .A1(n7684), .A2(H4phu6), .B1(n7595), .B2(n2646), .C1(n7255), .C2(Jyohu6), .ZN(n3734) );
  AOI221_X1 U6249 ( .B1(n7265), .B2(n7588), .C1(n7264), .C2(n7590), .A(n1828), 
        .ZN(n3573) );
  INV_X1 U6250 ( .A(n3626), .ZN(n1828) );
  AOI222_X1 U6251 ( .A1(n7589), .A2(n7267), .B1(n6575), .B2(n7268), .C1(n7604), 
        .C2(n7266), .ZN(n3626) );
  AOI221_X1 U6252 ( .B1(Zzohu6), .B2(n7669), .C1(n7273), .C2(n6578), .A(n2656), 
        .ZN(n3575) );
  INV_X1 U6253 ( .A(n3577), .ZN(n2656) );
  AOI222_X1 U6254 ( .A1(n7645), .A2(V4phu6), .B1(n7696), .B2(Uwdpw6), .C1(
        n7585), .C2(Y2phu6), .ZN(n3577) );
  OAI221_X1 U6255 ( .B1(n7671), .B2(n1858), .C1(n7672), .C2(n872), .A(n1863), 
        .ZN(n7981) );
  NAND2_X1 U6256 ( .A1(L6gpw6[22]), .A2(n866), .ZN(n1863) );
  OAI221_X1 U6257 ( .B1(n7543), .B2(n1858), .C1(n7353), .C2(n872), .A(n1883), 
        .ZN(n8001) );
  NAND2_X1 U6258 ( .A1(L6gpw6[1]), .A2(n866), .ZN(n1883) );
  OAI221_X1 U6259 ( .B1(n7289), .B2(n1858), .C1(n7290), .C2(n872), .A(n1864), 
        .ZN(n7982) );
  NAND2_X1 U6260 ( .A1(L6gpw6[21]), .A2(n866), .ZN(n1864) );
  OAI221_X1 U6261 ( .B1(n7538), .B2(n1858), .C1(n7539), .C2(n872), .A(n1871), 
        .ZN(n7989) );
  NAND2_X1 U6262 ( .A1(L6gpw6[14]), .A2(n866), .ZN(n1871) );
  OAI221_X1 U6263 ( .B1(n7536), .B2(n1858), .C1(n7537), .C2(n872), .A(n1870), 
        .ZN(n7988) );
  NAND2_X1 U6264 ( .A1(L6gpw6[15]), .A2(n866), .ZN(n1870) );
  OAI221_X1 U6265 ( .B1(n7365), .B2(n1858), .C1(n7366), .C2(n872), .A(n1874), 
        .ZN(n7992) );
  NAND2_X1 U6266 ( .A1(L6gpw6[10]), .A2(n866), .ZN(n1874) );
  OAI221_X1 U6267 ( .B1(n7542), .B2(n1858), .C1(n7642), .C2(n872), .A(n1882), 
        .ZN(n8000) );
  NAND2_X1 U6268 ( .A1(L6gpw6[2]), .A2(n1861), .ZN(n1882) );
  OAI221_X1 U6269 ( .B1(n7691), .B2(n1858), .C1(n7692), .C2(n872), .A(n1881), 
        .ZN(n7999) );
  NAND2_X1 U6270 ( .A1(L6gpw6[3]), .A2(n1861), .ZN(n1881) );
  OAI221_X1 U6271 ( .B1(n7686), .B2(n1858), .C1(n7687), .C2(n872), .A(n1880), 
        .ZN(n7998) );
  NAND2_X1 U6272 ( .A1(L6gpw6[4]), .A2(n1861), .ZN(n1880) );
  OAI221_X1 U6273 ( .B1(n7635), .B2(n1858), .C1(n7445), .C2(n872), .A(n1878), 
        .ZN(n7996) );
  NAND2_X1 U6274 ( .A1(L6gpw6[6]), .A2(n1861), .ZN(n1878) );
  OAI221_X1 U6275 ( .B1(n7402), .B2(n1858), .C1(n7403), .C2(n872), .A(n1876), 
        .ZN(n7994) );
  NAND2_X1 U6276 ( .A1(L6gpw6[8]), .A2(n1861), .ZN(n1876) );
  OAI221_X1 U6277 ( .B1(n7361), .B2(n1858), .C1(n7362), .C2(n872), .A(n1869), 
        .ZN(n7987) );
  NAND2_X1 U6278 ( .A1(L6gpw6[16]), .A2(n866), .ZN(n1869) );
  OAI221_X1 U6279 ( .B1(n7367), .B2(n1858), .C1(n7368), .C2(n872), .A(n1868), 
        .ZN(n7986) );
  NAND2_X1 U6280 ( .A1(L6gpw6[17]), .A2(n866), .ZN(n1868) );
  OAI221_X1 U6281 ( .B1(n7390), .B2(n1858), .C1(n7391), .C2(n872), .A(n1867), 
        .ZN(n7985) );
  NAND2_X1 U6282 ( .A1(L6gpw6[18]), .A2(n866), .ZN(n1867) );
  OAI221_X1 U6283 ( .B1(n7379), .B2(n1858), .C1(n7443), .C2(n872), .A(n1866), 
        .ZN(n7984) );
  NAND2_X1 U6284 ( .A1(L6gpw6[19]), .A2(n866), .ZN(n1866) );
  OAI221_X1 U6285 ( .B1(n7275), .B2(n1858), .C1(n7276), .C2(n872), .A(n1860), 
        .ZN(n7979) );
  NAND2_X1 U6286 ( .A1(L6gpw6[12]), .A2(n866), .ZN(n1860) );
  OAI221_X1 U6287 ( .B1(n7338), .B2(n1858), .C1(n7339), .C2(n872), .A(n1879), 
        .ZN(n7997) );
  NAND2_X1 U6288 ( .A1(L6gpw6[5]), .A2(n1861), .ZN(n1879) );
  INV_X1 U6289 ( .A(IRQ[28]), .ZN(n8333) );
  NAND3_X1 U6290 ( .A1(n2850), .A2(n2851), .A3(n1823), .ZN(Pfphu6) );
  INV_X1 U6291 ( .A(n2853), .ZN(n1823) );
  AOI21_X1 U6292 ( .B1(n118), .B2(n1407), .A(n6659), .ZN(n2853) );
  INV_X1 U6293 ( .A(IRQ[23]), .ZN(n8335) );
  INV_X1 U6294 ( .A(IRQ[7]), .ZN(n8348) );
  INV_X1 U6295 ( .A(IRQ[20]), .ZN(n8338) );
  INV_X1 U6296 ( .A(IRQ[22]), .ZN(n8336) );
  INV_X1 U6297 ( .A(IRQ[3]), .ZN(n8352) );
  INV_X1 U6298 ( .A(IRQ[4]), .ZN(n8351) );
  INV_X1 U6299 ( .A(IRQ[6]), .ZN(n8349) );
  INV_X1 U6300 ( .A(IRQ[18]), .ZN(n8340) );
  INV_X1 U6301 ( .A(IRQ[8]), .ZN(n8347) );
  INV_X1 U6302 ( .A(IRQ[16]), .ZN(n8342) );
  INV_X1 U6303 ( .A(IRQ[0]), .ZN(n8355) );
  INV_X1 U6304 ( .A(IRQ[9]), .ZN(n8346) );
  INV_X1 U6305 ( .A(IRQ[19]), .ZN(n8339) );
  INV_X1 U6306 ( .A(IRQ[21]), .ZN(n8337) );
  INV_X1 U6308 ( .A(IRQ[5]), .ZN(n8350) );
  INV_X1 U6309 ( .A(IRQ[17]), .ZN(n8341) );
  INV_X1 U6310 ( .A(IRQ[1]), .ZN(n8354) );
  INV_X1 U6311 ( .A(IRQ[29]), .ZN(n8332) );
  INV_X1 U6312 ( .A(IRQ[2]), .ZN(n8353) );
  INV_X1 U6313 ( .A(IRQ[15]), .ZN(n8343) );
  INV_X1 U6314 ( .A(HRDATA[5]), .ZN(n8324) );
  INV_X1 U6315 ( .A(HRDATA[3]), .ZN(n8326) );
  INV_X1 U6316 ( .A(HRDATA[22]), .ZN(n8308) );
  INV_X1 U6317 ( .A(HRDATA[31]), .ZN(n8299) );
  INV_X1 U6318 ( .A(HRDATA[24]), .ZN(n8306) );
  INV_X1 U6319 ( .A(HRDATA[27]), .ZN(n8303) );
  INV_X1 U6320 ( .A(HRDATA[26]), .ZN(n8304) );
  OAI221_X1 U6321 ( .B1(n7540), .B2(n1858), .C1(n7541), .C2(n872), .A(n1877), 
        .ZN(n7995) );
  NAND2_X1 U6322 ( .A1(L6gpw6[7]), .A2(n1861), .ZN(n1877) );
  OAI221_X1 U6323 ( .B1(n7698), .B2(n1858), .C1(n7699), .C2(n872), .A(n1875), 
        .ZN(n7993) );
  NAND2_X1 U6324 ( .A1(L6gpw6[9]), .A2(n866), .ZN(n1875) );
  OAI221_X1 U6325 ( .B1(n7327), .B2(n1858), .C1(n7444), .C2(n872), .A(n1873), 
        .ZN(n7991) );
  NAND2_X1 U6326 ( .A1(L6gpw6[11]), .A2(n866), .ZN(n1873) );
  OAI221_X1 U6327 ( .B1(n7287), .B2(n1858), .C1(n7288), .C2(n872), .A(n1872), 
        .ZN(n7990) );
  NAND2_X1 U6328 ( .A1(L6gpw6[13]), .A2(n866), .ZN(n1872) );
  OAI221_X1 U6329 ( .B1(n7277), .B2(n1858), .C1(n7278), .C2(n872), .A(n1865), 
        .ZN(n7983) );
  NAND2_X1 U6330 ( .A1(L6gpw6[20]), .A2(n866), .ZN(n1865) );
  OAI221_X1 U6331 ( .B1(n7351), .B2(n1858), .C1(n7352), .C2(n872), .A(n1884), 
        .ZN(n8002) );
  NAND2_X1 U6332 ( .A1(L6gpw6[0]), .A2(n866), .ZN(n1884) );
  INV_X1 U6333 ( .A(HRDATA[30]), .ZN(n8300) );
  INV_X1 U6334 ( .A(HRDATA[21]), .ZN(n8309) );
  INV_X1 U6335 ( .A(HRDATA[17]), .ZN(n8313) );
  INV_X1 U6336 ( .A(HRDATA[14]), .ZN(n8315) );
  INV_X1 U6337 ( .A(HRDATA[13]), .ZN(n8316) );
  INV_X1 U6338 ( .A(HRDATA[12]), .ZN(n8317) );
  INV_X1 U6339 ( .A(HRDATA[10]), .ZN(n8319) );
  INV_X1 U6340 ( .A(HRDATA[8]), .ZN(n8321) );
  OR2_X1 U6341 ( .A1(DBGRESTARTED), .A2(DBGRESTART), .ZN(n4059) );
  INV_X1 U6342 ( .A(n1007), .ZN(n1822) );
  OAI222_X1 U6343 ( .A1(n1008), .A2(n6659), .B1(n1009), .B2(n3115), .C1(n2965), 
        .C2(n8329), .ZN(n1007) );
  INV_X1 U6344 ( .A(n3941), .ZN(n2646) );
  OAI21_X1 U6345 ( .B1(n3942), .B2(n3943), .A(n2831), .ZN(n3941) );
  AOI22_X1 U6346 ( .A1(n7595), .A2(n2830), .B1(n226), .B2(HWDATA[25]), .ZN(
        n3943) );
  AND2_X1 U6347 ( .A1(n6589), .A2(IRQ[25]), .ZN(n3942) );
  OAI221_X1 U6349 ( .B1(n7526), .B2(n1921), .C1(n1922), .C2(n1916), .A(n1917), 
        .ZN(n8006) );
  AOI222_X1 U6350 ( .A1(n1918), .A2(n5042), .B1(n1919), .B2(n470), .C1(n1920), 
        .C2(n4910), .ZN(n1922) );
  AOI21_X1 U6351 ( .B1(n1924), .B2(n5065), .A(n1838), .ZN(n1921) );
  INV_X1 U6352 ( .A(n1914), .ZN(n1838) );
  OAI22_X1 U6353 ( .A1(n7401), .A2(n1859), .B1(n2859), .B2(n2860), .ZN(P9vhu6)
         );
  AOI21_X1 U6354 ( .B1(n2861), .B2(n2862), .A(n2863), .ZN(n2859) );
  INV_X1 U6355 ( .A(n2860), .ZN(n1859) );
  OAI21_X1 U6356 ( .B1(n2871), .B2(n2872), .A(N701), .ZN(n2860) );
  AOI221_X1 U6357 ( .B1(Npghu6), .B2(n7550), .C1(Nwdpw6), .C2(n7597), .A(n2647), .ZN(n3678) );
  INV_X1 U6358 ( .A(n3745), .ZN(n2647) );
  AOI22_X1 U6359 ( .A1(n7583), .A2(R2phu6), .B1(n7601), .B2(Qyohu6), .ZN(n3745) );
  INV_X1 U6360 ( .A(n1362), .ZN(n2100) );
  AOI221_X1 U6361 ( .B1(n7481), .B2(n1363), .C1(n1364), .C2(n1365), .A(n1366), 
        .ZN(n1362) );
  NOR2_X1 U6362 ( .A1(n4112), .A2(n4123), .ZN(n1363) );
  INV_X1 U6363 ( .A(n3655), .ZN(n2682) );
  AOI22_X1 U6364 ( .A1(n7591), .A2(n7262), .B1(n7689), .B2(n7263), .ZN(n3655)
         );
  NOR2_X1 U6365 ( .A1(n3859), .A2(n2937), .ZN(A4phu6) );
  INV_X1 U6366 ( .A(n5542), .ZN(n2937) );
  OAI211_X1 U6367 ( .C1(n8350), .C2(n8289), .A(n5543), .B(n3861), .ZN(n5542)
         );
  OAI21_X1 U6368 ( .B1(n4072), .B2(n672), .A(n6576), .ZN(n5543) );
  AOI221_X1 U6369 ( .B1(n7272), .B2(n6582), .C1(n7271), .C2(n7357), .A(n2674), 
        .ZN(n3574) );
  INV_X1 U6370 ( .A(n3603), .ZN(n2674) );
  AOI22_X1 U6371 ( .A1(n7594), .A2(n7269), .B1(n7596), .B2(n7270), .ZN(n3603)
         );
  NAND2_X1 U6372 ( .A1(n1961), .A2(n1962), .ZN(n8009) );
  OAI21_X1 U6373 ( .B1(n6887), .B2(n1963), .A(n8162), .ZN(n1962) );
  INV_X1 U6374 ( .A(n4120), .ZN(n2486) );
  OAI211_X1 U6375 ( .C1(n4121), .C2(n234), .A(n4122), .B(IRQ[27]), .ZN(n4120)
         );
  AOI211_X1 U6376 ( .C1(n3849), .C2(n6573), .A(n233), .B(n4023), .ZN(n4122) );
  INV_X1 U6377 ( .A(n4021), .ZN(n3849) );
  INV_X1 U6378 ( .A(n3777), .ZN(n2485) );
  OAI211_X1 U6379 ( .C1(n3778), .C2(n234), .A(n3779), .B(IRQ[24]), .ZN(n3777)
         );
  AOI211_X1 U6380 ( .C1(n3845), .C2(n6580), .A(n233), .B(n3758), .ZN(n3779) );
  INV_X1 U6381 ( .A(n3756), .ZN(n3845) );
  INV_X1 U6382 ( .A(n2300), .ZN(n2479) );
  OAI211_X1 U6383 ( .C1(n234), .C2(n2302), .A(n2303), .B(NMI), .ZN(n2300) );
  AOI21_X1 U6384 ( .B1(n3843), .B2(n7549), .A(n2305), .ZN(n2303) );
  NOR2_X1 U6385 ( .A1(n233), .A2(n3952), .ZN(n2302) );
  INV_X1 U6386 ( .A(STCALIB[5]), .ZN(n8360) );
  OAI222_X1 U6387 ( .A1(n8357), .A2(n4788), .B1(n2202), .B2(n7535), .C1(n1893), 
        .C2(n7369), .ZN(n5927) );
  INV_X1 U6388 ( .A(STCALIB[23]), .ZN(n8357) );
  NOR3_X1 U6389 ( .A1(n7414), .A2(n6836), .A3(n7456), .ZN(n2307) );
  NOR3_X1 U6390 ( .A1(n6836), .A2(n6643), .A3(n7414), .ZN(n2333) );
  NAND4_X1 U6391 ( .A1(n1311), .A2(n1344), .A3(n1345), .A4(n7411), .ZN(n1020)
         );
  NOR3_X1 U6392 ( .A1(n555), .A2(n7313), .A3(n548), .ZN(n663) );
  NOR2_X1 U6393 ( .A1(n4395), .A2(n7363), .ZN(n5406) );
  NOR4_X1 U6394 ( .A1(n7648), .A2(n7450), .A3(n4149), .A4(n969), .ZN(n938) );
  OR3_X1 U6395 ( .A1(n7428), .A2(n7387), .A3(n7427), .ZN(n969) );
  NAND4_X1 U6396 ( .A1(n5406), .A2(n7371), .A3(n4410), .A4(n4160), .ZN(n1893)
         );
  NOR3_X1 U6397 ( .A1(n2015), .A2(n7317), .A3(n4036), .ZN(n544) );
  NOR2_X1 U6398 ( .A1(n4406), .A2(n7438), .ZN(n1183) );
  NOR3_X1 U6399 ( .A1(n3623), .A2(n7399), .A3(n2243), .ZN(n1698) );
  OAI211_X1 U6400 ( .C1(n3107), .C2(n5570), .A(n6081), .B(n5577), .ZN(n4267)
         );
  NAND3_X1 U6401 ( .A1(n7703), .A2(n8175), .A3(n6040), .ZN(n6081) );
  OR2_X1 U6402 ( .A1(n948), .A2(n152), .ZN(n954) );
  NAND3_X1 U6403 ( .A1(n8164), .A2(n8172), .A3(n3894), .ZN(n953) );
  AOI21_X1 U6404 ( .B1(n1731), .B2(n3684), .A(n7399), .ZN(n5036) );
  AOI211_X1 U6405 ( .C1(n3828), .C2(n3800), .A(n2447), .B(n7332), .ZN(n5390)
         );
  OAI21_X1 U6406 ( .B1(n7505), .B2(n7393), .A(n7519), .ZN(n4220) );
  OAI21_X1 U6407 ( .B1(n2933), .B2(n7510), .A(n475), .ZN(n4221) );
  NOR3_X1 U6408 ( .A1(n7548), .A2(n7371), .A3(n4160), .ZN(n5483) );
  NOR2_X1 U6409 ( .A1(n5980), .A2(n7371), .ZN(n5345) );
  AOI21_X1 U6411 ( .B1(n429), .B2(n1943), .A(n1944), .ZN(n1942) );
  OAI21_X1 U6412 ( .B1(n254), .B2(n2524), .A(n1949), .ZN(n1943) );
  NAND3_X1 U6413 ( .A1(n1938), .A2(n1950), .A3(n7497), .ZN(n1949) );
  NOR2_X1 U6414 ( .A1(n4028), .A2(n7310), .ZN(n610) );
  NAND4_X1 U6415 ( .A1(n7387), .A2(n7427), .A3(n7428), .A4(n7648), .ZN(n152)
         );
  NOR4_X1 U6416 ( .A1(n3682), .A2(n2377), .A3(n1958), .A4(n7518), .ZN(n41) );
  NOR2_X1 U6417 ( .A1(n7534), .A2(n7363), .ZN(n5545) );
  NAND3_X1 U6418 ( .A1(n1344), .A2(n7411), .A3(n1969), .ZN(n1000) );
  NOR3_X1 U6419 ( .A1(n5070), .A2(n7529), .A3(n4261), .ZN(n4834) );
  NOR2_X1 U6420 ( .A1(n470), .A2(n7516), .ZN(n1595) );
  NOR3_X1 U6421 ( .A1(n7476), .A2(n228), .A3(n4194), .ZN(n2876) );
  NOR2_X1 U6422 ( .A1(n7510), .A2(n524), .ZN(n1744) );
  NOR2_X1 U6423 ( .A1(n2124), .A2(n7399), .ZN(n2921) );
  AOI211_X1 U6424 ( .C1(n6672), .C2(n6671), .A(n3135), .B(n641), .ZN(n620) );
  INV_X1 U6425 ( .A(n642), .ZN(n3135) );
  NAND2_X1 U6426 ( .A1(n7312), .A2(n7315), .ZN(n548) );
  NAND2_X1 U6427 ( .A1(n7460), .A2(n2307), .ZN(Frmhu6) );
  NAND2_X1 U6428 ( .A1(n7464), .A2(n2333), .ZN(G9khu6) );
  OAI222_X1 U6429 ( .A1(n6632), .A2(n4729), .B1(n6581), .B2(n4730), .C1(n7364), 
        .C2(n2825), .ZN(n1032) );
  NAND3_X1 U6430 ( .A1(n642), .A2(n4033), .A3(n7320), .ZN(n2159) );
  AOI222_X1 U6431 ( .A1(n2489), .A2(n2232), .B1(n7529), .B2(n2495), .C1(n2842), 
        .C2(n4993), .ZN(n2841) );
  NAND4_X1 U6432 ( .A1(n2129), .A2(HALTED), .A3(n7371), .A4(n4160), .ZN(n1419)
         );
  NOR3_X1 U6433 ( .A1(n7548), .A2(n7383), .A3(n3288), .ZN(n2129) );
  NOR2_X1 U6434 ( .A1(n3225), .A2(n7308), .ZN(n648) );
  AOI222_X1 U6435 ( .A1(n473), .A2(n1612), .B1(n1684), .B2(n7516), .C1(n1685), 
        .C2(n2262), .ZN(n1676) );
  NOR3_X1 U6436 ( .A1(n4688), .A2(n7492), .A3(n522), .ZN(n1533) );
  AOI221_X1 U6437 ( .B1(n7282), .B2(n1477), .C1(n1478), .C2(n7492), .A(n1479), 
        .ZN(n1471) );
  NAND2_X1 U6438 ( .A1(n1480), .A2(n3830), .ZN(n1479) );
  NAND2_X1 U6439 ( .A1(n5225), .A2(n1483), .ZN(n1477) );
  NAND3_X1 U6440 ( .A1(n1482), .A2(n516), .A3(n267), .ZN(n1480) );
  NAND2_X1 U6441 ( .A1(n5973), .A2(n7398), .ZN(n903) );
  OAI221_X1 U6442 ( .B1(n633), .B2(n548), .C1(n7312), .C2(n3202), .A(n634), 
        .ZN(n7839) );
  OAI21_X1 U6443 ( .B1(n4022), .B2(n3203), .A(n636), .ZN(n634) );
  NOR4_X1 U6444 ( .A1(n637), .A2(n638), .A3(n639), .A4(n620), .ZN(n633) );
  OAI21_X1 U6445 ( .B1(n7314), .B2(n645), .A(n3191), .ZN(n637) );
  NOR3_X1 U6446 ( .A1(n4160), .A2(n7548), .A3(n4182), .ZN(n5971) );
  OAI21_X1 U6447 ( .B1(n7318), .B2(n382), .A(n551), .ZN(n2183) );
  NAND4_X1 U6448 ( .A1(n1857), .A2(n7371), .A3(n4410), .A4(n4160), .ZN(n2151)
         );
  OAI221_X1 U6449 ( .B1(n7595), .B2(n4730), .C1(n7581), .C2(n4729), .A(n903), 
        .ZN(n1164) );
  NAND4_X1 U6450 ( .A1(n1538), .A2(n7433), .A3(n7399), .A4(n7510), .ZN(n3966)
         );
  NOR4_X1 U6451 ( .A1(n7424), .A2(n152), .A3(n947), .A4(n948), .ZN(n932) );
  OAI211_X1 U6452 ( .C1(n7510), .C2(n2371), .A(n2372), .B(n2373), .ZN(n1920)
         );
  OAI211_X1 U6453 ( .C1(n1744), .C2(n2375), .A(n230), .B(n2376), .ZN(n2372) );
  AOI21_X1 U6454 ( .B1(n518), .B2(n1457), .A(n2374), .ZN(n2373) );
  NOR3_X1 U6455 ( .A1(n7447), .A2(n7437), .A3(n7641), .ZN(n957) );
  NOR2_X1 U6456 ( .A1(n7310), .A2(n7309), .ZN(n619) );
  OAI222_X1 U6457 ( .A1(n2574), .A2(n2694), .B1(n7381), .B2(n2576), .C1(n7399), 
        .C2(n2699), .ZN(n2573) );
  NOR4_X1 U6458 ( .A1(n2587), .A2(n1683), .A3(n7433), .A4(n7523), .ZN(n2574)
         );
  AOI221_X1 U6459 ( .B1(n2577), .B2(n529), .C1(n1685), .C2(n2578), .A(n2579), 
        .ZN(n2576) );
  OAI211_X1 U6460 ( .C1(n2588), .C2(n2589), .A(n7381), .B(n7519), .ZN(n2587)
         );
  OAI221_X1 U6461 ( .B1(n7283), .B2(n4193), .C1(n508), .C2(n4628), .A(n6562), 
        .ZN(n6557) );
  AOI221_X1 U6462 ( .B1(n1463), .B2(n508), .C1(n5574), .C2(n272), .A(n2743), 
        .ZN(n6562) );
  OAI221_X1 U6463 ( .B1(n93), .B2(n2256), .C1(n2699), .C2(n4186), .A(n1583), 
        .ZN(n1579) );
  AOI222_X1 U6464 ( .A1(n1584), .A2(n1585), .B1(n1586), .B2(n1587), .C1(n1588), 
        .C2(n270), .ZN(n1583) );
  OAI221_X1 U6465 ( .B1(n7514), .B2(n1589), .C1(n7519), .C2(n5042), .A(n1591), 
        .ZN(n1585) );
  AOI221_X1 U6466 ( .B1(n1592), .B2(n7514), .C1(n1593), .C2(n464), .A(n1594), 
        .ZN(n1591) );
  OAI221_X1 U6467 ( .B1(n3113), .B2(n3715), .C1(n3716), .C2(n5225), .A(n3717), 
        .ZN(n699) );
  OAI211_X1 U6468 ( .C1(n810), .C2(n2113), .A(n7533), .B(n3718), .ZN(n3717) );
  NOR3_X1 U6469 ( .A1(n3719), .A2(n3720), .A3(n3721), .ZN(n3716) );
  NOR2_X1 U6470 ( .A1(n477), .A2(n7492), .ZN(n3718) );
  NOR2_X1 U6471 ( .A1(n2825), .A2(n7383), .ZN(n3687) );
  OAI22_X1 U6472 ( .A1(n7325), .A2(n7359), .B1(n7329), .B2(n3241), .ZN(n2999)
         );
  AOI221_X1 U6473 ( .B1(n1519), .B2(n1520), .C1(n7378), .C2(n1521), .A(n1522), 
        .ZN(n1499) );
  OAI22_X1 U6474 ( .A1(n4693), .A2(n4265), .B1(n3623), .B2(n1528), .ZN(n1521)
         );
  NOR3_X1 U6475 ( .A1(n4668), .A2(n1524), .A3(n4189), .ZN(n1522) );
  AOI221_X1 U6476 ( .B1(n4670), .B2(n4572), .C1(n7505), .C2(n5042), .A(n3530), 
        .ZN(n3529) );
  OAI21_X1 U6477 ( .B1(n4669), .B2(n5042), .A(n4555), .ZN(n3530) );
  AOI221_X1 U6478 ( .B1(n2806), .B2(n1706), .C1(n7524), .C2(n5065), .A(n3164), 
        .ZN(n3163) );
  OAI22_X1 U6479 ( .A1(n2807), .A2(n3566), .B1(n57), .B2(n3099), .ZN(n3164) );
  AOI221_X1 U6480 ( .B1(n1964), .B2(n4993), .C1(n1511), .C2(n1512), .A(n1513), 
        .ZN(n1501) );
  INV_X1 U6481 ( .A(n1518), .ZN(n1964) );
  AOI221_X1 U6482 ( .B1(n2893), .B2(n5047), .C1(n1907), .C2(n3526), .A(n3527), 
        .ZN(n3523) );
  OAI211_X1 U6483 ( .C1(n270), .C2(n4993), .A(n4669), .B(n7518), .ZN(n3526) );
  AOI22_X1 U6484 ( .A1(n7492), .A2(n2748), .B1(n2749), .B2(n230), .ZN(n2747)
         );
  NAND4_X1 U6485 ( .A1(n2750), .A2(n2751), .A3(n511), .A4(n2752), .ZN(n2749)
         );
  OAI21_X1 U6486 ( .B1(n1478), .B2(n7282), .A(n1615), .ZN(n2751) );
  OAI222_X1 U6487 ( .A1(n4237), .A2(n2547), .B1(n1622), .B2(n3549), .C1(n7283), 
        .C2(n1623), .ZN(n1548) );
  AOI21_X1 U6488 ( .B1(n1628), .B2(n265), .A(n1629), .ZN(n1622) );
  AOI221_X1 U6489 ( .B1(n2124), .B2(n1624), .C1(n1625), .C2(n1626), .A(n1627), 
        .ZN(n1623) );
  NOR3_X1 U6490 ( .A1(n2594), .A2(n522), .A3(n3628), .ZN(n1629) );
  NAND4_X1 U6491 ( .A1(n5022), .A2(n4685), .A3(n5023), .A4(n5024), .ZN(n3027)
         );
  OAI21_X1 U6492 ( .B1(n7516), .B2(n7433), .A(n2893), .ZN(n5022) );
  OAI21_X1 U6493 ( .B1(n521), .B2(n4932), .A(n479), .ZN(n5023) );
  AOI21_X1 U6494 ( .B1(n3077), .B2(n2262), .A(n3075), .ZN(n5024) );
  OAI222_X1 U6495 ( .A1(n6759), .A2(n2194), .B1(n6774), .B2(n2197), .C1(n7623), 
        .C2(n2196), .ZN(n5479) );
  NAND4_X1 U6497 ( .A1(n6082), .A2(n5600), .A3(n5575), .A4(n5569), .ZN(n4526)
         );
  NAND3_X1 U6498 ( .A1(n7626), .A2(n4694), .A3(n6040), .ZN(n6082) );
  NAND4_X1 U6499 ( .A1(n7316), .A2(n7319), .A3(n641), .A4(n600), .ZN(n2165) );
  AOI211_X1 U6500 ( .C1(n2494), .C2(n2495), .A(n2496), .B(n2497), .ZN(n2493)
         );
  XNOR2_X1 U6501 ( .A(n2499), .B(n5299), .ZN(n2494) );
  NOR3_X1 U6502 ( .A1(n4187), .A2(n7516), .A3(n2498), .ZN(n2497) );
  OR2_X1 U6503 ( .A1(n2501), .A2(n7530), .ZN(n2499) );
  NAND4_X1 U6504 ( .A1(n1488), .A2(n7492), .A3(n1457), .A4(n1489), .ZN(n1487)
         );
  OAI22_X1 U6505 ( .A1(n7518), .A2(n5037), .B1(n7516), .B2(n4566), .ZN(n1489)
         );
  AOI211_X1 U6506 ( .C1(n7519), .C2(n270), .A(n1595), .B(n1760), .ZN(n1759) );
  INV_X1 U6507 ( .A(n2007), .ZN(n3129) );
  AOI211_X1 U6508 ( .C1(n236), .C2(n6648), .A(n542), .B(n2008), .ZN(n2007) );
  OAI22_X1 U6509 ( .A1(n928), .A2(n7420), .B1(n917), .B2(n7337), .ZN(n2008) );
  INV_X1 U6510 ( .A(n1992), .ZN(n3128) );
  AOI211_X1 U6511 ( .C1(n236), .C2(n6654), .A(n542), .B(n1993), .ZN(n1992) );
  OAI22_X1 U6512 ( .A1(n928), .A2(n6625), .B1(n913), .B2(n6624), .ZN(n1993) );
  NOR2_X1 U6513 ( .A1(n3246), .A2(n7393), .ZN(n2996) );
  NAND3_X1 U6514 ( .A1(n7316), .A2(n7319), .A3(n663), .ZN(n2015) );
  OAI21_X1 U6515 ( .B1(n2700), .B2(n5111), .A(n4629), .ZN(n3425) );
  OR4_X1 U6516 ( .A1(n4651), .A2(n7628), .A3(n7375), .A4(n7279), .ZN(n4629) );
  NOR4_X1 U6517 ( .A1(n1647), .A2(n1648), .A3(n1649), .A4(n1475), .ZN(n1646)
         );
  OAI221_X1 U6518 ( .B1(n1651), .B2(n522), .C1(n4749), .C2(n3787), .A(n3744), 
        .ZN(n1647) );
  INV_X1 U6519 ( .A(n1653), .ZN(n3744) );
  OAI221_X1 U6520 ( .B1(n7519), .B2(n2235), .C1(n7329), .C2(n2254), .A(n3003), 
        .ZN(n2981) );
  AOI22_X1 U6521 ( .A1(n2247), .A2(n4908), .B1(n2489), .B2(n3065), .ZN(n3003)
         );
  NOR2_X1 U6522 ( .A1(n3200), .A2(n7311), .ZN(n2054) );
  NOR2_X1 U6523 ( .A1(n7480), .A2(n7481), .ZN(n2149) );
  OAI222_X1 U6524 ( .A1(n7416), .A2(n537), .B1(n908), .B2(n4048), .C1(n7420), 
        .C2(n917), .ZN(n8037) );
  OAI222_X1 U6525 ( .A1(n6672), .A2(n537), .B1(n7405), .B2(n908), .C1(n6671), 
        .C2(n917), .ZN(n7304) );
  OAI222_X1 U6526 ( .A1(n6612), .A2(n537), .B1(n6656), .B2(n908), .C1(n6611), 
        .C2(n917), .ZN(n7296) );
  OAI222_X1 U6527 ( .A1(n6609), .A2(n537), .B1(n6662), .B2(n908), .C1(n6623), 
        .C2(n917), .ZN(n7295) );
  OAI222_X1 U6528 ( .A1(n6620), .A2(n537), .B1(n6652), .B2(n908), .C1(n6619), 
        .C2(n917), .ZN(n7302) );
  OAI222_X1 U6529 ( .A1(n6616), .A2(n537), .B1(n6666), .B2(n908), .C1(n6615), 
        .C2(n917), .ZN(n7299) );
  OAI222_X1 U6530 ( .A1(n6671), .A2(n537), .B1(n6651), .B2(n908), .C1(n6621), 
        .C2(n917), .ZN(n7303) );
  OAI222_X1 U6531 ( .A1(n6617), .A2(n537), .B1(n6667), .B2(n908), .C1(n6616), 
        .C2(n917), .ZN(n7300) );
  OAI222_X1 U6532 ( .A1(n6613), .A2(n537), .B1(n7389), .B2(n908), .C1(n6612), 
        .C2(n917), .ZN(n7297) );
  OAI222_X1 U6533 ( .A1(n6614), .A2(n537), .B1(n6664), .B2(n908), .C1(n6613), 
        .C2(n917), .ZN(n7298) );
  OAI222_X1 U6534 ( .A1(n6618), .A2(n537), .B1(n6665), .B2(n908), .C1(n6617), 
        .C2(n917), .ZN(n7301) );
  OAI22_X1 U6535 ( .A1(n7537), .A2(n1893), .B1(n7536), .B2(n2202), .ZN(n5979)
         );
  NAND2_X1 U6536 ( .A1(n7459), .A2(n2307), .ZN(Ypmhu6) );
  NAND2_X1 U6537 ( .A1(n7463), .A2(n2333), .ZN(Y7khu6) );
  OAI22_X1 U6538 ( .A1(n7518), .A2(n2244), .B1(n2272), .B2(n2990), .ZN(n2982)
         );
  XNOR2_X1 U6539 ( .A(n3697), .B(n2503), .ZN(n2990) );
  OAI221_X1 U6540 ( .B1(n7505), .B2(n2235), .C1(n7325), .C2(n2254), .A(n3248), 
        .ZN(n3229) );
  AOI22_X1 U6541 ( .A1(n2247), .A2(n3690), .B1(n2489), .B2(n4841), .ZN(n3248)
         );
  OAI22_X1 U6542 ( .A1(n7399), .A2(n2697), .B1(n475), .B2(n2256), .ZN(n1753)
         );
  OAI221_X1 U6543 ( .B1(n3180), .B2(n6622), .C1(n2015), .C2(n7320), .A(n3190), 
        .ZN(n2014) );
  OAI22_X1 U6544 ( .A1(n7374), .A2(n4738), .B1(n7518), .B2(n4241), .ZN(n4238)
         );
  OAI22_X1 U6545 ( .A1(n7543), .A2(n2202), .B1(n3968), .B2(n2825), .ZN(n4771)
         );
  OAI22_X1 U6546 ( .A1(n7691), .A2(n2202), .B1(n5088), .B2(n2825), .ZN(n5670)
         );
  OAI22_X1 U6547 ( .A1(n7542), .A2(n2202), .B1(n5111), .B2(n2825), .ZN(n4712)
         );
  OAI22_X1 U6548 ( .A1(n7538), .A2(n2202), .B1(n6627), .B2(n4729), .ZN(n5469)
         );
  NOR2_X1 U6549 ( .A1(n4054), .A2(n7451), .ZN(n1311) );
  OAI21_X1 U6550 ( .B1(n2650), .B2(n2818), .A(n1794), .ZN(n7957) );
  OAI221_X1 U6551 ( .B1(n352), .B2(n2818), .C1(n1796), .C2(n3851), .A(n6681), 
        .ZN(n1794) );
  OAI221_X1 U6552 ( .B1(n1022), .B2(n1000), .C1(n6852), .C2(n990), .A(n1023), 
        .ZN(n1015) );
  NOR2_X1 U6553 ( .A1(n3786), .A2(n2519), .ZN(n1022) );
  NOR2_X1 U6554 ( .A1(n918), .A2(n7424), .ZN(n920) );
  NAND4_X1 U6555 ( .A1(n7378), .A2(n1538), .A3(n7355), .A4(n7354), .ZN(n1534)
         );
  AOI21_X1 U6556 ( .B1(n3244), .B2(n7505), .A(n3240), .ZN(n3243) );
  NAND4_X1 U6557 ( .A1(n4317), .A2(n7518), .A3(n475), .A4(n1840), .ZN(n4316)
         );
  NAND3_X1 U6558 ( .A1(n1672), .A2(n7492), .A3(n1754), .ZN(n1750) );
  AOI221_X1 U6559 ( .B1(n1755), .B2(n1756), .C1(n7399), .C2(n1757), .A(n1758), 
        .ZN(n1754) );
  NOR3_X1 U6560 ( .A1(n1739), .A2(n7505), .A3(n3625), .ZN(n1758) );
  OAI222_X1 U6561 ( .A1(n7381), .A2(n5037), .B1(n1759), .B2(n2262), .C1(n7433), 
        .C2(n7510), .ZN(n1757) );
  AOI21_X1 U6562 ( .B1(n3246), .B2(n7393), .A(n2996), .ZN(n3245) );
  NOR2_X1 U6563 ( .A1(n4024), .A2(n7314), .ZN(n655) );
  AOI22_X1 U6564 ( .A1(n7399), .A2(n2375), .B1(n1584), .B2(n7518), .ZN(n5038)
         );
  NAND4_X1 U6565 ( .A1(n2784), .A2(n2785), .A3(n3127), .A4(n4035), .ZN(n532)
         );
  NAND2_X1 U6566 ( .A1(n7318), .A2(n2057), .ZN(n2785) );
  NOR3_X1 U6567 ( .A1(n2697), .A2(n7433), .A3(n270), .ZN(n2764) );
  NAND4_X1 U6568 ( .A1(n1970), .A2(n1900), .A3(n3260), .A4(n3261), .ZN(n3217)
         );
  AOI22_X1 U6569 ( .A1(n2875), .A2(n7259), .B1(n496), .B2(n7282), .ZN(n3260)
         );
  INV_X1 U6570 ( .A(n3270), .ZN(n1900) );
  AOI221_X1 U6572 ( .B1(n1488), .B2(n3262), .C1(n1672), .C2(n3263), .A(n3264), 
        .ZN(n3261) );
  XNOR2_X1 U6573 ( .A(n7359), .B(n7325), .ZN(n3241) );
  OAI22_X1 U6574 ( .A1(n7384), .A2(n4729), .B1(n6575), .B2(n4730), .ZN(n5398)
         );
  NAND2_X1 U6575 ( .A1(n4751), .A2(n2165), .ZN(n556) );
  NAND4_X1 U6576 ( .A1(n6673), .A2(n7336), .A3(n7417), .A4(n534), .ZN(n4751)
         );
  XNOR2_X1 U6577 ( .A(n3894), .B(n7423), .ZN(n923) );
  XNOR2_X1 U6578 ( .A(n8253), .B(n7437), .ZN(n944) );
  OAI221_X1 U6579 ( .B1(n1554), .B2(n4693), .C1(n1555), .C2(n3623), .A(n1556), 
        .ZN(n1549) );
  AOI221_X1 U6580 ( .B1(n1567), .B2(n1620), .C1(n1621), .C2(n513), .A(n1462), 
        .ZN(n1554) );
  AOI221_X1 U6581 ( .B1(n1615), .B2(n4932), .C1(n3549), .C2(n529), .A(n1617), 
        .ZN(n1555) );
  AOI22_X1 U6583 ( .A1(n1557), .A2(n230), .B1(n7510), .B2(n90), .ZN(n1556) );
  OAI22_X1 U6584 ( .A1(n1835), .A2(n800), .B1(n7536), .B2(n799), .ZN(n7716) );
  OAI22_X1 U6587 ( .A1(n1835), .A2(n2897), .B1(n7567), .B2(n2105), .ZN(n7717)
         );
  OAI22_X1 U6588 ( .A1(n1835), .A2(n2989), .B1(n7618), .B2(n2101), .ZN(n7715)
         );
  OAI22_X1 U6589 ( .A1(n1835), .A2(n2983), .B1(n7606), .B2(n2099), .ZN(n7714)
         );
  OAI22_X1 U6591 ( .A1(n1835), .A2(n2992), .B1(n7562), .B2(n2095), .ZN(n7713)
         );
  OAI22_X1 U6592 ( .A1(n1835), .A2(n2885), .B1(n7622), .B2(n2093), .ZN(n7712)
         );
  OAI22_X1 U6593 ( .A1(n1835), .A2(n2906), .B1(n7611), .B2(n2091), .ZN(n7711)
         );
  OAI22_X1 U6594 ( .A1(n1835), .A2(n2987), .B1(n7553), .B2(n2097), .ZN(n7710)
         );
  OAI22_X1 U6595 ( .A1(n1835), .A2(n2883), .B1(n7556), .B2(n2089), .ZN(n7709)
         );
  XNOR2_X1 U6596 ( .A(n6604), .B(n6675), .ZN(n2168) );
  NAND2_X1 U6597 ( .A1(n7505), .A2(n464), .ZN(n1948) );
  OAI21_X1 U6598 ( .B1(n3113), .B2(n492), .A(n7492), .ZN(n1483) );
  OAI211_X1 U6599 ( .C1(n922), .C2(n3886), .A(n957), .B(n7450), .ZN(n947) );
  OAI22_X1 U6600 ( .A1(n7414), .A2(n3007), .B1(n1832), .B2(n2446), .ZN(W0xhu6)
         );
  OAI21_X1 U6601 ( .B1(n7519), .B2(n2244), .A(n3235), .ZN(n3230) );
  OAI211_X1 U6602 ( .C1(n3236), .C2(n3237), .A(n2846), .B(n3001), .ZN(n3235)
         );
  OAI21_X1 U6603 ( .B1(n6430), .B2(n3804), .A(n6431), .ZN(n4557) );
  NOR3_X1 U6604 ( .A1(n4563), .A2(n5550), .A3(n4562), .ZN(n6430) );
  NAND4_X1 U6606 ( .A1(n7326), .A2(n7529), .A3(n7286), .A4(n6432), .ZN(n6431)
         );
  NOR4_X1 U6607 ( .A1(n5070), .A2(n516), .A3(n3860), .A4(n3083), .ZN(n6432) );
  OAI22_X1 U6608 ( .A1(n2671), .A2(n800), .B1(n7671), .B2(n799), .ZN(n6984) );
  OAI22_X1 U6609 ( .A1(n2676), .A2(n800), .B1(n7535), .B2(n799), .ZN(n7199) );
  OAI22_X1 U6610 ( .A1(n2671), .A2(n2883), .B1(n7678), .B2(n2089), .ZN(n6977)
         );
  OAI22_X1 U6611 ( .A1(n2671), .A2(n2906), .B1(n7677), .B2(n2091), .ZN(n6978)
         );
  OAI22_X1 U6612 ( .A1(n2671), .A2(n2885), .B1(n6735), .B2(n2093), .ZN(n6979)
         );
  OAI22_X1 U6613 ( .A1(n2671), .A2(n2992), .B1(n7676), .B2(n2095), .ZN(n6980)
         );
  OAI22_X1 U6614 ( .A1(n2671), .A2(n2987), .B1(n7675), .B2(n2097), .ZN(n6981)
         );
  OAI22_X1 U6615 ( .A1(n2671), .A2(n2983), .B1(n7674), .B2(n2099), .ZN(n6982)
         );
  OAI22_X1 U6616 ( .A1(n2671), .A2(n2989), .B1(n7673), .B2(n2101), .ZN(n6983)
         );
  OAI22_X1 U6617 ( .A1(n2671), .A2(n2897), .B1(n7670), .B2(n2105), .ZN(n6985)
         );
  OAI22_X1 U6618 ( .A1(n2676), .A2(n2883), .B1(n7557), .B2(n2089), .ZN(n7010)
         );
  OAI22_X1 U6619 ( .A1(n2676), .A2(n2987), .B1(n7554), .B2(n2097), .ZN(n7014)
         );
  OAI22_X1 U6620 ( .A1(n2676), .A2(n2897), .B1(n7566), .B2(n2105), .ZN(n7034)
         );
  OAI22_X1 U6621 ( .A1(n2676), .A2(n2992), .B1(n7563), .B2(n2095), .ZN(n7040)
         );
  OAI22_X1 U6622 ( .A1(n2676), .A2(n2989), .B1(n7619), .B2(n2101), .ZN(n7046)
         );
  OAI22_X1 U6623 ( .A1(n2676), .A2(n2885), .B1(n6777), .B2(n2093), .ZN(n7047)
         );
  OAI22_X1 U6624 ( .A1(n2676), .A2(n2983), .B1(n7607), .B2(n2099), .ZN(n7056)
         );
  OAI22_X1 U6625 ( .A1(n2676), .A2(n2906), .B1(n7612), .B2(n2091), .ZN(n7060)
         );
  OAI22_X1 U6626 ( .A1(n7606), .A2(n2198), .B1(n7556), .B2(n2193), .ZN(n5977)
         );
  OAI22_X1 U6627 ( .A1(n7566), .A2(n2200), .B1(n7619), .B2(n2199), .ZN(n5925)
         );
  OAI22_X1 U6628 ( .A1(n7567), .A2(n2200), .B1(n7618), .B2(n2199), .ZN(n5975)
         );
  OAI22_X1 U6629 ( .A1(n356), .A2(n2883), .B1(n7558), .B2(n2089), .ZN(n7008)
         );
  OAI22_X1 U6630 ( .A1(n356), .A2(n2987), .B1(n7555), .B2(n2097), .ZN(n7012)
         );
  OAI22_X1 U6631 ( .A1(n356), .A2(n2897), .B1(n7565), .B2(n2105), .ZN(n7036)
         );
  OAI22_X1 U6632 ( .A1(n356), .A2(n2992), .B1(n7564), .B2(n2095), .ZN(n7038)
         );
  OAI22_X1 U6633 ( .A1(n356), .A2(n2989), .B1(n7620), .B2(n2101), .ZN(n7044)
         );
  OAI22_X1 U6634 ( .A1(n356), .A2(n2885), .B1(n7624), .B2(n2093), .ZN(n7049)
         );
  OAI22_X1 U6635 ( .A1(n356), .A2(n2983), .B1(n7609), .B2(n2099), .ZN(n7054)
         );
  OAI22_X1 U6636 ( .A1(n356), .A2(n2906), .B1(n7614), .B2(n2091), .ZN(n7058)
         );
  AOI21_X1 U6637 ( .B1(n2297), .B2(n4047), .A(n7455), .ZN(Edkhu6) );
  AOI21_X1 U6638 ( .B1(n733), .B2(n4047), .A(n7454), .ZN(Avmhu6) );
  NOR2_X1 U6639 ( .A1(n4324), .A2(n7425), .ZN(n1287) );
  NAND2_X1 U6640 ( .A1(n3066), .A2(n4584), .ZN(n101) );
  NAND3_X1 U6641 ( .A1(n7400), .A2(n4458), .A3(n7530), .ZN(n4584) );
  OAI22_X1 U6642 ( .A1(n6772), .A2(n2200), .B1(n6776), .B2(n2199), .ZN(n5486)
         );
  OAI22_X1 U6643 ( .A1(n7617), .A2(n2199), .B1(n6702), .B2(n2196), .ZN(n5466)
         );
  OAI22_X1 U6644 ( .A1(n7674), .A2(n2198), .B1(n7678), .B2(n2193), .ZN(n5525)
         );
  OAI22_X1 U6645 ( .A1(n7670), .A2(n2200), .B1(n7673), .B2(n2199), .ZN(n5524)
         );
  NAND2_X1 U6646 ( .A1(n7318), .A2(n4033), .ZN(n600) );
  OAI22_X1 U6647 ( .A1(n7607), .A2(n2198), .B1(n7557), .B2(n2193), .ZN(n5926)
         );
  OAI22_X1 U6648 ( .A1(n6712), .A2(n2197), .B1(n7610), .B2(n2195), .ZN(n5936)
         );
  OAI22_X1 U6649 ( .A1(n7679), .A2(n2106), .B1(n2671), .B2(n2865), .ZN(n6976)
         );
  OAI22_X1 U6650 ( .A1(n7434), .A2(n2106), .B1(n2676), .B2(n2865), .ZN(n7211)
         );
  NAND2_X1 U6651 ( .A1(n7458), .A2(n2307), .ZN(Romhu6) );
  NAND2_X1 U6652 ( .A1(n7462), .A2(n2333), .ZN(Q6khu6) );
  OAI22_X1 U6653 ( .A1(n7318), .A2(n788), .B1(n6569), .B2(n791), .ZN(n7214) );
  OAI22_X1 U6654 ( .A1(n349), .A2(n2883), .B1(n6758), .B2(n2089), .ZN(n7009)
         );
  OAI22_X1 U6655 ( .A1(n349), .A2(n2987), .B1(n6759), .B2(n2097), .ZN(n7013)
         );
  OAI22_X1 U6656 ( .A1(n349), .A2(n2897), .B1(n6772), .B2(n2105), .ZN(n7035)
         );
  OAI22_X1 U6657 ( .A1(n349), .A2(n2992), .B1(n6774), .B2(n2095), .ZN(n7039)
         );
  OAI22_X1 U6658 ( .A1(n349), .A2(n2989), .B1(n6776), .B2(n2101), .ZN(n7045)
         );
  OAI22_X1 U6659 ( .A1(n349), .A2(n2885), .B1(n7623), .B2(n2093), .ZN(n7048)
         );
  OAI22_X1 U6660 ( .A1(n349), .A2(n2983), .B1(n7608), .B2(n2099), .ZN(n7055)
         );
  OAI22_X1 U6661 ( .A1(n349), .A2(n2906), .B1(n7613), .B2(n2091), .ZN(n7059)
         );
  NOR2_X1 U6662 ( .A1(n4410), .A2(n7398), .ZN(n5978) );
  OAI22_X1 U6663 ( .A1(n7613), .A2(n2195), .B1(n7257), .B2(n2151), .ZN(n5480)
         );
  OAI22_X1 U6664 ( .A1(n7331), .A2(n2106), .B1(n356), .B2(n2865), .ZN(n7041)
         );
  OAI22_X1 U6665 ( .A1(n7615), .A2(n2972), .B1(n356), .B2(n2127), .ZN(n7052)
         );
  AOI22_X1 U6666 ( .A1(n1672), .A2(n2265), .B1(n2760), .B2(n449), .ZN(n2744)
         );
  OAI221_X1 U6667 ( .B1(n3547), .B2(n2696), .C1(n7354), .C2(n2614), .A(n2761), 
        .ZN(n2760) );
  INV_X1 U6668 ( .A(n2768), .ZN(n2265) );
  AOI211_X1 U6669 ( .C1(n1576), .C2(n2762), .A(n2763), .B(n2764), .ZN(n2761)
         );
  AOI222_X1 U6670 ( .A1(n7406), .A2(n8164), .B1(n929), .B2(n930), .C1(n7490), 
        .C2(n3895), .ZN(n927) );
  OAI211_X1 U6671 ( .C1(n932), .C2(n933), .A(Jshpw6[6]), .B(n935), .ZN(n930)
         );
  NAND4_X1 U6672 ( .A1(n7407), .A2(n7632), .A3(n7422), .A4(n949), .ZN(n929) );
  NOR3_X1 U6673 ( .A1(n7631), .A2(n7397), .A3(n7422), .ZN(n935) );
  AOI22_X1 U6674 ( .A1(n1532), .A2(n56), .B1(n1533), .B2(n7378), .ZN(n1531) );
  NAND2_X1 U6675 ( .A1(n7317), .A2(n642), .ZN(n535) );
  NAND2_X1 U6676 ( .A1(n2784), .A2(n7318), .ZN(n579) );
  NAND3_X1 U6677 ( .A1(n1612), .A2(n7518), .A3(n7414), .ZN(n1611) );
  AOI21_X1 U6678 ( .B1(n936), .B2(n937), .A(n7407), .ZN(n933) );
  OAI22_X1 U6679 ( .A1(n940), .A2(Jshpw6[5]), .B1(n942), .B2(n938), .ZN(n936)
         );
  NAND3_X1 U6680 ( .A1(n938), .A2(n918), .A3(n939), .ZN(n937) );
  OAI22_X1 U6681 ( .A1(n332), .A2(n800), .B1(n7538), .B2(n799), .ZN(n6938) );
  NAND3_X1 U6682 ( .A1(n649), .A2(n605), .A3(n3138), .ZN(n7840) );
  INV_X1 U6683 ( .A(n651), .ZN(n3138) );
  NAND3_X1 U6684 ( .A1(n663), .A2(n554), .A3(n7321), .ZN(n649) );
  OAI22_X1 U6685 ( .A1(n548), .A2(n652), .B1(n3202), .B2(n653), .ZN(n651) );
  NAND3_X1 U6686 ( .A1(n2377), .A2(n2378), .A3(n2379), .ZN(n1919) );
  AOI22_X1 U6687 ( .A1(n2380), .A2(n230), .B1(n7510), .B2(n90), .ZN(n2379) );
  OAI21_X1 U6688 ( .B1(n3547), .B2(n2243), .A(n2381), .ZN(n2380) );
  OAI221_X1 U6689 ( .B1(n7510), .B2(n1600), .C1(n4670), .C2(n4725), .A(n1601), 
        .ZN(n1577) );
  AOI221_X1 U6690 ( .B1(n1592), .B2(n7514), .C1(n5063), .C2(n464), .A(n1609), 
        .ZN(n1600) );
  AOI22_X1 U6691 ( .A1(n270), .A2(n1602), .B1(n3676), .B2(n2262), .ZN(n1601)
         );
  OAI21_X1 U6692 ( .B1(n270), .B2(n5002), .A(n1611), .ZN(n1609) );
  OAI22_X1 U6693 ( .A1(n332), .A2(n2883), .B1(n6700), .B2(n2089), .ZN(n6931)
         );
  OAI22_X1 U6694 ( .A1(n332), .A2(n2906), .B1(n6701), .B2(n2091), .ZN(n6932)
         );
  OAI22_X1 U6695 ( .A1(n332), .A2(n2885), .B1(n6702), .B2(n2093), .ZN(n6933)
         );
  OAI22_X1 U6696 ( .A1(n332), .A2(n2992), .B1(n7561), .B2(n2095), .ZN(n6934)
         );
  OAI22_X1 U6697 ( .A1(n332), .A2(n2987), .B1(n7552), .B2(n2097), .ZN(n6935)
         );
  OAI22_X1 U6698 ( .A1(n332), .A2(n2983), .B1(n7605), .B2(n2099), .ZN(n6936)
         );
  OAI22_X1 U6699 ( .A1(n332), .A2(n2989), .B1(n7617), .B2(n2101), .ZN(n6937)
         );
  OAI22_X1 U6700 ( .A1(n332), .A2(n2897), .B1(n7568), .B2(n2105), .ZN(n6939)
         );
  NAND2_X1 U6701 ( .A1(n1840), .A2(n4105), .ZN(n1972) );
  OAI22_X1 U6702 ( .A1(n6743), .A2(n698), .B1(n6837), .B2(n1436), .ZN(n4105)
         );
  OAI22_X1 U6703 ( .A1(n7257), .A2(n2106), .B1(n349), .B2(n2865), .ZN(n7042)
         );
  OAI22_X1 U6704 ( .A1(n7616), .A2(n2972), .B1(n349), .B2(n2127), .ZN(n7051)
         );
  OAI22_X1 U6705 ( .A1(n7676), .A2(n2197), .B1(n7677), .B2(n2195), .ZN(n5508)
         );
  OAI22_X1 U6706 ( .A1(n6691), .A2(n818), .B1(n6692), .B2(n2085), .ZN(n6923)
         );
  OAI22_X1 U6707 ( .A1(n6790), .A2(n818), .B1(n6882), .B2(n2085), .ZN(n7072)
         );
  OAI22_X1 U6708 ( .A1(n6791), .A2(n818), .B1(n6884), .B2(n2085), .ZN(n7073)
         );
  OAI22_X1 U6709 ( .A1(n6793), .A2(n818), .B1(n6885), .B2(n815), .ZN(n7076) );
  OAI22_X1 U6710 ( .A1(n6794), .A2(n818), .B1(n6887), .B2(n2085), .ZN(n7077)
         );
  OAI22_X1 U6711 ( .A1(n6795), .A2(n818), .B1(n6889), .B2(n2085), .ZN(n7078)
         );
  OAI22_X1 U6712 ( .A1(n6797), .A2(n818), .B1(n6908), .B2(n2085), .ZN(n7080)
         );
  OAI22_X1 U6713 ( .A1(n6798), .A2(n818), .B1(n6906), .B2(n2085), .ZN(n7081)
         );
  OAI22_X1 U6714 ( .A1(n6799), .A2(n818), .B1(n6903), .B2(n2085), .ZN(n7082)
         );
  OAI22_X1 U6715 ( .A1(n6800), .A2(n818), .B1(n6894), .B2(n2085), .ZN(n7083)
         );
  OAI22_X1 U6716 ( .A1(n6801), .A2(n818), .B1(n6915), .B2(n2085), .ZN(n7084)
         );
  OAI22_X1 U6717 ( .A1(n6802), .A2(n818), .B1(n6897), .B2(n2085), .ZN(n7085)
         );
  OAI221_X1 U6718 ( .B1(n7417), .B2(n3180), .C1(n908), .C2(n8284), .A(n3147), 
        .ZN(n8051) );
  INV_X1 U6719 ( .A(n2036), .ZN(n3147) );
  OAI22_X1 U6720 ( .A1(n537), .A2(n7322), .B1(n913), .B2(n6672), .ZN(n2036) );
  OAI221_X1 U6721 ( .B1(n7656), .B2(n3180), .C1(n6658), .C2(n908), .A(n3146), 
        .ZN(n7294) );
  INV_X1 U6722 ( .A(n2174), .ZN(n3146) );
  OAI22_X1 U6723 ( .A1(n537), .A2(n7652), .B1(n913), .B2(n7651), .ZN(n2174) );
  NAND2_X1 U6724 ( .A1(n7306), .A2(n556), .ZN(n559) );
  OAI22_X1 U6725 ( .A1(n4134), .A2(n800), .B1(n7540), .B2(n799), .ZN(n6947) );
  OAI22_X1 U6726 ( .A1(n4126), .A2(n800), .B1(n7635), .B2(n799), .ZN(n7197) );
  OAI22_X1 U6727 ( .A1(n4134), .A2(n2897), .B1(n7569), .B2(n2105), .ZN(n6946)
         );
  OAI22_X1 U6728 ( .A1(n4134), .A2(n2989), .B1(n6710), .B2(n2101), .ZN(n6948)
         );
  OAI22_X1 U6729 ( .A1(n4134), .A2(n2983), .B1(n6711), .B2(n2099), .ZN(n6949)
         );
  OAI22_X1 U6730 ( .A1(n4134), .A2(n2987), .B1(n7551), .B2(n2097), .ZN(n6950)
         );
  OAI22_X1 U6731 ( .A1(n4134), .A2(n2992), .B1(n6712), .B2(n2095), .ZN(n6951)
         );
  OAI22_X1 U6732 ( .A1(n4134), .A2(n2885), .B1(n7621), .B2(n2093), .ZN(n6952)
         );
  OAI22_X1 U6733 ( .A1(n4134), .A2(n2906), .B1(n7610), .B2(n2091), .ZN(n6953)
         );
  OAI22_X1 U6734 ( .A1(n4134), .A2(n2883), .B1(n7323), .B2(n2089), .ZN(n6954)
         );
  OAI22_X1 U6735 ( .A1(n4126), .A2(n2883), .B1(n7639), .B2(n2089), .ZN(n7007)
         );
  OAI22_X1 U6736 ( .A1(n4126), .A2(n2987), .B1(n7636), .B2(n2097), .ZN(n7011)
         );
  OAI22_X1 U6737 ( .A1(n4126), .A2(n2897), .B1(n7634), .B2(n2105), .ZN(n7033)
         );
  OAI22_X1 U6738 ( .A1(n4126), .A2(n2992), .B1(n6773), .B2(n2095), .ZN(n7037)
         );
  OAI22_X1 U6739 ( .A1(n4126), .A2(n2989), .B1(n6775), .B2(n2101), .ZN(n7043)
         );
  OAI22_X1 U6740 ( .A1(n4126), .A2(n2885), .B1(n7637), .B2(n2093), .ZN(n7050)
         );
  OAI22_X1 U6741 ( .A1(n4126), .A2(n2983), .B1(n6778), .B2(n2099), .ZN(n7053)
         );
  OAI22_X1 U6742 ( .A1(n4126), .A2(n2906), .B1(n7638), .B2(n2091), .ZN(n7057)
         );
  NAND2_X1 U6743 ( .A1(n7708), .A2(n2307), .ZN(Knmhu6) );
  NAND2_X1 U6744 ( .A1(n7707), .A2(n2333), .ZN(I5khu6) );
  NOR3_X1 U6745 ( .A1(n528), .A2(n7335), .A3(n7482), .ZN(n2177) );
  NOR2_X1 U6746 ( .A1(n3244), .A2(n7505), .ZN(n3240) );
  NAND4_X1 U6747 ( .A1(n604), .A2(n605), .A3(n606), .A4(n607), .ZN(n7838) );
  OAI211_X1 U6748 ( .C1(n630), .C2(n609), .A(n4028), .B(n7310), .ZN(n606) );
  AOI22_X1 U6749 ( .A1(n4015), .A2(n608), .B1(n609), .B2(n610), .ZN(n607) );
  NOR2_X1 U6750 ( .A1(n4024), .A2(n3142), .ZN(n630) );
  AOI22_X1 U6751 ( .A1(n70), .A2(n3702), .B1(n72), .B2(n73), .ZN(n69) );
  INV_X1 U6752 ( .A(n77), .ZN(n3702) );
  OAI22_X1 U6753 ( .A1(n505), .A2(n4193), .B1(n3123), .B2(n3837), .ZN(n73) );
  AOI21_X1 U6754 ( .B1(n4572), .B2(n7516), .A(n79), .ZN(n77) );
  NAND4_X1 U6755 ( .A1(n6575), .A2(n6578), .A3(n6581), .A4(n6582), .ZN(n5519)
         );
  AOI22_X1 U6756 ( .A1(n7423), .A2(n958), .B1(n959), .B2(n960), .ZN(n951) );
  AND3_X1 U6757 ( .A1(n945), .A2(n7447), .A3(n7437), .ZN(n959) );
  AOI211_X1 U6758 ( .C1(n918), .C2(n923), .A(n152), .B(n3890), .ZN(n960) );
  OAI21_X1 U6759 ( .B1(Jshpw6[4]), .B2(n4146), .A(n965), .ZN(n958) );
  NAND2_X1 U6760 ( .A1(vis_ipsr_o[1]), .A2(n5244), .ZN(n2113) );
  NAND4_X1 U6761 ( .A1(n1558), .A2(n1559), .A3(n1560), .A4(n1561), .ZN(n1557)
         );
  AOI221_X1 U6762 ( .B1(n1562), .B2(n1563), .C1(n1564), .C2(n1565), .A(n1566), 
        .ZN(n1561) );
  AOI222_X1 U6763 ( .A1(n2124), .A2(n529), .B1(n1613), .B2(n7518), .C1(n1584), 
        .C2(n4187), .ZN(n1558) );
  AOI222_X1 U6764 ( .A1(n1576), .A2(n1577), .B1(n1462), .B2(n1578), .C1(n7354), 
        .C2(n1579), .ZN(n1559) );
  NAND4_X1 U6765 ( .A1(n7585), .A2(n7586), .A3(n7587), .A4(n7588), .ZN(n5517)
         );
  AOI21_X1 U6766 ( .B1(n6660), .B2(n903), .A(n4723), .ZN(n5482) );
  NAND3_X1 U6767 ( .A1(n7305), .A2(n3158), .A3(n4752), .ZN(n534) );
  NOR3_X1 U6768 ( .A1(n7482), .A2(n7250), .A3(n7335), .ZN(n4752) );
  AOI22_X1 U6769 ( .A1(n497), .A2(n498), .B1(n499), .B2(n228), .ZN(n494) );
  NAND2_X1 U6770 ( .A1(n2124), .A2(n500), .ZN(n498) );
  OAI211_X1 U6771 ( .C1(n501), .C2(n7259), .A(n4341), .B(n7399), .ZN(n500) );
  OAI211_X1 U6772 ( .C1(n2594), .C2(n1619), .A(n2256), .B(n2698), .ZN(n1617)
         );
  NAND2_X1 U6773 ( .A1(n7399), .A2(n265), .ZN(n1619) );
  AOI21_X1 U6774 ( .B1(n7701), .B2(n903), .A(n4723), .ZN(n5965) );
  NAND4_X1 U6775 ( .A1(n7593), .A2(n7594), .A3(n7595), .A4(n7596), .ZN(n5515)
         );
  OAI22_X1 U6776 ( .A1(n905), .A2(n800), .B1(n7542), .B2(n799), .ZN(n7722) );
  OAI22_X1 U6777 ( .A1(n905), .A2(n3002), .B1(n7442), .B2(n2112), .ZN(n7723)
         );
  OAI22_X1 U6778 ( .A1(n905), .A2(n2123), .B1(n7560), .B2(n2967), .ZN(n7721)
         );
  NAND4_X1 U6779 ( .A1(n7255), .A2(n7357), .A3(n7583), .A4(n7584), .ZN(n5518)
         );
  NAND4_X1 U6780 ( .A1(n7597), .A2(n7598), .A3(n7599), .A4(n7601), .ZN(n5514)
         );
  OAI22_X1 U6781 ( .A1(n7316), .A2(n788), .B1(n6572), .B2(n794), .ZN(n7221) );
  AOI21_X1 U6782 ( .B1(n7354), .B2(n1679), .A(n4187), .ZN(n1678) );
  OAI211_X1 U6783 ( .C1(n4672), .C2(n5002), .A(n3701), .B(n1682), .ZN(n1679)
         );
  AOI21_X1 U6784 ( .B1(n1683), .B2(n7514), .A(n7381), .ZN(n1682) );
  NAND4_X1 U6785 ( .A1(n7602), .A2(n7604), .A3(n7645), .A4(n7669), .ZN(n5513)
         );
  OAI22_X1 U6786 ( .A1(n6815), .A2(n847), .B1(n6906), .B2(n836), .ZN(n7100) );
  OAI22_X1 U6787 ( .A1(n6868), .A2(n863), .B1(n6906), .B2(n2077), .ZN(n7170)
         );
  OAI22_X1 U6788 ( .A1(n6892), .A2(n854), .B1(n6906), .B2(n2079), .ZN(n7191)
         );
  NAND4_X1 U6789 ( .A1(n7684), .A2(n7689), .A3(n7696), .A4(n3645), .ZN(n5512)
         );
  OAI22_X1 U6790 ( .A1(n6615), .A2(n788), .B1(n6906), .B2(n794), .ZN(n7226) );
  OAI22_X1 U6791 ( .A1(n1515), .A2(n841), .B1(n6885), .B2(n836), .ZN(n7095) );
  OAI22_X1 U6792 ( .A1(n6811), .A2(n841), .B1(n6887), .B2(n836), .ZN(n7096) );
  OAI22_X1 U6793 ( .A1(n1119), .A2(n857), .B1(n6885), .B2(n855), .ZN(n7165) );
  OAI22_X1 U6794 ( .A1(n6864), .A2(n857), .B1(n6887), .B2(n2077), .ZN(n7166)
         );
  OAI22_X1 U6795 ( .A1(n1256), .A2(n850), .B1(n6885), .B2(n848), .ZN(n7187) );
  OAI22_X1 U6796 ( .A1(n6888), .A2(n850), .B1(n6887), .B2(n2079), .ZN(n7188)
         );
  OAI22_X1 U6797 ( .A1(n7420), .A2(n788), .B1(n6887), .B2(n794), .ZN(n7234) );
  OAI22_X1 U6798 ( .A1(n7416), .A2(n2155), .B1(n6885), .B2(n791), .ZN(n7244)
         );
  OAI21_X1 U6799 ( .B1(n7564), .B2(n2197), .A(n5958), .ZN(n5957) );
  NAND3_X1 U6800 ( .A1(n2969), .A2(n4454), .A3(n5483), .ZN(n5958) );
  NAND3_X1 U6801 ( .A1(n1607), .A2(n2952), .A3(n7523), .ZN(n1686) );
  OAI22_X1 U6802 ( .A1(n6726), .A2(n818), .B1(n6727), .B2(n815), .ZN(n6968) );
  OAI22_X1 U6803 ( .A1(n7431), .A2(n788), .B1(n6727), .B2(n791), .ZN(n7243) );
  OAI22_X1 U6804 ( .A1(n6687), .A2(n857), .B1(n6692), .B2(n855), .ZN(n6919) );
  OAI22_X1 U6805 ( .A1(n6688), .A2(n850), .B1(n6692), .B2(n848), .ZN(n6920) );
  OAI22_X1 U6806 ( .A1(n6736), .A2(n863), .B1(n6741), .B2(n855), .ZN(n6986) );
  OAI22_X1 U6807 ( .A1(n6737), .A2(n854), .B1(n6741), .B2(n848), .ZN(n6987) );
  OAI22_X1 U6808 ( .A1(n6738), .A2(n847), .B1(n6741), .B2(n2081), .ZN(n6988)
         );
  OAI22_X1 U6809 ( .A1(n6740), .A2(n818), .B1(n6741), .B2(n815), .ZN(n6990) );
  OAI22_X1 U6810 ( .A1(n6720), .A2(n857), .B1(n6904), .B2(n855), .ZN(n6962) );
  OAI22_X1 U6811 ( .A1(n6721), .A2(n850), .B1(n6904), .B2(n848), .ZN(n6963) );
  OAI22_X1 U6812 ( .A1(n6722), .A2(n841), .B1(n6904), .B2(n2081), .ZN(n6964)
         );
  OAI22_X1 U6813 ( .A1(n6724), .A2(n818), .B1(n6904), .B2(n815), .ZN(n6966) );
  OAI22_X1 U6814 ( .A1(n6744), .A2(n863), .B1(n6750), .B2(n855), .ZN(n6993) );
  OAI22_X1 U6815 ( .A1(n6745), .A2(n854), .B1(n6750), .B2(n848), .ZN(n6994) );
  OAI22_X1 U6816 ( .A1(n6746), .A2(n847), .B1(n6750), .B2(n2081), .ZN(n6995)
         );
  OAI22_X1 U6817 ( .A1(n6748), .A2(n824), .B1(n6750), .B2(n815), .ZN(n6997) );
  OAI22_X1 U6818 ( .A1(n6713), .A2(n863), .B1(n6718), .B2(n2077), .ZN(n6956)
         );
  OAI22_X1 U6819 ( .A1(n6714), .A2(n854), .B1(n6718), .B2(n2079), .ZN(n6957)
         );
  OAI22_X1 U6820 ( .A1(n6717), .A2(n818), .B1(n6718), .B2(n2085), .ZN(n6960)
         );
  OAI22_X1 U6821 ( .A1(n6788), .A2(n824), .B1(n6905), .B2(n815), .ZN(n7070) );
  OAI22_X1 U6822 ( .A1(n6807), .A2(n847), .B1(n6905), .B2(n2081), .ZN(n7090)
         );
  OAI22_X1 U6823 ( .A1(n6860), .A2(n863), .B1(n6905), .B2(n855), .ZN(n7160) );
  OAI22_X1 U6824 ( .A1(n6880), .A2(n854), .B1(n6905), .B2(n848), .ZN(n7182) );
  OAI22_X1 U6825 ( .A1(n7651), .A2(n788), .B1(n6692), .B2(n794), .ZN(n7227) );
  OAI22_X1 U6826 ( .A1(n6609), .A2(n788), .B1(n6741), .B2(n794), .ZN(n7238) );
  NAND4_X1 U6827 ( .A1(n611), .A2(n3204), .A3(n612), .A4(n613), .ZN(n608) );
  NAND3_X1 U6828 ( .A1(n626), .A2(n4027), .A3(n3197), .ZN(n611) );
  OAI21_X1 U6829 ( .B1(n621), .B2(n622), .A(n4022), .ZN(n612) );
  AOI211_X1 U6830 ( .C1(n586), .C2(n7318), .A(n603), .B(n614), .ZN(n613) );
  OAI22_X1 U6831 ( .A1(n6612), .A2(n788), .B1(n6904), .B2(n794), .ZN(n7232) );
  OAI22_X1 U6832 ( .A1(n6621), .A2(n2155), .B1(n6750), .B2(n791), .ZN(n7247)
         );
  OAI22_X1 U6833 ( .A1(n6611), .A2(n788), .B1(n6718), .B2(n791), .ZN(n7223) );
  OAI22_X1 U6834 ( .A1(n6614), .A2(n788), .B1(n6905), .B2(n794), .ZN(n7216) );
  OAI22_X1 U6835 ( .A1(n6809), .A2(n841), .B1(n6882), .B2(n836), .ZN(n7092) );
  OAI22_X1 U6836 ( .A1(n6862), .A2(n857), .B1(n6882), .B2(n2077), .ZN(n7162)
         );
  OAI22_X1 U6837 ( .A1(n6883), .A2(n850), .B1(n6882), .B2(n2079), .ZN(n7184)
         );
  OAI22_X1 U6838 ( .A1(n6817), .A2(n841), .B1(n6894), .B2(n836), .ZN(n7102) );
  OAI22_X1 U6839 ( .A1(n6870), .A2(n857), .B1(n6894), .B2(n2077), .ZN(n7172)
         );
  OAI22_X1 U6840 ( .A1(n6895), .A2(n850), .B1(n6894), .B2(n2079), .ZN(n7193)
         );
  OAI22_X1 U6841 ( .A1(n7346), .A2(n2155), .B1(n6882), .B2(n791), .ZN(n7217)
         );
  OAI22_X1 U6842 ( .A1(n6625), .A2(n788), .B1(n6894), .B2(n794), .ZN(n7220) );
  OAI22_X1 U6843 ( .A1(n7468), .A2(n841), .B1(n6897), .B2(n836), .ZN(n7104) );
  OAI22_X1 U6844 ( .A1(n7470), .A2(n857), .B1(n6897), .B2(n2077), .ZN(n7173)
         );
  OAI22_X1 U6845 ( .A1(n7472), .A2(n850), .B1(n6897), .B2(n2079), .ZN(n7195)
         );
  OAI22_X1 U6846 ( .A1(n700), .A2(n800), .B1(n7543), .B2(n799), .ZN(n7719) );
  OAI22_X1 U6847 ( .A1(n7409), .A2(n788), .B1(n6897), .B2(n794), .ZN(n7233) );
  OAI22_X1 U6848 ( .A1(n700), .A2(n3002), .B1(n7570), .B2(n2112), .ZN(n7720)
         );
  OAI22_X1 U6849 ( .A1(n700), .A2(n2123), .B1(n7559), .B2(n2967), .ZN(n7718)
         );
  OAI22_X1 U6850 ( .A1(n6786), .A2(n824), .B1(n6907), .B2(n815), .ZN(n7068) );
  OAI22_X1 U6851 ( .A1(n6805), .A2(n847), .B1(n6907), .B2(n2081), .ZN(n7088)
         );
  OAI22_X1 U6852 ( .A1(n6858), .A2(n863), .B1(n6907), .B2(n855), .ZN(n7158) );
  OAI22_X1 U6853 ( .A1(n6878), .A2(n854), .B1(n6907), .B2(n848), .ZN(n7180) );
  OAI22_X1 U6854 ( .A1(n6729), .A2(n857), .B1(n6912), .B2(n855), .ZN(n6970) );
  OAI22_X1 U6855 ( .A1(n6730), .A2(n850), .B1(n6912), .B2(n848), .ZN(n6971) );
  OAI22_X1 U6856 ( .A1(n6731), .A2(n841), .B1(n6912), .B2(n2081), .ZN(n6972)
         );
  OAI22_X1 U6857 ( .A1(n6733), .A2(n824), .B1(n6912), .B2(n815), .ZN(n6974) );
  OAI22_X1 U6858 ( .A1(n6816), .A2(n841), .B1(n6903), .B2(n836), .ZN(n7101) );
  OAI22_X1 U6859 ( .A1(n6869), .A2(n857), .B1(n6903), .B2(n2077), .ZN(n7171)
         );
  OAI22_X1 U6860 ( .A1(n6893), .A2(n850), .B1(n6903), .B2(n2079), .ZN(n7192)
         );
  OAI22_X1 U6861 ( .A1(n6787), .A2(n824), .B1(n7653), .B2(n815), .ZN(n7069) );
  OAI22_X1 U6862 ( .A1(n6806), .A2(n847), .B1(n7653), .B2(n836), .ZN(n7089) );
  OAI22_X1 U6863 ( .A1(n6859), .A2(n863), .B1(n7653), .B2(n855), .ZN(n7159) );
  OAI22_X1 U6864 ( .A1(n6879), .A2(n854), .B1(n7653), .B2(n848), .ZN(n7181) );
  OAI22_X1 U6865 ( .A1(n6610), .A2(n2155), .B1(n6907), .B2(n791), .ZN(n7248)
         );
  OAI22_X1 U6866 ( .A1(n6623), .A2(n788), .B1(n6912), .B2(n794), .ZN(n7230) );
  OAI22_X1 U6867 ( .A1(n6613), .A2(n788), .B1(n6903), .B2(n794), .ZN(n7241) );
  OAI22_X1 U6868 ( .A1(n7483), .A2(n841), .B1(n6884), .B2(n836), .ZN(n7093) );
  OAI22_X1 U6869 ( .A1(n6818), .A2(n841), .B1(n6915), .B2(n836), .ZN(n7103) );
  OAI22_X1 U6870 ( .A1(n7486), .A2(n857), .B1(n6884), .B2(n2077), .ZN(n7163)
         );
  OAI22_X1 U6871 ( .A1(n7485), .A2(n850), .B1(n6884), .B2(n2079), .ZN(n7185)
         );
  OAI22_X1 U6872 ( .A1(n6896), .A2(n850), .B1(n6915), .B2(n2079), .ZN(n7194)
         );
  OAI22_X1 U6873 ( .A1(n6916), .A2(n857), .B1(n6915), .B2(n2077), .ZN(n7212)
         );
  OAI22_X1 U6874 ( .A1(n7652), .A2(n788), .B1(n7653), .B2(n794), .ZN(Qixhu6)
         );
  OAI22_X1 U6875 ( .A1(n7334), .A2(n2155), .B1(n6884), .B2(n791), .ZN(n7242)
         );
  OAI22_X1 U6876 ( .A1(n6624), .A2(n2155), .B1(n6915), .B2(n791), .ZN(n7246)
         );
  OAI221_X1 U6877 ( .B1(n3219), .B2(n548), .C1(n6670), .C2(n913), .A(n665), 
        .ZN(n7841) );
  AOI21_X1 U6878 ( .B1(n666), .B2(n556), .A(n663), .ZN(n665) );
  OAI22_X1 U6879 ( .A1(n7440), .A2(n3007), .B1(n3012), .B2(n2446), .ZN(P0xhu6)
         );
  OAI22_X1 U6880 ( .A1(n6694), .A2(n857), .B1(n6902), .B2(n2077), .ZN(n6925)
         );
  OAI22_X1 U6881 ( .A1(n6695), .A2(n850), .B1(n6902), .B2(n2079), .ZN(n6926)
         );
  OAI22_X1 U6882 ( .A1(n6698), .A2(n824), .B1(n6902), .B2(n2085), .ZN(n6929)
         );
  OAI22_X1 U6883 ( .A1(n6789), .A2(n824), .B1(n6900), .B2(n815), .ZN(n7071) );
  OAI22_X1 U6884 ( .A1(n6808), .A2(n847), .B1(n6900), .B2(n836), .ZN(n7091) );
  OAI22_X1 U6885 ( .A1(n6812), .A2(n841), .B1(n6889), .B2(n836), .ZN(n7097) );
  OAI22_X1 U6886 ( .A1(n6861), .A2(n863), .B1(n6900), .B2(n855), .ZN(n7161) );
  OAI22_X1 U6887 ( .A1(n6865), .A2(n857), .B1(n6889), .B2(n2077), .ZN(n7167)
         );
  OAI22_X1 U6888 ( .A1(n6881), .A2(n850), .B1(n6900), .B2(n2079), .ZN(n7183)
         );
  OAI22_X1 U6889 ( .A1(n6890), .A2(n850), .B1(n6889), .B2(n2079), .ZN(n7189)
         );
  OAI22_X1 U6890 ( .A1(n6785), .A2(n824), .B1(n6901), .B2(n815), .ZN(n7067) );
  OAI22_X1 U6891 ( .A1(n6804), .A2(n847), .B1(n6901), .B2(n2081), .ZN(n7087)
         );
  OAI22_X1 U6892 ( .A1(n6857), .A2(n863), .B1(n6901), .B2(n855), .ZN(n7157) );
  OAI22_X1 U6893 ( .A1(n6877), .A2(n854), .B1(n6901), .B2(n848), .ZN(n7179) );
  OAI22_X1 U6894 ( .A1(n6672), .A2(n2155), .B1(n6902), .B2(n794), .ZN(n7231)
         );
  OAI22_X1 U6895 ( .A1(n6703), .A2(n857), .B1(n6708), .B2(n2077), .ZN(n6940)
         );
  OAI22_X1 U6896 ( .A1(n6704), .A2(n850), .B1(n6708), .B2(n2079), .ZN(n6941)
         );
  OAI22_X1 U6897 ( .A1(n6707), .A2(n818), .B1(n6708), .B2(n2085), .ZN(n6944)
         );
  OAI22_X1 U6898 ( .A1(n6751), .A2(n863), .B1(n6756), .B2(n855), .ZN(n7001) );
  OAI22_X1 U6899 ( .A1(n6752), .A2(n854), .B1(n6756), .B2(n848), .ZN(n7002) );
  OAI22_X1 U6900 ( .A1(n6753), .A2(n847), .B1(n6756), .B2(n2081), .ZN(n7003)
         );
  OAI22_X1 U6901 ( .A1(n6755), .A2(n824), .B1(n6756), .B2(n815), .ZN(n7005) );
  OAI22_X1 U6902 ( .A1(n6761), .A2(n863), .B1(n6766), .B2(n855), .ZN(n7016) );
  OAI22_X1 U6903 ( .A1(n6762), .A2(n854), .B1(n6766), .B2(n848), .ZN(n7017) );
  OAI22_X1 U6904 ( .A1(n6763), .A2(n847), .B1(n6766), .B2(n2081), .ZN(n7018)
         );
  OAI22_X1 U6905 ( .A1(n6765), .A2(n824), .B1(n6766), .B2(n815), .ZN(n7020) );
  OAI22_X1 U6906 ( .A1(n6796), .A2(n824), .B1(n6875), .B2(n2085), .ZN(n7079)
         );
  OAI22_X1 U6907 ( .A1(n6813), .A2(n841), .B1(n6875), .B2(n836), .ZN(n7098) );
  OAI22_X1 U6908 ( .A1(n6814), .A2(n841), .B1(n6908), .B2(n836), .ZN(n7099) );
  OAI22_X1 U6909 ( .A1(n6866), .A2(n857), .B1(n6875), .B2(n2077), .ZN(n7168)
         );
  OAI22_X1 U6910 ( .A1(n6867), .A2(n857), .B1(n6908), .B2(n2077), .ZN(n7169)
         );
  OAI22_X1 U6911 ( .A1(n6876), .A2(n854), .B1(n6875), .B2(n848), .ZN(n7178) );
  OAI22_X1 U6912 ( .A1(n6891), .A2(n850), .B1(n6908), .B2(n2079), .ZN(n7190)
         );
  OAI22_X1 U6913 ( .A1(n6779), .A2(n863), .B1(n6911), .B2(n855), .ZN(n7061) );
  OAI22_X1 U6914 ( .A1(n6780), .A2(n854), .B1(n6911), .B2(n848), .ZN(n7062) );
  OAI22_X1 U6915 ( .A1(n6781), .A2(n847), .B1(n6911), .B2(n2081), .ZN(n7063)
         );
  OAI22_X1 U6916 ( .A1(n6783), .A2(n824), .B1(n6911), .B2(n815), .ZN(n7065) );
  OAI22_X1 U6917 ( .A1(n7477), .A2(n788), .B1(n6900), .B2(n794), .ZN(n7215) );
  OAI22_X1 U6918 ( .A1(n7322), .A2(n788), .B1(n6889), .B2(n794), .ZN(n7239) );
  OAI22_X1 U6919 ( .A1(n6671), .A2(n788), .B1(n6901), .B2(n791), .ZN(n7222) );
  OAI22_X1 U6920 ( .A1(n6617), .A2(n2155), .B1(n6708), .B2(n791), .ZN(n7245)
         );
  OAI22_X1 U6921 ( .A1(n6620), .A2(n788), .B1(n6756), .B2(n794), .ZN(n7237) );
  OAI22_X1 U6922 ( .A1(n6616), .A2(n2155), .B1(n6766), .B2(n794), .ZN(n7235)
         );
  OAI22_X1 U6923 ( .A1(n6619), .A2(n788), .B1(n6875), .B2(n794), .ZN(n7229) );
  OAI22_X1 U6924 ( .A1(n6618), .A2(n2155), .B1(n6908), .B2(n791), .ZN(n7219)
         );
  OAI22_X1 U6925 ( .A1(n7337), .A2(n2155), .B1(n6911), .B2(n791), .ZN(n7225)
         );
  AND2_X1 U6926 ( .A1(n7363), .A2(n4395), .ZN(n1857) );
  AOI21_X1 U6927 ( .B1(n2507), .B2(vis_apsr_o[1]), .A(n470), .ZN(n2945) );
  OAI22_X1 U6928 ( .A1(n2679), .A2(n800), .B1(n7367), .B2(n799), .ZN(n7203) );
  OAI22_X1 U6929 ( .A1(n2686), .A2(n800), .B1(n7379), .B2(n2103), .ZN(n7202)
         );
  OAI22_X1 U6930 ( .A1(n2689), .A2(n800), .B1(n7277), .B2(n799), .ZN(n6955) );
  OAI22_X1 U6931 ( .A1(n2691), .A2(n800), .B1(n7289), .B2(n799), .ZN(n7205) );
  AOI21_X1 U6932 ( .B1(n5510), .B2(n5511), .A(n2825), .ZN(n5509) );
  NOR4_X1 U6933 ( .A1(n5516), .A2(n5517), .A3(n5518), .A4(n5519), .ZN(n5510)
         );
  NOR4_X1 U6934 ( .A1(n5512), .A2(n5513), .A3(n5514), .A4(n5515), .ZN(n5511)
         );
  NAND4_X1 U6935 ( .A1(n7589), .A2(n7590), .A3(n7591), .A4(n7592), .ZN(n5516)
         );
  AND2_X1 U6936 ( .A1(n1287), .A2(n7451), .ZN(n1969) );
  OAI22_X1 U6937 ( .A1(n7321), .A2(n3136), .B1(n7293), .B2(n2159), .ZN(Tgxhu6)
         );
  OAI22_X1 U6938 ( .A1(n7478), .A2(n2665), .B1(n3133), .B2(n3770), .ZN(Isxhu6)
         );
  OAI21_X1 U6939 ( .B1(n3771), .B2(n3772), .A(n3884), .ZN(n3770) );
  NOR3_X1 U6940 ( .A1(n7477), .A2(n7322), .A3(n7337), .ZN(n3771) );
  AOI21_X1 U6941 ( .B1(n513), .B2(n514), .A(n515), .ZN(n512) );
  NOR3_X1 U6942 ( .A1(n2698), .A2(n7433), .A3(n1967), .ZN(n515) );
  OAI22_X1 U6943 ( .A1(n2665), .A2(n4044), .B1(n3772), .B2(n3133), .ZN(Avxhu6)
         );
  OAI22_X1 U6944 ( .A1(n7347), .A2(n3136), .B1(n7346), .B2(n2159), .ZN(Fgxhu6)
         );
  OAI22_X1 U6945 ( .A1(n2664), .A2(n800), .B1(n7361), .B2(n799), .ZN(n7204) );
  OAI22_X1 U6946 ( .A1(n2667), .A2(n800), .B1(n7390), .B2(n799), .ZN(n7201) );
  OAI22_X1 U6947 ( .A1(n6608), .A2(n3136), .B1(n7409), .B2(n2159), .ZN(n7251)
         );
  OAI22_X1 U6948 ( .A1(n2776), .A2(n800), .B1(n7686), .B2(n799), .ZN(n7028) );
  OAI22_X1 U6949 ( .A1(n1831), .A2(n800), .B1(n7351), .B2(n799), .ZN(n7030) );
  OAI22_X1 U6950 ( .A1(n7656), .A2(n3136), .B1(n7652), .B2(n2159), .ZN(Mgxhu6)
         );
  OAI22_X1 U6951 ( .A1(n1831), .A2(n3002), .B1(n6760), .B2(n2112), .ZN(n7015)
         );
  OAI22_X1 U6952 ( .A1(n2776), .A2(n2123), .B1(n7688), .B2(n2967), .ZN(n7029)
         );
  OAI22_X1 U6953 ( .A1(n339), .A2(n800), .B1(n7698), .B2(n799), .ZN(n7198) );
  OAI22_X1 U6954 ( .A1(n335), .A2(n800), .B1(n7402), .B2(n799), .ZN(n7200) );
  OAI22_X1 U6955 ( .A1(n339), .A2(n892), .B1(n7697), .B2(n1853), .ZN(n7978) );
  NOR2_X1 U6956 ( .A1(n703), .A2(n339), .ZN(n1853) );
  OAI22_X1 U6957 ( .A1(n335), .A2(n892), .B1(n6635), .B2(n1771), .ZN(n7949) );
  NOR2_X1 U6958 ( .A1(n703), .A2(n335), .ZN(n1771) );
  OAI22_X1 U6959 ( .A1(n7293), .A2(n3133), .B1(n7320), .B2(n2665), .ZN(Sqxhu6)
         );
  OAI211_X1 U6960 ( .C1(n7396), .C2(n908), .A(n3190), .B(n3153), .ZN(n8041) );
  INV_X1 U6961 ( .A(n2017), .ZN(n3153) );
  OAI22_X1 U6962 ( .A1(n928), .A2(n6621), .B1(n917), .B2(n6620), .ZN(n2017) );
  OAI22_X1 U6963 ( .A1(n4028), .A2(n3202), .B1(n583), .B2(n548), .ZN(n7837) );
  NOR4_X1 U6964 ( .A1(n584), .A2(n585), .A3(n586), .A4(n3216), .ZN(n583) );
  OAI221_X1 U6965 ( .B1(n597), .B2(n601), .C1(n7314), .C2(n3215), .A(n3143), 
        .ZN(n584) );
  OAI21_X1 U6966 ( .B1(n7313), .B2(n587), .A(n588), .ZN(n585) );
  OAI22_X1 U6967 ( .A1(n7415), .A2(n3007), .B1(n4052), .B2(n2446), .ZN(I0xhu6)
         );
  OAI211_X1 U6968 ( .C1(n7650), .C2(n908), .A(n3190), .B(n3006), .ZN(n8047) );
  INV_X1 U6969 ( .A(n2029), .ZN(n3006) );
  OAI22_X1 U6970 ( .A1(n537), .A2(n7651), .B1(n917), .B2(n7346), .ZN(n2029) );
  OAI211_X1 U6971 ( .C1(n7662), .C2(n908), .A(n3190), .B(n3151), .ZN(n8044) );
  INV_X1 U6972 ( .A(n2023), .ZN(n3151) );
  OAI22_X1 U6973 ( .A1(n537), .A2(n6611), .B1(n917), .B2(n6610), .ZN(n2023) );
  OAI211_X1 U6974 ( .C1(n7659), .C2(n908), .A(n3190), .B(n3154), .ZN(n8020) );
  INV_X1 U6975 ( .A(n1995), .ZN(n3154) );
  OAI22_X1 U6976 ( .A1(n928), .A2(n6623), .B1(n917), .B2(n6625), .ZN(n1995) );
  OAI211_X1 U6977 ( .C1(n7449), .C2(n908), .A(n3190), .B(n3045), .ZN(n8042) );
  INV_X1 U6978 ( .A(n2019), .ZN(n3045) );
  OAI22_X1 U6979 ( .A1(n537), .A2(n6619), .B1(n917), .B2(n6618), .ZN(n2019) );
  OAI211_X1 U6980 ( .C1(n7386), .C2(n908), .A(n3190), .B(n3152), .ZN(n8043) );
  INV_X1 U6981 ( .A(n2021), .ZN(n3152) );
  OAI22_X1 U6982 ( .A1(n537), .A2(n6615), .B1(n917), .B2(n6614), .ZN(n2021) );
  OAI211_X1 U6983 ( .C1(n7665), .C2(n908), .A(n3190), .B(n3150), .ZN(n8045) );
  INV_X1 U6984 ( .A(n2025), .ZN(n3150) );
  OAI22_X1 U6985 ( .A1(n537), .A2(n6610), .B1(n917), .B2(n6609), .ZN(n2025) );
  OAI211_X1 U6986 ( .C1(n7413), .C2(n908), .A(n3190), .B(n3149), .ZN(n8046) );
  INV_X1 U6987 ( .A(n2027), .ZN(n3149) );
  OAI22_X1 U6988 ( .A1(n537), .A2(n6624), .B1(n917), .B2(n7652), .ZN(n2027) );
  OAI22_X1 U6989 ( .A1(n7317), .A2(n2155), .B1(n6592), .B2(n794), .ZN(n7236)
         );
  OAI22_X1 U6991 ( .A1(n2657), .A2(n892), .B1(n7574), .B2(n1816), .ZN(n7965)
         );
  NOR2_X1 U6992 ( .A1(n703), .A2(n2657), .ZN(n1816) );
  OAI22_X1 U6993 ( .A1(n2653), .A2(n800), .B1(n7365), .B2(n799), .ZN(n6999) );
  OAI22_X1 U6994 ( .A1(n2655), .A2(n800), .B1(n7327), .B2(n799), .ZN(n7000) );
  OAI22_X1 U6995 ( .A1(n2654), .A2(n800), .B1(n7275), .B2(n799), .ZN(n7022) );
  OAI22_X1 U6996 ( .A1(n2657), .A2(n800), .B1(n7287), .B2(n2103), .ZN(n7206)
         );
  OAI22_X1 U6997 ( .A1(n2653), .A2(n892), .B1(n6633), .B2(n1776), .ZN(n7951)
         );
  NOR2_X1 U6998 ( .A1(n891), .A2(n2653), .ZN(n1776) );
  OAI22_X1 U6999 ( .A1(n2655), .A2(n892), .B1(n6630), .B2(n1792), .ZN(n7956)
         );
  NOR2_X1 U7000 ( .A1(n891), .A2(n2655), .ZN(n1792) );
  OAI22_X1 U7001 ( .A1(n2654), .A2(n892), .B1(n6629), .B2(n1806), .ZN(n7961)
         );
  NOR2_X1 U7002 ( .A1(n891), .A2(n2654), .ZN(n1806) );
  OAI21_X1 U7003 ( .B1(n2455), .B2(n57), .A(n1455), .ZN(n2452) );
  NOR3_X1 U7004 ( .A1(n1706), .A2(n237), .A3(n7400), .ZN(n2455) );
  NAND2_X1 U7005 ( .A1(n1274), .A2(n7411), .ZN(n1083) );
  OAI22_X1 U7006 ( .A1(n7253), .A2(n788), .B1(n6872), .B2(n791), .ZN(n7228) );
  OAI22_X1 U7007 ( .A1(n7439), .A2(n788), .B1(n6898), .B2(n794), .ZN(n7218) );
  OAI22_X1 U7008 ( .A1(n7293), .A2(n788), .B1(n6910), .B2(n791), .ZN(n7224) );
  OAI22_X1 U7009 ( .A1(n3769), .A2(n800), .B1(n7691), .B2(n799), .ZN(n7031) );
  OAI22_X1 U7010 ( .A1(n4072), .A2(n800), .B1(n7338), .B2(n799), .ZN(n7210) );
  OAI211_X1 U7011 ( .C1(n531), .C2(n532), .A(n533), .B(n534), .ZN(n7832) );
  OAI21_X1 U7012 ( .B1(n7439), .B2(n535), .A(n3233), .ZN(n533) );
  OAI21_X1 U7013 ( .B1(n5946), .B2(n538), .A(n4650), .ZN(n5783) );
  AOI21_X1 U7014 ( .B1(n7703), .B2(n7626), .A(n508), .ZN(n5946) );
  OAI22_X1 U7015 ( .A1(n6622), .A2(n2160), .B1(n554), .B2(n3145), .ZN(n7252)
         );
  INV_X1 U7016 ( .A(n2160), .ZN(n3145) );
  NOR3_X1 U7017 ( .A1(n528), .A2(n7318), .A3(n3156), .ZN(n2160) );
  OAI21_X1 U7018 ( .B1(n2644), .B2(n892), .A(n1850), .ZN(n7977) );
  OAI21_X1 U7019 ( .B1(n891), .B2(n2644), .A(n8152), .ZN(n1850) );
  OAI21_X1 U7020 ( .B1(n6631), .B2(n4723), .A(n903), .ZN(n4722) );
  INV_X1 U7021 ( .A(n962), .ZN(n3890) );
  OAI21_X1 U7022 ( .B1(n920), .B2(n939), .A(n7423), .ZN(n962) );
  OAI21_X1 U7023 ( .B1(n344), .B2(n892), .A(n1784), .ZN(n7953) );
  OAI21_X1 U7024 ( .B1(n891), .B2(n344), .A(n8140), .ZN(n1784) );
  NAND3_X1 U7025 ( .A1(n1482), .A2(n3851), .A3(n4462), .ZN(n4461) );
  OAI21_X1 U7026 ( .B1(n4463), .B2(n4464), .A(n3981), .ZN(n4462) );
  NOR3_X1 U7027 ( .A1(n3763), .A2(n7400), .A3(n7530), .ZN(n4463) );
  NAND3_X1 U7028 ( .A1(n3701), .A2(n270), .A3(n2580), .ZN(n2578) );
  AOI211_X1 U7029 ( .C1(n2581), .C2(n1592), .A(n4554), .B(n2583), .ZN(n2580)
         );
  NOR2_X1 U7030 ( .A1(n7518), .A2(n5042), .ZN(n2581) );
  INV_X1 U7031 ( .A(n1495), .ZN(n4554) );
  NAND2_X1 U7032 ( .A1(n556), .A2(n2162), .ZN(n554) );
  NAND4_X1 U7033 ( .A1(n4136), .A2(n3127), .A3(n2165), .A4(n2166), .ZN(n2162)
         );
  AOI21_X1 U7034 ( .B1(n528), .B2(n4138), .A(n2168), .ZN(n2166) );
  NAND2_X1 U7035 ( .A1(n7363), .A2(n7534), .ZN(n3288) );
  OAI21_X1 U7036 ( .B1(n4072), .B2(n894), .A(n1824), .ZN(n7968) );
  OAI21_X1 U7037 ( .B1(n703), .B2(n4072), .A(n8281), .ZN(n1824) );
  OAI22_X1 U7038 ( .A1(n4018), .A2(n579), .B1(n7417), .B2(n580), .ZN(n7836) );
  NOR2_X1 U7039 ( .A1(n7416), .A2(n535), .ZN(n580) );
  AND2_X1 U7040 ( .A1(\add_3107/B[1] ), .A2(Tnhpw6[0]), .ZN(n408) );
  OR2_X1 U7041 ( .A1(n988), .A2(n7412), .ZN(n420) );
  XNOR2_X1 U7042 ( .A(n6675), .B(n791), .ZN(n7830) );
  OR4_X1 U7043 ( .A1(n5564), .A2(n426), .A3(n7626), .A4(n267), .ZN(n5577) );
  AND2_X1 U7044 ( .A1(n5978), .A2(n7371), .ZN(n5972) );
  OAI21_X1 U7045 ( .B1(n6597), .B2(n791), .A(n2156), .ZN(n7240) );
  OAI21_X1 U7046 ( .B1(n2157), .B2(n6596), .A(n791), .ZN(n2156) );
  OAI21_X1 U7047 ( .B1(n7479), .B2(n791), .A(n2359), .ZN(Xpxhu6) );
  OR3_X1 U7048 ( .A1(n2157), .A2(n7478), .A3(n788), .ZN(n2359) );
  NOR2_X1 U7049 ( .A1(n6803), .A2(n2439), .ZN(Wbkhu6) );
  OAI211_X1 U7050 ( .C1(n524), .C2(n4573), .A(n4574), .B(n4575), .ZN(n4530) );
  AOI21_X1 U7051 ( .B1(n2742), .B2(n7283), .A(n4583), .ZN(n4573) );
  NAND3_X1 U7052 ( .A1(n1642), .A2(n538), .A3(n4582), .ZN(n4574) );
  NOR2_X1 U7053 ( .A1(n4576), .A2(n2935), .ZN(n4575) );
  NOR2_X1 U7054 ( .A1(n6856), .A2(n2439), .ZN(Ttmhu6) );
  OR4_X1 U7055 ( .A1(n3114), .A2(n4261), .A3(n3083), .A4(n7400), .ZN(n4384) );
  NAND3_X1 U7056 ( .A1(n1451), .A2(n1452), .A3(n1453), .ZN(n1444) );
  NAND4_X1 U7057 ( .A1(n435), .A2(n1454), .A3(n1455), .A4(n433), .ZN(n1453) );
  NAND4_X1 U7058 ( .A1(n1456), .A2(n417), .A3(n7433), .A4(n1457), .ZN(n1451)
         );
  NAND3_X1 U7059 ( .A1(n1433), .A2(n2548), .A3(n225), .ZN(n7940) );
  OR3_X1 U7060 ( .A1(n3710), .A2(n6653), .A3(n1435), .ZN(n1433) );
  INV_X1 U7061 ( .A(n1436), .ZN(n3710) );
  AND4_X1 U7062 ( .A1(n7309), .A2(n556), .A3(n4015), .A4(n4750), .ZN(n2784) );
  NOR2_X1 U7063 ( .A1(n3144), .A2(n3212), .ZN(n4750) );
  AND2_X1 U7064 ( .A1(Jshpw6[7]), .A2(n425), .ZN(n421) );
  AND2_X1 U7065 ( .A1(Jshpw6[4]), .A2(n424), .ZN(n422) );
  AND2_X1 U7066 ( .A1(Jshpw6[5]), .A2(n422), .ZN(n423) );
  AND2_X1 U7067 ( .A1(Tnhpw6[3]), .A2(\add_3107/carry[4] ), .ZN(n424) );
  AND2_X1 U7068 ( .A1(Jshpw6[6]), .A2(n423), .ZN(n425) );
  NAND2_X1 U7069 ( .A1(n7452), .A2(n7453), .ZN(n2297) );
  OR3_X1 U7070 ( .A1(n3259), .A2(n6910), .A3(n2446), .ZN(n2850) );
  OR3_X1 U7071 ( .A1(n1958), .A2(n4223), .A3(n2273), .ZN(n67) );
  AOI21_X1 U7072 ( .B1(n4672), .B2(n1594), .A(n7510), .ZN(n4223) );
  NAND2_X1 U7073 ( .A1(n6873), .A2(n6874), .ZN(n2264) );
  AOI211_X1 U7074 ( .C1(n8278), .C2(n2836), .A(n2856), .B(n5991), .ZN(n1091)
         );
  OAI22_X1 U7075 ( .A1(n4730), .A2(n7599), .B1(n2825), .B2(n3775), .ZN(n5991)
         );
  INV_X1 U7076 ( .A(n4723), .ZN(n2836) );
  NAND2_X1 U7077 ( .A1(n1634), .A2(n1635), .ZN(n7943) );
  OAI221_X1 U7078 ( .B1(n1636), .B2(n3851), .C1(n7383), .C2(n1638), .A(n8291), 
        .ZN(n1635) );
  NAND3_X1 U7079 ( .A1(n4098), .A2(n4099), .A3(n4100), .ZN(n2446) );
  AND4_X1 U7080 ( .A1(n6897), .A2(n6894), .A3(n6882), .A4(n6692), .ZN(n4098)
         );
  NOR4_X1 U7081 ( .A1(n4101), .A2(n4102), .A3(n7412), .A4(n4123), .ZN(n4100)
         );
  AND3_X1 U7082 ( .A1(n4104), .A2(n6912), .A3(n6907), .ZN(n4099) );
  INV_X1 U7083 ( .A(n4305), .ZN(n1970) );
  OAI211_X1 U7084 ( .C1(n3730), .C2(n2506), .A(n4307), .B(n4308), .ZN(n4305)
         );
  NAND4_X1 U7085 ( .A1(n1576), .A2(n7433), .A3(n5063), .A4(n449), .ZN(n4307)
         );
  AOI22_X1 U7086 ( .A1(n2875), .A2(n7373), .B1(n1511), .B2(n2921), .ZN(n4308)
         );
  OR3_X1 U7087 ( .A1(n1947), .A2(n7393), .A3(n42), .ZN(n1486) );
  INV_X1 U7088 ( .A(n1727), .ZN(n2128) );
  AOI222_X1 U7089 ( .A1(n1728), .A2(n497), .B1(n1729), .B2(n1626), .C1(n4263), 
        .C2(n1533), .ZN(n1727) );
  OAI21_X1 U7090 ( .B1(n485), .B2(n1730), .A(n492), .ZN(n1729) );
  OR4_X1 U7091 ( .A1(n7399), .A2(n7476), .A3(n449), .A4(n1731), .ZN(n1728) );
  OAI22_X1 U7092 ( .A1(n7335), .A2(n2665), .B1(n3852), .B2(n3853), .ZN(Hvxhu6)
         );
  NAND4_X1 U7093 ( .A1(n6624), .A2(n6625), .A3(n7334), .A4(n7346), .ZN(n3853)
         );
  NAND4_X1 U7094 ( .A1(n7409), .A2(n7431), .A3(n3854), .A4(n7651), .ZN(n3852)
         );
  AND2_X1 U7095 ( .A1(n2665), .A2(n7652), .ZN(n3854) );
  AND2_X1 U7096 ( .A1(Jshpw6[8]), .A2(n421), .ZN(n430) );
  AND3_X1 U7097 ( .A1(n7653), .A2(n3479), .A3(n6915), .ZN(n4104) );
  AOI21_X1 U7098 ( .B1(n7305), .B2(n3982), .A(n7482), .ZN(Fwohu6) );
  OR2_X1 U7099 ( .A1(n535), .A2(n7293), .ZN(n3982) );
  OAI221_X1 U7100 ( .B1(n7306), .B2(n546), .C1(n3126), .C2(n548), .A(n549), 
        .ZN(n7834) );
  NAND3_X1 U7101 ( .A1(n1826), .A2(n551), .A3(n7306), .ZN(n549) );
  AOI21_X1 U7102 ( .B1(n552), .B2(n551), .A(n560), .ZN(n546) );
  INV_X1 U7103 ( .A(n553), .ZN(n3126) );
  OAI221_X1 U7104 ( .B1(n7293), .B2(n928), .C1(n7253), .C2(n913), .A(n1825), 
        .ZN(n7843) );
  INV_X1 U7105 ( .A(n673), .ZN(n1825) );
  OAI221_X1 U7106 ( .B1(n908), .B2(n7292), .C1(n3180), .C2(n7321), .A(n3190), 
        .ZN(n673) );
  OAI221_X1 U7107 ( .B1(n7337), .B2(n928), .C1(n7477), .C2(n913), .A(n3131), 
        .ZN(n8039) );
  INV_X1 U7108 ( .A(n2010), .ZN(n3131) );
  OAI221_X1 U7109 ( .B1(n908), .B2(n7640), .C1(n3180), .C2(n7336), .A(n3190), 
        .ZN(n2010) );
  OAI221_X1 U7110 ( .B1(n7253), .B2(n928), .C1(n7439), .C2(n913), .A(n3132), 
        .ZN(n7842) );
  INV_X1 U7111 ( .A(n668), .ZN(n3132) );
  OAI221_X1 U7112 ( .B1(n908), .B2(n7646), .C1(n3180), .C2(n6673), .A(n3190), 
        .ZN(n668) );
  AND3_X1 U7113 ( .A1(n3034), .A2(n3035), .A3(IRQ[13]), .ZN(Nothu6) );
  AOI221_X1 U7114 ( .B1(n3841), .B2(n6587), .C1(n762), .C2(n3986), .A(n233), 
        .ZN(n3034) );
  INV_X1 U7115 ( .A(n3038), .ZN(n3841) );
  AND3_X1 U7116 ( .A1(n2829), .A2(n2830), .A3(IRQ[25]), .ZN(Ppthu6) );
  AOI221_X1 U7117 ( .B1(n2831), .B2(n6589), .C1(n762), .C2(n3983), .A(n233), 
        .ZN(n2829) );
  AND3_X1 U7118 ( .A1(n2668), .A2(n2669), .A3(IRQ[10]), .ZN(Snthu6) );
  AOI221_X1 U7119 ( .B1(n3846), .B2(n6594), .C1(n762), .C2(n3939), .A(n233), 
        .ZN(n2668) );
  INV_X1 U7120 ( .A(n2672), .ZN(n3846) );
  AND3_X1 U7121 ( .A1(n2240), .A2(n2241), .A3(IRQ[11]), .ZN(Znthu6) );
  AOI221_X1 U7122 ( .B1(n3840), .B2(n6606), .C1(n762), .C2(n3959), .A(n233), 
        .ZN(n2240) );
  INV_X1 U7123 ( .A(n2245), .ZN(n3840) );
  INV_X1 U7124 ( .A(n5533), .ZN(n2901) );
  OAI22_X1 U7125 ( .A1(n6773), .A2(n2197), .B1(n7638), .B2(n2195), .ZN(n5533)
         );
  NAND2_X1 U7126 ( .A1(n571), .A2(n3137), .ZN(n7835) );
  INV_X1 U7127 ( .A(n573), .ZN(n3137) );
  OAI21_X1 U7128 ( .B1(n7420), .B2(n535), .A(n3242), .ZN(n571) );
  AOI211_X1 U7129 ( .C1(n574), .C2(n7312), .A(n244), .B(n7321), .ZN(n573) );
  NAND2_X1 U7130 ( .A1(n1972), .A2(n1973), .ZN(n8012) );
  OAI21_X1 U7131 ( .B1(n6885), .B2(n1963), .A(n8285), .ZN(n1973) );
  INV_X1 U7132 ( .A(n1605), .ZN(n3676) );
  AOI22_X1 U7133 ( .A1(n4572), .A2(n3682), .B1(n1607), .B2(n7393), .ZN(n1605)
         );
  INV_X1 U7134 ( .A(n4087), .ZN(n2616) );
  OAI22_X1 U7135 ( .A1(n4068), .A2(n6874), .B1(n2617), .B2(n6873), .ZN(n4087)
         );
  INV_X1 U7136 ( .A(n2011), .ZN(n3130) );
  AOI211_X1 U7137 ( .C1(n4042), .C2(n244), .A(n2013), .B(n2014), .ZN(n2011) );
  OAI22_X1 U7138 ( .A1(n908), .A2(n6649), .B1(n928), .B2(n7477), .ZN(n2013) );
  INV_X1 U7139 ( .A(n4067), .ZN(n2615) );
  OAI22_X1 U7140 ( .A1(n4068), .A2(n7452), .B1(n2617), .B2(n7453), .ZN(n4067)
         );
  OAI21_X1 U7141 ( .B1(n7482), .B2(n525), .A(n1819), .ZN(n7831) );
  AOI21_X1 U7142 ( .B1(n528), .B2(n4034), .A(n530), .ZN(n525) );
  INV_X1 U7143 ( .A(n527), .ZN(n1819) );
  NAND2_X1 U7144 ( .A1(n6661), .A2(n902), .ZN(n7880) );
  OR3_X1 U7145 ( .A1(n903), .A2(n904), .A3(n905), .ZN(n902) );
  INV_X1 U7146 ( .A(n2179), .ZN(n3139) );
  AOI22_X1 U7147 ( .A1(n2180), .A2(SWDITMS), .B1(n4022), .B2(n3140), .ZN(n2179) );
  INV_X1 U7148 ( .A(n2180), .ZN(n3140) );
  OAI211_X1 U7149 ( .C1(n2182), .C2(n4016), .A(n2183), .B(n7312), .ZN(n2180)
         );
  NOR3_X1 U7150 ( .A1(n4406), .A2(n7425), .A3(n1248), .ZN(n1075) );
  NOR2_X1 U7151 ( .A1(n1005), .A2(n7412), .ZN(n2137) );
  NOR2_X1 U7152 ( .A1(n984), .A2(n7412), .ZN(n2141) );
  NAND2_X1 U7153 ( .A1(n497), .A2(n7359), .ZN(n2864) );
  NOR4_X1 U7154 ( .A1(n7349), .A2(n7348), .A3(n7347), .A4(n7249), .ZN(n531) );
  NOR2_X1 U7155 ( .A1(n991), .A2(n7412), .ZN(n2108) );
  NOR2_X1 U7156 ( .A1(n2151), .A2(n7383), .ZN(n2106) );
  NOR3_X1 U7157 ( .A1(n3208), .A2(n7309), .A3(n2049), .ZN(n592) );
  NOR2_X1 U7158 ( .A1(n1008), .A2(n7412), .ZN(n118) );
  NOR3_X1 U7159 ( .A1(n6675), .A2(n6604), .A3(n4041), .ZN(n2157) );
  NOR2_X1 U7160 ( .A1(n7448), .A2(n7388), .ZN(n1344) );
  NOR2_X1 U7161 ( .A1(n113), .A2(n7412), .ZN(n2144) );
  NAND3_X1 U7162 ( .A1(n1344), .A2(n1183), .A3(n2854), .ZN(n1008) );
  NOR3_X1 U7163 ( .A1(n4405), .A2(n7425), .A3(n3913), .ZN(n2854) );
  NOR2_X1 U7164 ( .A1(n125), .A2(n7412), .ZN(n2192) );
  NOR2_X1 U7165 ( .A1(n1894), .A2(n7383), .ZN(n2112) );
  AOI21_X1 U7166 ( .B1(n3203), .B2(n4022), .A(n7312), .ZN(n636) );
  XNOR2_X1 U7167 ( .A(n7306), .B(n4022), .ZN(n2057) );
  NOR4_X1 U7168 ( .A1(n980), .A2(n981), .A3(n982), .A4(n983), .ZN(n979) );
  NAND3_X1 U7169 ( .A1(n993), .A2(n994), .A3(n3480), .ZN(n980) );
  OAI222_X1 U7170 ( .A1(n6856), .A2(n990), .B1(n6837), .B2(n991), .C1(n7457), 
        .C2(n992), .ZN(n981) );
  OAI222_X1 U7171 ( .A1(n4324), .A2(n987), .B1(n6803), .B2(n988), .C1(n7469), 
        .C2(n989), .ZN(n982) );
  NOR4_X1 U7172 ( .A1(n3696), .A2(Tzfpw6[7]), .A3(Tzfpw6[22]), .A4(Tzfpw6[2]), 
        .ZN(n3695) );
  NAND3_X1 U7173 ( .A1(n7692), .A2(n7699), .A3(n7687), .ZN(n3696) );
  AOI22_X1 U7174 ( .A1(n4022), .A2(n4011), .B1(SWDO), .B2(n570), .ZN(n552) );
  INV_X1 U7175 ( .A(n570), .ZN(n4011) );
  NOR2_X1 U7176 ( .A1(n913), .A2(n7318), .ZN(n570) );
  NOR4_X1 U7177 ( .A1(n7283), .A2(n7375), .A3(n2568), .A4(n4738), .ZN(n2892)
         );
  NOR2_X1 U7178 ( .A1(n7425), .A2(n7411), .ZN(n1290) );
  NOR2_X1 U7179 ( .A1(n4329), .A2(n7419), .ZN(n1346) );
  NOR4_X1 U7180 ( .A1(n590), .A2(n591), .A3(n592), .A4(n593), .ZN(n587) );
  OAI221_X1 U7181 ( .B1(n594), .B2(n595), .C1(n596), .C2(n597), .A(n598), .ZN(
        n590) );
  NOR2_X1 U7182 ( .A1(n596), .A2(n7306), .ZN(n594) );
  AND2_X1 U7183 ( .A1(n4032), .A2(n600), .ZN(n596) );
  NOR3_X1 U7184 ( .A1(n3226), .A2(n7308), .A3(n3208), .ZN(n593) );
  NOR3_X1 U7185 ( .A1(n7411), .A2(n7388), .A3(n3882), .ZN(n1304) );
  NOR3_X1 U7186 ( .A1(n3201), .A2(n7311), .A3(n3223), .ZN(n656) );
  NOR3_X1 U7187 ( .A1(n7314), .A2(n7310), .A3(n7315), .ZN(n662) );
  AOI221_X1 U7188 ( .B1(n3479), .B2(n1144), .C1(n3474), .C2(n4408), .A(n1146), 
        .ZN(n1142) );
  OAI22_X1 U7189 ( .A1(n7462), .A2(n984), .B1(n7455), .B2(n988), .ZN(n1146) );
  NOR3_X1 U7190 ( .A1(n3142), .A2(n7318), .A3(n3215), .ZN(n666) );
  NAND4_X1 U7191 ( .A1(n2045), .A2(n2046), .A3(n7318), .A4(n4028), .ZN(n604)
         );
  NOR3_X1 U7192 ( .A1(n4405), .A2(n7425), .A3(n4301), .ZN(n2132) );
  AOI221_X1 U7193 ( .B1(n7310), .B2(n7308), .C1(n610), .C2(n4024), .A(n648), 
        .ZN(n645) );
  NOR2_X1 U7194 ( .A1(n7518), .A2(n7510), .ZN(n2848) );
  NAND3_X1 U7195 ( .A1(n7425), .A2(n3913), .A3(n1344), .ZN(n1283) );
  OAI221_X1 U7196 ( .B1(n616), .B2(n3144), .C1(n7313), .C2(n555), .A(n618), 
        .ZN(n603) );
  AOI21_X1 U7197 ( .B1(n619), .B2(n7313), .A(n610), .ZN(n616) );
  OAI21_X1 U7198 ( .B1(n7318), .B2(n2056), .A(n4018), .ZN(n601) );
  AOI221_X1 U7199 ( .B1(n1333), .B2(n3479), .C1(n1290), .C2(n1334), .A(n1335), 
        .ZN(n1332) );
  NOR2_X1 U7200 ( .A1(n7414), .A2(n7440), .ZN(n1333) );
  OAI21_X1 U7201 ( .B1(n7448), .B2(n1337), .A(n1338), .ZN(n1334) );
  OAI22_X1 U7202 ( .A1(n6845), .A2(n990), .B1(n4054), .B2(n993), .ZN(n1335) );
  NOR2_X1 U7203 ( .A1(n7438), .A2(n7419), .ZN(n1310) );
  OAI222_X1 U7204 ( .A1(n7707), .A2(n984), .B1(n7471), .B2(n985), .C1(n6874), 
        .C2(n113), .ZN(n983) );
  OAI222_X1 U7205 ( .A1(n1004), .A2(n7475), .B1(n1005), .B2(n7708), .C1(n1006), 
        .C2(n7473), .ZN(n1003) );
  OAI222_X1 U7206 ( .A1(n6816), .A2(n989), .B1(n6799), .B2(n988), .C1(n6869), 
        .C2(n985), .ZN(n1016) );
  OAI222_X1 U7207 ( .A1(n1006), .A2(n6888), .B1(n984), .B2(n7465), .C1(n1005), 
        .C2(n7461), .ZN(n1280) );
  OAI222_X1 U7208 ( .A1(n1009), .A2(n7627), .B1(n113), .B2(n6873), .C1(n1005), 
        .C2(n7458), .ZN(n1147) );
  OAI222_X1 U7209 ( .A1(n6790), .A2(n988), .B1(n6843), .B2(n990), .C1(n6809), 
        .C2(n989), .ZN(n1097) );
  NOR2_X1 U7210 ( .A1(n2202), .A2(n7383), .ZN(n2103) );
  NAND3_X1 U7211 ( .A1(n7314), .A2(n4029), .A3(n610), .ZN(n618) );
  NOR2_X1 U7212 ( .A1(n1893), .A2(n7383), .ZN(n1886) );
  NAND3_X1 U7213 ( .A1(n2054), .A2(n7309), .A3(n7310), .ZN(n597) );
  INV_X1 U7214 ( .A(n2005), .ZN(n3009) );
  AOI211_X1 U7215 ( .C1(n236), .C2(n6644), .A(n542), .B(n2006), .ZN(n2005) );
  OAI22_X1 U7216 ( .A1(n537), .A2(n7439), .B1(n917), .B2(n7416), .ZN(n2006) );
  OAI22_X1 U7217 ( .A1(n7313), .A2(n598), .B1(n644), .B2(n4022), .ZN(n658) );
  NOR2_X1 U7218 ( .A1(n3686), .A2(n7259), .ZN(n3074) );
  OAI221_X1 U7219 ( .B1(n7519), .B2(n2256), .C1(n7525), .C2(n2572), .A(n4215), 
        .ZN(n2802) );
  NAND3_X1 U7220 ( .A1(n7388), .A2(n4405), .A3(n1291), .ZN(n1248) );
  NOR3_X1 U7221 ( .A1(n7448), .A2(n7411), .A3(n7438), .ZN(n1291) );
  NAND3_X1 U7222 ( .A1(n2054), .A2(n4028), .A3(n7310), .ZN(n595) );
  NOR3_X1 U7223 ( .A1(n4670), .A2(n7516), .A3(n4993), .ZN(n1743) );
  NAND2_X1 U7224 ( .A1(n474), .A2(n3234), .ZN(n2843) );
  OAI21_X1 U7225 ( .B1(n7329), .B2(n485), .A(n3709), .ZN(n3234) );
  NAND4_X1 U7226 ( .A1(n1290), .A2(n7448), .A3(n4405), .A4(n3470), .ZN(n987)
         );
  NOR2_X1 U7227 ( .A1(n2049), .A2(n7311), .ZN(n2045) );
  OAI21_X1 U7228 ( .B1(n6836), .B2(n2108), .A(n2134), .ZN(n7125) );
  NAND3_X1 U7229 ( .A1(n1371), .A2(n3388), .A3(n2108), .ZN(n2134) );
  OAI22_X1 U7230 ( .A1(n7451), .A2(n1345), .B1(n4405), .B2(n1275), .ZN(n1309)
         );
  NOR3_X1 U7231 ( .A1(n7533), .A2(n237), .A3(n7492), .ZN(n3720) );
  NAND3_X1 U7232 ( .A1(n1274), .A2(n7451), .A3(n1290), .ZN(n1247) );
  OAI211_X1 U7233 ( .C1(n1592), .C2(n4987), .A(n2918), .B(n2919), .ZN(n1756)
         );
  NOR2_X1 U7234 ( .A1(n7516), .A2(n7518), .ZN(n2919) );
  OAI21_X1 U7235 ( .B1(n7519), .B2(n7505), .A(n4987), .ZN(n2918) );
  NOR3_X1 U7236 ( .A1(n3528), .A2(n7519), .A3(n7523), .ZN(n3521) );
  OAI21_X1 U7237 ( .B1(n4993), .B2(n4978), .A(n7514), .ZN(n3528) );
  NAND3_X1 U7238 ( .A1(n7398), .A2(n4182), .A3(n2129), .ZN(n2127) );
  NAND2_X1 U7239 ( .A1(n7311), .A2(n7314), .ZN(n589) );
  OAI211_X1 U7240 ( .C1(n7318), .C2(n7319), .A(n4033), .B(n4032), .ZN(n626) );
  XNOR2_X1 U7241 ( .A(n7423), .B(Jshpw6[4]), .ZN(n948) );
  NAND2_X1 U7242 ( .A1(n1589), .A2(n7259), .ZN(n1731) );
  NAND2_X1 U7243 ( .A1(n1442), .A2(n5026), .ZN(n3029) );
  OAI211_X1 U7244 ( .C1(n5027), .C2(n2262), .A(n5028), .B(n2267), .ZN(n5026)
         );
  AOI22_X1 U7245 ( .A1(n7399), .A2(n4635), .B1(n7510), .B2(n7381), .ZN(n5027)
         );
  NAND3_X1 U7246 ( .A1(n5042), .A2(n2262), .A3(n2893), .ZN(n5028) );
  NAND3_X1 U7247 ( .A1(n7505), .A2(n4987), .A3(n7519), .ZN(n42) );
  NOR3_X1 U7248 ( .A1(n943), .A2(n152), .A3(n944), .ZN(n942) );
  OAI22_X1 U7249 ( .A1(n7447), .A2(n7450), .B1(n945), .B2(n4145), .ZN(n943) );
  OAI21_X1 U7250 ( .B1(n1990), .B2(n1991), .A(n2233), .ZN(\sub_3151/A[0] ) );
  NAND4_X1 U7251 ( .A1(n7501), .A2(n7502), .A3(n7503), .A4(n7504), .ZN(n1990)
         );
  NAND4_X1 U7252 ( .A1(n7496), .A2(n7498), .A3(n7499), .A4(n7500), .ZN(n1991)
         );
  OAI21_X1 U7253 ( .B1(n7519), .B2(n5042), .A(n7514), .ZN(n1602) );
  NAND3_X1 U7254 ( .A1(n7319), .A2(n4032), .A3(n7317), .ZN(n2056) );
  OAI22_X1 U7255 ( .A1(n1006), .A2(n6780), .B1(n1004), .B2(n6782), .ZN(n1065)
         );
  OAI22_X1 U7256 ( .A1(n1006), .A2(n6890), .B1(n1004), .B2(n6828), .ZN(n1230)
         );
  NOR2_X1 U7257 ( .A1(n4123), .A2(n6885), .ZN(n1391) );
  NOR2_X1 U7258 ( .A1(n4123), .A2(n6887), .ZN(n1379) );
  NAND2_X1 U7259 ( .A1(n7425), .A2(n1271), .ZN(n994) );
  OAI221_X1 U7260 ( .B1(n4406), .B2(n1248), .C1(n4324), .C2(n1272), .A(n1273), 
        .ZN(n1271) );
  NAND4_X1 U7261 ( .A1(n1274), .A2(n7451), .A3(n1275), .A4(n3913), .ZN(n1273)
         );
  AOI221_X1 U7262 ( .B1(n5040), .B2(n529), .C1(n5041), .C2(n1744), .A(n1511), 
        .ZN(n5039) );
  NOR2_X1 U7263 ( .A1(n7381), .A2(n475), .ZN(n5041) );
  OAI21_X1 U7264 ( .B1(n7519), .B2(n4187), .A(n4186), .ZN(n5040) );
  NOR3_X1 U7265 ( .A1(n3192), .A2(n7316), .A3(n624), .ZN(n621) );
  NOR3_X1 U7266 ( .A1(n4035), .A2(n7317), .A3(n7318), .ZN(n624) );
  NOR3_X1 U7267 ( .A1(n3202), .A2(n7314), .A3(n4016), .ZN(n2061) );
  INV_X1 U7268 ( .A(n1253), .ZN(n3450) );
  OAI22_X1 U7269 ( .A1(n1006), .A2(n6881), .B1(n1004), .B2(n6824), .ZN(n1253)
         );
  OAI221_X1 U7270 ( .B1(n6870), .B2(n985), .C1(n7694), .C2(n113), .A(n3451), 
        .ZN(n1177) );
  INV_X1 U7271 ( .A(n1189), .ZN(n3451) );
  OAI22_X1 U7272 ( .A1(n1006), .A2(n6895), .B1(n1004), .B2(n6833), .ZN(n1189)
         );
  OAI22_X1 U7273 ( .A1(n7318), .A2(n3141), .B1(n7319), .B2(n2184), .ZN(n7724)
         );
  OAI22_X1 U7274 ( .A1(n7313), .A2(n3141), .B1(n7316), .B2(n2184), .ZN(Yvohu6)
         );
  OAI22_X1 U7275 ( .A1(n7317), .A2(n3141), .B1(n7318), .B2(n2184), .ZN(n7725)
         );
  OAI22_X1 U7276 ( .A1(n7316), .A2(n3141), .B1(n7317), .B2(n2184), .ZN(Rvohu6)
         );
  NAND2_X1 U7277 ( .A1(n7310), .A2(n4029), .ZN(n2049) );
  NOR3_X1 U7278 ( .A1(n2186), .A2(n656), .A3(n2187), .ZN(n2182) );
  AOI211_X1 U7279 ( .C1(n7311), .C2(n2188), .A(n3212), .B(n3200), .ZN(n2187)
         );
  OAI22_X1 U7280 ( .A1(n7310), .A2(n3144), .B1(n3226), .B2(n4024), .ZN(n2186)
         );
  NAND2_X1 U7281 ( .A1(n7309), .A2(n7318), .ZN(n2188) );
  OAI221_X1 U7282 ( .B1(n2043), .B2(n3202), .C1(n2044), .C2(n548), .A(n604), 
        .ZN(n8053) );
  AOI21_X1 U7283 ( .B1(n3225), .B2(n4029), .A(n2048), .ZN(n2043) );
  NOR3_X1 U7285 ( .A1(n2047), .A2(n658), .A3(n657), .ZN(n2044) );
  OAI221_X1 U7286 ( .B1(n7313), .B2(n2050), .C1(n2049), .C2(n589), .A(n618), 
        .ZN(n2047) );
  NOR2_X1 U7287 ( .A1(n7285), .A2(n7503), .ZN(Vnfpw6[6]) );
  OAI22_X1 U7288 ( .A1(n6883), .A2(n1006), .B1(n6862), .B2(n985), .ZN(n1098)
         );
  OAI22_X1 U7289 ( .A1(n6693), .A2(n807), .B1(n6692), .B2(n2087), .ZN(n6924)
         );
  OAI22_X1 U7290 ( .A1(n6843), .A2(n807), .B1(n6882), .B2(n2087), .ZN(n7132)
         );
  OAI22_X1 U7291 ( .A1(n6844), .A2(n807), .B1(n6884), .B2(n2087), .ZN(n7133)
         );
  OAI22_X1 U7292 ( .A1(n6846), .A2(n807), .B1(n6885), .B2(n803), .ZN(n7136) );
  OAI22_X1 U7293 ( .A1(n6847), .A2(n807), .B1(n6887), .B2(n2087), .ZN(n7137)
         );
  OAI22_X1 U7295 ( .A1(n6848), .A2(n807), .B1(n6889), .B2(n2087), .ZN(n7138)
         );
  OAI22_X1 U7296 ( .A1(n6850), .A2(n807), .B1(n6908), .B2(n2087), .ZN(n7140)
         );
  OAI22_X1 U7297 ( .A1(n6851), .A2(n807), .B1(n6906), .B2(n2087), .ZN(n7141)
         );
  OAI22_X1 U7298 ( .A1(n6852), .A2(n807), .B1(n6903), .B2(n2087), .ZN(n7142)
         );
  OAI22_X1 U7299 ( .A1(n6853), .A2(n807), .B1(n6894), .B2(n2087), .ZN(n7143)
         );
  OAI22_X1 U7300 ( .A1(n6854), .A2(n807), .B1(n6915), .B2(n2087), .ZN(n7144)
         );
  OAI22_X1 U7301 ( .A1(n6855), .A2(n807), .B1(n6897), .B2(n2087), .ZN(n7145)
         );
  NAND3_X1 U7302 ( .A1(n7448), .A2(n4405), .A3(n1310), .ZN(n1338) );
  NOR2_X1 U7303 ( .A1(n7285), .A2(n7496), .ZN(Vnfpw6[0]) );
  NOR2_X1 U7304 ( .A1(n7285), .A2(n7501), .ZN(Vnfpw6[4]) );
  NOR2_X1 U7305 ( .A1(n7285), .A2(n7499), .ZN(Vnfpw6[2]) );
  OAI22_X1 U7306 ( .A1(n2953), .A2(n3547), .B1(n2954), .B2(n3548), .ZN(n2920)
         );
  AOI21_X1 U7307 ( .B1(n475), .B2(n4635), .A(n2262), .ZN(n2954) );
  NOR4_X1 U7308 ( .A1(n2956), .A2(n2957), .A3(n470), .A4(n4635), .ZN(n2953) );
  OAI22_X1 U7309 ( .A1(n4572), .A2(n4670), .B1(n7518), .B2(n4672), .ZN(n2957)
         );
  AOI21_X1 U7310 ( .B1(n7451), .B2(n7419), .A(n4306), .ZN(n1337) );
  OAI211_X1 U7311 ( .C1(n6653), .C2(n1000), .A(n2136), .B(n1180), .ZN(n1179)
         );
  XNOR2_X1 U7312 ( .A(n2585), .B(n7516), .ZN(n2956) );
  NAND2_X1 U7313 ( .A1(n3269), .A2(n7519), .ZN(n1494) );
  AOI22_X1 U7314 ( .A1(n2051), .A2(n2052), .B1(n619), .B2(n2053), .ZN(n2050)
         );
  NOR2_X1 U7315 ( .A1(n7316), .A2(n7317), .ZN(n2051) );
  OAI22_X1 U7316 ( .A1(n7318), .A2(n3192), .B1(n7306), .B2(n595), .ZN(n2052)
         );
  NOR2_X1 U7317 ( .A1(n7285), .A2(n7504), .ZN(Vnfpw6[7]) );
  OAI22_X1 U7318 ( .A1(n6837), .A2(n2108), .B1(n1832), .B2(n3419), .ZN(n7126)
         );
  OAI22_X1 U7319 ( .A1(n7452), .A2(n2192), .B1(n1832), .B2(n3471), .ZN(Z5xhu6)
         );
  OAI22_X1 U7320 ( .A1(n6874), .A2(n2144), .B1(n1832), .B2(n3473), .ZN(n7177)
         );
  OAI22_X1 U7321 ( .A1(n7457), .A2(n2147), .B1(n1832), .B2(n3444), .ZN(n7208)
         );
  INV_X1 U7322 ( .A(n2147), .ZN(n3444) );
  NOR2_X1 U7323 ( .A1(n992), .A2(n7412), .ZN(n2147) );
  OAI22_X1 U7324 ( .A1(n6831), .A2(n833), .B1(n6906), .B2(n828), .ZN(n7119) );
  OAI22_X1 U7325 ( .A1(n1397), .A2(n830), .B1(n6885), .B2(n828), .ZN(n7114) );
  OAI22_X1 U7326 ( .A1(n6827), .A2(n830), .B1(n6887), .B2(n828), .ZN(n7115) );
  OAI22_X1 U7327 ( .A1(n6728), .A2(n807), .B1(n6727), .B2(n803), .ZN(n6969) );
  OAI22_X1 U7328 ( .A1(n1832), .A2(n420), .B1(n6803), .B2(n818), .ZN(n7086) );
  OAI22_X1 U7329 ( .A1(n1832), .A2(n431), .B1(n6856), .B2(n807), .ZN(n7146) );
  OAI22_X1 U7330 ( .A1(n1832), .A2(n3460), .B1(n7708), .B2(n2137), .ZN(n7147)
         );
  OAI22_X1 U7331 ( .A1(n1832), .A2(n3454), .B1(n7707), .B2(n2141), .ZN(n7152)
         );
  OAI22_X1 U7332 ( .A1(n1832), .A2(n247), .B1(n7469), .B2(n841), .ZN(n7094) );
  OAI22_X1 U7333 ( .A1(n1832), .A2(n249), .B1(n7475), .B2(n830), .ZN(n7113) );
  OAI22_X1 U7334 ( .A1(n1832), .A2(n250), .B1(n7471), .B2(n857), .ZN(n7164) );
  OAI22_X1 U7335 ( .A1(n1832), .A2(n253), .B1(n7473), .B2(n850), .ZN(n7186) );
  AOI21_X1 U7336 ( .B1(n118), .B2(n119), .A(n7466), .ZN(n117) );
  OAI22_X1 U7337 ( .A1(n6689), .A2(n841), .B1(n6692), .B2(n2081), .ZN(n6921)
         );
  OAI22_X1 U7338 ( .A1(n6690), .A2(n830), .B1(n6692), .B2(n828), .ZN(n6922) );
  OAI22_X1 U7339 ( .A1(n6739), .A2(n833), .B1(n6741), .B2(n2083), .ZN(n6989)
         );
  OAI22_X1 U7340 ( .A1(n6742), .A2(n807), .B1(n6741), .B2(n803), .ZN(n6991) );
  OAI22_X1 U7341 ( .A1(n6723), .A2(n830), .B1(n6904), .B2(n2083), .ZN(n6965)
         );
  OAI22_X1 U7342 ( .A1(n6725), .A2(n807), .B1(n6904), .B2(n803), .ZN(n6967) );
  OAI22_X1 U7343 ( .A1(n6747), .A2(n833), .B1(n6750), .B2(n2083), .ZN(n6996)
         );
  OAI22_X1 U7344 ( .A1(n6749), .A2(n809), .B1(n6750), .B2(n803), .ZN(n6998) );
  OAI22_X1 U7345 ( .A1(n6715), .A2(n847), .B1(n6718), .B2(n2081), .ZN(n6958)
         );
  OAI22_X1 U7346 ( .A1(n6716), .A2(n833), .B1(n6718), .B2(n828), .ZN(n6959) );
  OAI22_X1 U7347 ( .A1(n6719), .A2(n807), .B1(n6718), .B2(n2087), .ZN(n6961)
         );
  OAI22_X1 U7348 ( .A1(n6823), .A2(n833), .B1(n6905), .B2(n2083), .ZN(n7109)
         );
  OAI22_X1 U7349 ( .A1(n6841), .A2(n809), .B1(n6905), .B2(n803), .ZN(n7130) );
  OAI22_X1 U7350 ( .A1(n6825), .A2(n830), .B1(n6882), .B2(n828), .ZN(n7111) );
  OAI22_X1 U7351 ( .A1(n6833), .A2(n830), .B1(n6894), .B2(n828), .ZN(n7121) );
  OAI22_X1 U7352 ( .A1(n7474), .A2(n830), .B1(n6897), .B2(n828), .ZN(n7123) );
  OAI22_X1 U7353 ( .A1(n6821), .A2(n833), .B1(n6907), .B2(n2083), .ZN(n7107)
         );
  OAI22_X1 U7354 ( .A1(n6839), .A2(n809), .B1(n6907), .B2(n803), .ZN(n7128) );
  OAI22_X1 U7355 ( .A1(n6732), .A2(n830), .B1(n6912), .B2(n2083), .ZN(n6973)
         );
  OAI22_X1 U7356 ( .A1(n6734), .A2(n809), .B1(n6912), .B2(n803), .ZN(n6975) );
  OAI22_X1 U7357 ( .A1(n6832), .A2(n830), .B1(n6903), .B2(n828), .ZN(n7120) );
  OAI22_X1 U7358 ( .A1(n6822), .A2(n833), .B1(n7653), .B2(n2083), .ZN(n7108)
         );
  OAI22_X1 U7359 ( .A1(n6840), .A2(n809), .B1(n7653), .B2(n803), .ZN(n7129) );
  OAI22_X1 U7360 ( .A1(n7484), .A2(n830), .B1(n6884), .B2(n2083), .ZN(n7112)
         );
  OAI22_X1 U7361 ( .A1(n6834), .A2(n830), .B1(n6915), .B2(n2083), .ZN(n7122)
         );
  OAI22_X1 U7362 ( .A1(n6696), .A2(n841), .B1(n6902), .B2(n2081), .ZN(n6927)
         );
  OAI22_X1 U7363 ( .A1(n6697), .A2(n830), .B1(n6902), .B2(n828), .ZN(n6928) );
  OAI22_X1 U7364 ( .A1(n6699), .A2(n809), .B1(n6902), .B2(n2087), .ZN(n6930)
         );
  OAI22_X1 U7365 ( .A1(n7456), .A2(n2144), .B1(n3012), .B2(n3473), .ZN(n7176)
         );
  OAI22_X1 U7366 ( .A1(n6824), .A2(n833), .B1(n6900), .B2(n828), .ZN(n7110) );
  OAI22_X1 U7367 ( .A1(n6828), .A2(n830), .B1(n6889), .B2(n828), .ZN(n7116) );
  OAI22_X1 U7368 ( .A1(n6842), .A2(n809), .B1(n6900), .B2(n803), .ZN(n7131) );
  OAI22_X1 U7369 ( .A1(n6820), .A2(n833), .B1(n6901), .B2(n2083), .ZN(n7106)
         );
  OAI22_X1 U7370 ( .A1(n6838), .A2(n809), .B1(n6901), .B2(n803), .ZN(n7127) );
  OAI22_X1 U7371 ( .A1(n6705), .A2(n841), .B1(n6708), .B2(n2081), .ZN(n6942)
         );
  OAI22_X1 U7372 ( .A1(n6706), .A2(n830), .B1(n6708), .B2(n828), .ZN(n6943) );
  OAI22_X1 U7373 ( .A1(n6709), .A2(n807), .B1(n6708), .B2(n2087), .ZN(n6945)
         );
  OAI22_X1 U7374 ( .A1(n6754), .A2(n833), .B1(n6756), .B2(n2083), .ZN(n7004)
         );
  OAI22_X1 U7375 ( .A1(n6757), .A2(n809), .B1(n6756), .B2(n803), .ZN(n7006) );
  OAI22_X1 U7376 ( .A1(n6764), .A2(n833), .B1(n6766), .B2(n2083), .ZN(n7019)
         );
  OAI22_X1 U7377 ( .A1(n6767), .A2(n809), .B1(n6766), .B2(n803), .ZN(n7021) );
  OAI22_X1 U7378 ( .A1(n6829), .A2(n830), .B1(n6875), .B2(n828), .ZN(n7117) );
  OAI22_X1 U7379 ( .A1(n6830), .A2(n830), .B1(n6908), .B2(n2083), .ZN(n7118)
         );
  OAI22_X1 U7380 ( .A1(n6849), .A2(n809), .B1(n6875), .B2(n2087), .ZN(n7139)
         );
  OAI22_X1 U7381 ( .A1(n6782), .A2(n833), .B1(n6911), .B2(n2083), .ZN(n7064)
         );
  OAI22_X1 U7382 ( .A1(n6784), .A2(n809), .B1(n6911), .B2(n803), .ZN(n7066) );
  NAND2_X1 U7383 ( .A1(n2045), .A2(n7309), .ZN(n557) );
  OAI221_X1 U7384 ( .B1(n1755), .B2(n475), .C1(n4572), .C2(n2262), .A(n2765), 
        .ZN(n2762) );
  AOI21_X1 U7385 ( .B1(n7381), .B2(n2766), .A(n2577), .ZN(n2765) );
  NAND2_X1 U7386 ( .A1(n7518), .A2(n1840), .ZN(n2766) );
  AND2_X1 U7387 ( .A1(n7319), .A2(n2178), .ZN(n528) );
  NAND3_X1 U7388 ( .A1(n4033), .A2(n4032), .A3(n4034), .ZN(n2178) );
  NOR2_X1 U7389 ( .A1(n1959), .A2(n6684), .ZN(n1960) );
  AOI21_X1 U7390 ( .B1(n643), .B2(n644), .A(n7313), .ZN(n638) );
  OAI22_X1 U7391 ( .A1(n7349), .A2(n4135), .B1(n7348), .B2(n2292), .ZN(Ytxhu6)
         );
  INV_X1 U7392 ( .A(n2292), .ZN(n4135) );
  NAND2_X1 U7393 ( .A1(n6675), .A2(n6604), .ZN(n2292) );
  NAND4_X1 U7394 ( .A1(n1904), .A2(n1905), .A3(n1906), .A4(n4685), .ZN(n1898)
         );
  OAI211_X1 U7395 ( .C1(n1909), .C2(n417), .A(n476), .B(n3549), .ZN(n1905) );
  OAI21_X1 U7396 ( .B1(n1912), .B2(n417), .A(n2124), .ZN(n1904) );
  OR4_X1 U7397 ( .A1(n1687), .A2(n4572), .A3(n4512), .A4(n7414), .ZN(n1906) );
  OAI22_X1 U7398 ( .A1(n6873), .A2(n2144), .B1(n3259), .B2(n3473), .ZN(n7175)
         );
  NOR2_X1 U7399 ( .A1(n8253), .A2(n7450), .ZN(n945) );
  OAI22_X1 U7400 ( .A1(n3012), .A2(n420), .B1(n6792), .B2(n818), .ZN(n7075) );
  OAI22_X1 U7401 ( .A1(n3012), .A2(n247), .B1(n1516), .B2(n841), .ZN(n7105) );
  OAI22_X1 U7402 ( .A1(n3012), .A2(n249), .B1(n1399), .B2(n830), .ZN(n7124) );
  OAI22_X1 U7403 ( .A1(n3012), .A2(n431), .B1(n6845), .B2(n807), .ZN(n7135) );
  OAI22_X1 U7404 ( .A1(n3012), .A2(n3460), .B1(n7459), .B2(n2137), .ZN(n7150)
         );
  OAI22_X1 U7405 ( .A1(n3012), .A2(n3454), .B1(n7463), .B2(n2141), .ZN(n7155)
         );
  OAI22_X1 U7406 ( .A1(n3012), .A2(n250), .B1(n1122), .B2(n857), .ZN(n7174) );
  OAI22_X1 U7407 ( .A1(n3012), .A2(n253), .B1(n1257), .B2(n850), .ZN(n7196) );
  OAI22_X1 U7408 ( .A1(n3012), .A2(n3471), .B1(n6643), .B2(n2192), .ZN(n7350)
         );
  OAI22_X1 U7409 ( .A1(n3259), .A2(n3471), .B1(n7453), .B2(n2192), .ZN(L5xhu6)
         );
  OAI22_X1 U7410 ( .A1(n3259), .A2(n3904), .B1(n7490), .B2(n2434), .ZN(Wexhu6)
         );
  OAI22_X1 U7411 ( .A1(n3259), .A2(n3460), .B1(n7458), .B2(n2137), .ZN(n7151)
         );
  OAI22_X1 U7412 ( .A1(n3259), .A2(n3454), .B1(n7462), .B2(n2141), .ZN(n7156)
         );
  OAI22_X1 U7413 ( .A1(n3259), .A2(n431), .B1(n7454), .B2(n807), .ZN(n7134) );
  OAI22_X1 U7414 ( .A1(n3259), .A2(n420), .B1(n7455), .B2(n818), .ZN(n7074) );
  OAI22_X1 U7415 ( .A1(n7461), .A2(n2137), .B1(n4117), .B2(n3460), .ZN(n7148)
         );
  OAI22_X1 U7416 ( .A1(n7460), .A2(n2137), .B1(n4052), .B2(n3460), .ZN(n7149)
         );
  OAI22_X1 U7417 ( .A1(n7465), .A2(n2141), .B1(n4117), .B2(n3454), .ZN(n7153)
         );
  OAI22_X1 U7418 ( .A1(n7464), .A2(n2141), .B1(n4052), .B2(n3454), .ZN(n7154)
         );
  OAI22_X1 U7419 ( .A1(n7347), .A2(n7348), .B1(n520), .B2(n1817), .ZN(n7829)
         );
  NOR2_X1 U7420 ( .A1(n4041), .A2(n4040), .ZN(n520) );
  OAI22_X1 U7421 ( .A1(n6913), .A2(n2149), .B1(n6914), .B2(n4115), .ZN(n7209)
         );
  OAI22_X1 U7422 ( .A1(n7489), .A2(n2434), .B1(n3904), .B2(n3469), .ZN(Kfxhu6)
         );
  NAND2_X1 U7423 ( .A1(n1407), .A2(n3259), .ZN(n3469) );
  OAI22_X1 U7424 ( .A1(n7421), .A2(n2434), .B1(n4117), .B2(n3904), .ZN(Dfxhu6)
         );
  AOI22_X1 U7425 ( .A1(n4219), .A2(n3181), .B1(n4635), .B2(n476), .ZN(n4218)
         );
  NOR2_X1 U7426 ( .A1(n7433), .A2(n7516), .ZN(n4219) );
  OR2_X1 U7427 ( .A1(n990), .A2(n7412), .ZN(n431) );
  OAI21_X1 U7428 ( .B1(n6743), .B2(n2108), .A(n2109), .ZN(n6992) );
  OR3_X1 U7429 ( .A1(n4123), .A2(n6750), .A3(n3419), .ZN(n2109) );
  NAND3_X1 U7430 ( .A1(n7290), .A2(n7339), .A3(n7288), .ZN(n3708) );
  NAND3_X1 U7431 ( .A1(n7537), .A2(n7539), .A3(n7445), .ZN(n3700) );
  NAND3_X1 U7432 ( .A1(n7369), .A2(n7391), .A3(n7368), .ZN(n3704) );
  AND3_X1 U7433 ( .A1(n7337), .A2(n7477), .A3(n7322), .ZN(n3772) );
  OR4_X1 U7435 ( .A1(n6727), .A2(n6718), .A3(n6741), .A4(n4103), .ZN(n4101) );
  OR2_X1 U7436 ( .A1(n6884), .A2(n6903), .ZN(n4103) );
  OAI21_X1 U7437 ( .B1(n6655), .B2(n1435), .A(n1436), .ZN(n7281) );
  NAND3_X1 U7438 ( .A1(n604), .A2(n3156), .A3(n2038), .ZN(n8052) );
  AOI22_X1 U7439 ( .A1(n2039), .A2(n609), .B1(n4015), .B2(n2040), .ZN(n2038)
         );
  XNOR2_X1 U7440 ( .A(n648), .B(n7311), .ZN(n2039) );
  OAI211_X1 U7441 ( .C1(n597), .C2(n601), .A(n3219), .B(n3195), .ZN(n2040) );
  OR3_X1 U7442 ( .A1(n6905), .A2(n6904), .A3(n6906), .ZN(n4102) );
  OR3_X1 U7443 ( .A1(n4028), .A2(n7308), .A3(n589), .ZN(n588) );
  INV_X1 U7444 ( .A(n2042), .ZN(n3195) );
  OAI222_X1 U7445 ( .A1(n4022), .A2(n643), .B1(n3223), .B2(n589), .C1(n618), 
        .C2(n7311), .ZN(n2042) );
  INV_X1 U7446 ( .A(n1191), .ZN(n3468) );
  OAI22_X1 U7447 ( .A1(n988), .A2(n6800), .B1(n989), .B2(n6817), .ZN(n1191) );
  OR2_X1 U7448 ( .A1(n7285), .A2(n7498), .ZN(n432) );
  OR2_X1 U7449 ( .A1(n7285), .A2(n7502), .ZN(n436) );
  OR2_X1 U7450 ( .A1(n7285), .A2(n7500), .ZN(n437) );
  INV_X1 U7451 ( .A(n1315), .ZN(n3456) );
  OAI21_X1 U7452 ( .B1(n984), .B2(n7464), .A(n1316), .ZN(n1315) );
  OR3_X1 U7453 ( .A1(n1283), .A2(n4405), .A3(n4324), .ZN(n1316) );
  INV_X1 U7454 ( .A(n1341), .ZN(n3472) );
  OAI22_X1 U7455 ( .A1(n6643), .A2(n125), .B1(n7466), .B2(n1008), .ZN(n1341)
         );
  INV_X1 U7456 ( .A(n1292), .ZN(n3467) );
  OAI22_X1 U7457 ( .A1(n989), .A2(n6811), .B1(n985), .B2(n6864), .ZN(n1292) );
  OR2_X1 U7458 ( .A1(n717), .A2(n718), .ZN(n7853) );
  AOI21_X1 U7459 ( .B1(n118), .B2(n710), .A(n7467), .ZN(n718) );
  NOR3_X4 U7460 ( .A1(n2964), .A2(n7332), .A3(n5786), .ZN(n4705) );
  NOR3_X4 U7461 ( .A1(n5786), .A2(n7332), .A3(n1342), .ZN(n4691) );
  INV_X1 U7462 ( .A(n4154), .ZN(n438) );
  INV_X1 U7463 ( .A(n438), .ZN(n439) );
  NOR3_X4 U7464 ( .A1(n3858), .A2(n7279), .A3(n1528), .ZN(n4424) );
  NOR3_X4 U7465 ( .A1(n386), .A2(n3394), .A3(n5712), .ZN(n2239) );
  NOR3_X4 U7466 ( .A1(n100), .A2(n3416), .A3(n5106), .ZN(n2321) );
  NOR3_X4 U7467 ( .A1(n402), .A2(n3425), .A3(n4613), .ZN(n2399) );
  NOR3_X4 U7468 ( .A1(n3410), .A2(n2150), .A3(n302), .ZN(n2209) );
  NOR3_X4 U7469 ( .A1(n3440), .A2(n2150), .A3(n276), .ZN(n2271) );
  AOI211_X4 U7470 ( .C1(n479), .C2(n4749), .A(n1851), .B(n483), .ZN(n241) );
  BUF_X1 U7471 ( .A(n7373), .Z(n502) );
  INV_X1 U7472 ( .A(n7355), .ZN(n516) );
  BUF_X1 U7473 ( .A(n523), .Z(n522) );
  BUF_X1 U7474 ( .A(n7282), .Z(n536) );
  INV_X1 U7475 ( .A(n387), .ZN(n568) );
  INV_X1 U7476 ( .A(n4763), .ZN(n631) );
  BUF_X1 U7477 ( .A(n660), .Z(n659) );
  INV_X1 U7478 ( .A(n242), .ZN(n667) );
  INV_X1 U7479 ( .A(n242), .ZN(n669) );
  BUF_X1 U7480 ( .A(n2611), .Z(n678) );
  BUF_X1 U7481 ( .A(n2362), .Z(n681) );
  BUF_X1 U7482 ( .A(n683), .Z(n682) );
  INV_X1 U7483 ( .A(n681), .ZN(n683) );
  BUF_X1 U7484 ( .A(n686), .Z(n685) );
  INV_X1 U7485 ( .A(n2348), .ZN(n686) );
  BUF_X1 U7486 ( .A(n2344), .Z(n687) );
  BUF_X1 U7487 ( .A(n690), .Z(n688) );
  INV_X1 U7488 ( .A(n687), .ZN(n690) );
  BUF_X1 U7489 ( .A(n695), .Z(n694) );
  INV_X1 U7490 ( .A(n2315), .ZN(n695) );
  BUF_X1 U7491 ( .A(n701), .Z(n697) );
  INV_X1 U7492 ( .A(n2297), .ZN(n701) );
  BUF_X1 U7493 ( .A(n2289), .Z(n704) );
  BUF_X1 U7494 ( .A(n709), .Z(n706) );
  INV_X1 U7495 ( .A(n704), .ZN(n709) );
  BUF_X1 U7496 ( .A(n2285), .Z(n712) );
  BUF_X1 U7497 ( .A(n714), .Z(n713) );
  INV_X1 U7498 ( .A(n712), .ZN(n714) );
  BUF_X1 U7499 ( .A(n736), .Z(n734) );
  INV_X1 U7500 ( .A(n2264), .ZN(n736) );
  BUF_X1 U7501 ( .A(n739), .Z(n738) );
  INV_X1 U7502 ( .A(n2253), .ZN(n739) );
  BUF_X1 U7503 ( .A(n2249), .Z(n740) );
  BUF_X1 U7504 ( .A(n744), .Z(n743) );
  INV_X1 U7505 ( .A(n740), .ZN(n744) );
  BUF_X1 U7506 ( .A(n2237), .Z(n747) );
  BUF_X1 U7507 ( .A(n749), .Z(n748) );
  INV_X1 U7508 ( .A(n747), .ZN(n749) );
  BUF_X1 U7509 ( .A(n2231), .Z(n751) );
  BUF_X1 U7510 ( .A(n755), .Z(n753) );
  INV_X1 U7511 ( .A(n751), .ZN(n755) );
  BUF_X1 U7512 ( .A(n761), .Z(n760) );
  INV_X1 U7513 ( .A(n2229), .ZN(n761) );
  BUF_X1 U7514 ( .A(n768), .Z(n767) );
  INV_X1 U7515 ( .A(n2218), .ZN(n768) );
  BUF_X1 U7516 ( .A(n2214), .Z(n771) );
  BUF_X1 U7517 ( .A(n775), .Z(n772) );
  INV_X1 U7518 ( .A(n771), .ZN(n775) );
  BUF_X1 U7519 ( .A(n780), .Z(n779) );
  INV_X1 U7520 ( .A(n2210), .ZN(n780) );
  INV_X1 U7521 ( .A(n431), .ZN(n807) );
  INV_X1 U7522 ( .A(n420), .ZN(n818) );
  INV_X1 U7523 ( .A(n741), .ZN(n883) );
  INV_X1 U7524 ( .A(n719), .ZN(n890) );
  INV_X1 U7525 ( .A(N701), .ZN(n963) );
  NOR2_X1 U7526 ( .A1(Vnfpw6[0]), .A2(\sub_3151/A[0] ), .ZN(n972) );
  AOI21_X1 U7527 ( .B1(\sub_3151/A[0] ), .B2(Vnfpw6[0]), .A(n972), .ZN(n964)
         );
  INV_X1 U7528 ( .A(n964), .ZN(Xlfpw6[1]) );
  NAND2_X1 U7529 ( .A1(n972), .A2(n432), .ZN(n974) );
  OAI21_X1 U7530 ( .B1(n972), .B2(n432), .A(n974), .ZN(Xlfpw6[2]) );
  NOR2_X1 U7531 ( .A1(n974), .A2(Vnfpw6[2]), .ZN(n976) );
  AOI21_X1 U7532 ( .B1(n974), .B2(Vnfpw6[2]), .A(n976), .ZN(n975) );
  INV_X1 U7533 ( .A(n975), .ZN(Xlfpw6[3]) );
  NAND2_X1 U7534 ( .A1(n976), .A2(n437), .ZN(n977) );
  OAI21_X1 U7535 ( .B1(n976), .B2(n437), .A(n977), .ZN(Xlfpw6[4]) );
  NOR2_X1 U7536 ( .A1(n977), .A2(Vnfpw6[4]), .ZN(n995) );
  AOI21_X1 U7537 ( .B1(n977), .B2(Vnfpw6[4]), .A(n995), .ZN(n986) );
  INV_X1 U7538 ( .A(n986), .ZN(Xlfpw6[5]) );
  NAND2_X1 U7539 ( .A1(n995), .A2(n436), .ZN(n1001) );
  OAI21_X1 U7540 ( .B1(n995), .B2(n436), .A(n1001), .ZN(Xlfpw6[6]) );
  XNOR2_X1 U7541 ( .A(Vnfpw6[6]), .B(n1001), .ZN(Xlfpw6[7]) );
  NOR2_X1 U7542 ( .A1(Vnfpw6[6]), .A2(n1001), .ZN(n1010) );
  XOR2_X1 U7543 ( .A(Vnfpw6[7]), .B(n1010), .Z(Xlfpw6[8]) );
  MUX2_X1 U7544 ( .A(Oodhu6), .B(PORESETn), .S(N427), .Z(Fmdhu6) );
  XNOR2_X1 U7545 ( .A(Togpw6[24]), .B(\eq_3147/A[22] ), .ZN(n1019) );
  XNOR2_X1 U7546 ( .A(Togpw6[23]), .B(\eq_3147/A[21] ), .ZN(n1014) );
  XNOR2_X1 U7547 ( .A(Togpw6[25]), .B(\eq_3147/A[23] ), .ZN(n1013) );
  NAND3_X1 U7548 ( .A1(n1019), .A2(n1014), .A3(n1013), .ZN(n1033) );
  XOR2_X1 U7549 ( .A(Togpw6[28]), .B(\eq_3147/A[26] ), .Z(n1031) );
  XOR2_X1 U7550 ( .A(Togpw6[26]), .B(\eq_3147/A[24] ), .Z(n1025) );
  XOR2_X1 U7551 ( .A(Togpw6[27]), .B(\eq_3147/A[25] ), .Z(n1024) );
  NOR4_X1 U7552 ( .A1(n1033), .A2(n1031), .A3(n1025), .A4(n1024), .ZN(n1117)
         );
  XNOR2_X1 U7553 ( .A(Togpw6[19]), .B(\eq_3147/A[17] ), .ZN(n1046) );
  XNOR2_X1 U7554 ( .A(Togpw6[18]), .B(\eq_3147/A[16] ), .ZN(n1041) );
  XNOR2_X1 U7555 ( .A(Togpw6[17]), .B(\eq_3147/A[15] ), .ZN(n1040) );
  XNOR2_X1 U7556 ( .A(Togpw6[16]), .B(\eq_3147/A[14] ), .ZN(n1038) );
  NAND4_X1 U7557 ( .A1(n1046), .A2(n1041), .A3(n1040), .A4(n1038), .ZN(n1060)
         );
  XOR2_X1 U7558 ( .A(Togpw6[22]), .B(\eq_3147/A[20] ), .Z(n1057) );
  XOR2_X1 U7559 ( .A(Togpw6[20]), .B(\eq_3147/A[18] ), .Z(n1049) );
  XOR2_X1 U7560 ( .A(Togpw6[21]), .B(\eq_3147/A[19] ), .Z(n1048) );
  NOR4_X1 U7561 ( .A1(n1060), .A2(n1057), .A3(n1049), .A4(n1048), .ZN(n1115)
         );
  XNOR2_X1 U7562 ( .A(Togpw6[12]), .B(\eq_3147/A[10] ), .ZN(n1068) );
  XNOR2_X1 U7563 ( .A(Togpw6[11]), .B(\eq_3147/A[9] ), .ZN(n1067) );
  XNOR2_X1 U7564 ( .A(Togpw6[10]), .B(\eq_3147/A[8] ), .ZN(n1063) );
  XNOR2_X1 U7565 ( .A(Togpw6[9]), .B(\eq_3147/A[7] ), .ZN(n1061) );
  NAND4_X1 U7566 ( .A1(n1068), .A2(n1067), .A3(n1063), .A4(n1061), .ZN(n1081)
         );
  XOR2_X1 U7567 ( .A(Togpw6[15]), .B(\eq_3147/A[13] ), .Z(n1078) );
  XOR2_X1 U7568 ( .A(Togpw6[13]), .B(\eq_3147/A[11] ), .Z(n1072) );
  XOR2_X1 U7569 ( .A(Togpw6[14]), .B(\eq_3147/A[12] ), .Z(n1071) );
  NOR4_X1 U7570 ( .A1(n1081), .A2(n1078), .A3(n1072), .A4(n1071), .ZN(n1114)
         );
  XNOR2_X1 U7571 ( .A(Togpw6[5]), .B(\eq_3147/A[3] ), .ZN(n1099) );
  XNOR2_X1 U7572 ( .A(Togpw6[4]), .B(\eq_3147/A[2] ), .ZN(n1096) );
  NOR2_X1 U7573 ( .A1(n1122), .A2(\eq_3147/A[0] ), .ZN(n1084) );
  OAI22_X1 U7574 ( .A1(n1084), .A2(n1798), .B1(Togpw6[3]), .B2(n1084), .ZN(
        n1095) );
  AND2_X1 U7575 ( .A1(\eq_3147/A[0] ), .A2(n1122), .ZN(n1088) );
  OAI22_X1 U7576 ( .A1(\eq_3147/A[1] ), .A2(n1088), .B1(n1088), .B2(n1119), 
        .ZN(n1092) );
  NAND4_X1 U7577 ( .A1(n1099), .A2(n1096), .A3(n1095), .A4(n1092), .ZN(n1112)
         );
  XOR2_X1 U7578 ( .A(Togpw6[8]), .B(\eq_3147/A[6] ), .Z(n1105) );
  XOR2_X1 U7579 ( .A(Togpw6[6]), .B(\eq_3147/A[4] ), .Z(n1103) );
  XOR2_X1 U7580 ( .A(Togpw6[7]), .B(\eq_3147/A[5] ), .Z(n1100) );
  NOR4_X1 U7581 ( .A1(n1112), .A2(n1105), .A3(n1103), .A4(n1100), .ZN(n1113)
         );
  XNOR2_X1 U7582 ( .A(Gqgpw6[24]), .B(\eq_3147/A[22] ), .ZN(n1130) );
  XNOR2_X1 U7583 ( .A(Gqgpw6[23]), .B(\eq_3147/A[21] ), .ZN(n1128) );
  XNOR2_X1 U7584 ( .A(Gqgpw6[25]), .B(\eq_3147/A[23] ), .ZN(n1126) );
  NAND3_X1 U7585 ( .A1(n1130), .A2(n1128), .A3(n1126), .ZN(n1141) );
  XOR2_X1 U7586 ( .A(Gqgpw6[28]), .B(\eq_3147/A[26] ), .Z(n1138) );
  XOR2_X1 U7587 ( .A(Gqgpw6[26]), .B(\eq_3147/A[24] ), .Z(n1134) );
  XOR2_X1 U7588 ( .A(Gqgpw6[27]), .B(\eq_3147/A[25] ), .Z(n1132) );
  NOR4_X1 U7589 ( .A1(n1141), .A2(n1138), .A3(n1134), .A4(n1132), .ZN(n1254)
         );
  XNOR2_X1 U7590 ( .A(Gqgpw6[19]), .B(\eq_3147/A[17] ), .ZN(n1155) );
  XNOR2_X1 U7591 ( .A(Gqgpw6[18]), .B(\eq_3147/A[16] ), .ZN(n1150) );
  XNOR2_X1 U7592 ( .A(Gqgpw6[17]), .B(\eq_3147/A[15] ), .ZN(n1145) );
  XNOR2_X1 U7593 ( .A(Gqgpw6[16]), .B(\eq_3147/A[14] ), .ZN(n1143) );
  NAND4_X1 U7594 ( .A1(n1155), .A2(n1150), .A3(n1145), .A4(n1143), .ZN(n1163)
         );
  XOR2_X1 U7595 ( .A(Gqgpw6[22]), .B(\eq_3147/A[20] ), .Z(n1161) );
  XOR2_X1 U7596 ( .A(Gqgpw6[20]), .B(\eq_3147/A[18] ), .Z(n1159) );
  XOR2_X1 U7597 ( .A(Gqgpw6[21]), .B(\eq_3147/A[19] ), .Z(n1157) );
  NOR4_X1 U7598 ( .A1(n1163), .A2(n1161), .A3(n1159), .A4(n1157), .ZN(n1252)
         );
  XNOR2_X1 U7599 ( .A(Gqgpw6[12]), .B(\eq_3147/A[10] ), .ZN(n1184) );
  XNOR2_X1 U7600 ( .A(Gqgpw6[11]), .B(\eq_3147/A[9] ), .ZN(n1175) );
  XNOR2_X1 U7601 ( .A(Gqgpw6[10]), .B(\eq_3147/A[8] ), .ZN(n1170) );
  XNOR2_X1 U7602 ( .A(Gqgpw6[9]), .B(\eq_3147/A[7] ), .ZN(n1168) );
  NAND4_X1 U7603 ( .A1(n1184), .A2(n1175), .A3(n1170), .A4(n1168), .ZN(n1190)
         );
  XOR2_X1 U7604 ( .A(Gqgpw6[15]), .B(\eq_3147/A[13] ), .Z(n1188) );
  XOR2_X1 U7605 ( .A(Gqgpw6[13]), .B(\eq_3147/A[11] ), .Z(n1187) );
  XOR2_X1 U7606 ( .A(Gqgpw6[14]), .B(\eq_3147/A[12] ), .Z(n1185) );
  NOR4_X1 U7607 ( .A1(n1190), .A2(n1188), .A3(n1187), .A4(n1185), .ZN(n1250)
         );
  XNOR2_X1 U7608 ( .A(Gqgpw6[5]), .B(\eq_3147/A[3] ), .ZN(n1221) );
  XNOR2_X1 U7609 ( .A(Gqgpw6[4]), .B(\eq_3147/A[2] ), .ZN(n1212) );
  NOR2_X1 U7610 ( .A1(n1257), .A2(\eq_3147/A[0] ), .ZN(n1197) );
  OAI22_X1 U7611 ( .A1(n1197), .A2(n1798), .B1(Gqgpw6[3]), .B2(n1197), .ZN(
        n1210) );
  AND2_X1 U7612 ( .A1(\eq_3147/A[0] ), .A2(n1257), .ZN(n1198) );
  OAI22_X1 U7613 ( .A1(\eq_3147/A[1] ), .A2(n1198), .B1(n1198), .B2(n1256), 
        .ZN(n1205) );
  NAND4_X1 U7614 ( .A1(n1221), .A2(n1212), .A3(n1210), .A4(n1205), .ZN(n1236)
         );
  XOR2_X1 U7615 ( .A(Gqgpw6[8]), .B(\eq_3147/A[6] ), .Z(n1233) );
  XOR2_X1 U7616 ( .A(Gqgpw6[6]), .B(\eq_3147/A[4] ), .Z(n1231) );
  XOR2_X1 U7617 ( .A(Gqgpw6[7]), .B(\eq_3147/A[5] ), .Z(n1226) );
  NOR4_X1 U7618 ( .A1(n1236), .A2(n1233), .A3(n1231), .A4(n1226), .ZN(n1243)
         );
  XNOR2_X1 U7619 ( .A(Trgpw6[24]), .B(\eq_3147/A[22] ), .ZN(n1268) );
  XNOR2_X1 U7620 ( .A(Trgpw6[23]), .B(\eq_3147/A[21] ), .ZN(n1261) );
  XNOR2_X1 U7621 ( .A(Trgpw6[25]), .B(\eq_3147/A[23] ), .ZN(n1259) );
  NAND3_X1 U7622 ( .A1(n1268), .A2(n1261), .A3(n1259), .ZN(n1286) );
  XOR2_X1 U7623 ( .A(Trgpw6[28]), .B(\eq_3147/A[26] ), .Z(n1285) );
  XOR2_X1 U7624 ( .A(Trgpw6[26]), .B(\eq_3147/A[24] ), .Z(n1279) );
  XOR2_X1 U7625 ( .A(Trgpw6[27]), .B(\eq_3147/A[25] ), .Z(n1276) );
  NOR4_X1 U7626 ( .A1(n1286), .A2(n1285), .A3(n1279), .A4(n1276), .ZN(n1395)
         );
  XNOR2_X1 U7627 ( .A(Trgpw6[19]), .B(\eq_3147/A[17] ), .ZN(n1306) );
  XNOR2_X1 U7628 ( .A(Trgpw6[18]), .B(\eq_3147/A[16] ), .ZN(n1305) );
  XNOR2_X1 U7629 ( .A(Trgpw6[17]), .B(\eq_3147/A[15] ), .ZN(n1289) );
  XNOR2_X1 U7630 ( .A(Trgpw6[16]), .B(\eq_3147/A[14] ), .ZN(n1288) );
  NAND4_X1 U7631 ( .A1(n1306), .A2(n1305), .A3(n1289), .A4(n1288), .ZN(n1314)
         );
  XOR2_X1 U7632 ( .A(Trgpw6[22]), .B(\eq_3147/A[20] ), .Z(n1312) );
  XOR2_X1 U7633 ( .A(Trgpw6[20]), .B(\eq_3147/A[18] ), .Z(n1308) );
  XOR2_X1 U7634 ( .A(Trgpw6[21]), .B(\eq_3147/A[19] ), .Z(n1307) );
  NOR4_X1 U7635 ( .A1(n1314), .A2(n1312), .A3(n1308), .A4(n1307), .ZN(n1393)
         );
  XNOR2_X1 U7636 ( .A(Trgpw6[12]), .B(\eq_3147/A[10] ), .ZN(n1331) );
  XNOR2_X1 U7637 ( .A(Trgpw6[11]), .B(\eq_3147/A[9] ), .ZN(n1326) );
  XNOR2_X1 U7638 ( .A(Trgpw6[10]), .B(\eq_3147/A[8] ), .ZN(n1322) );
  XNOR2_X1 U7639 ( .A(Trgpw6[9]), .B(\eq_3147/A[7] ), .ZN(n1317) );
  NAND4_X1 U7640 ( .A1(n1331), .A2(n1326), .A3(n1322), .A4(n1317), .ZN(n1349)
         );
  XOR2_X1 U7641 ( .A(Trgpw6[15]), .B(\eq_3147/A[13] ), .Z(n1340) );
  XOR2_X1 U7642 ( .A(Trgpw6[13]), .B(\eq_3147/A[11] ), .Z(n1339) );
  XOR2_X1 U7643 ( .A(Trgpw6[14]), .B(\eq_3147/A[12] ), .Z(n1336) );
  NOR4_X1 U7644 ( .A1(n1349), .A2(n1340), .A3(n1339), .A4(n1336), .ZN(n1388)
         );
  XNOR2_X1 U7645 ( .A(Trgpw6[5]), .B(\eq_3147/A[3] ), .ZN(n1375) );
  XNOR2_X1 U7646 ( .A(Trgpw6[4]), .B(\eq_3147/A[2] ), .ZN(n1372) );
  NOR2_X1 U7647 ( .A1(n1399), .A2(\eq_3147/A[0] ), .ZN(n1350) );
  OAI22_X1 U7648 ( .A1(n1350), .A2(n1798), .B1(Trgpw6[3]), .B2(n1350), .ZN(
        n1370) );
  AND2_X1 U7649 ( .A1(\eq_3147/A[0] ), .A2(n1399), .ZN(n1367) );
  OAI22_X1 U7650 ( .A1(\eq_3147/A[1] ), .A2(n1367), .B1(n1367), .B2(n1397), 
        .ZN(n1368) );
  NAND4_X1 U7651 ( .A1(n1375), .A2(n1372), .A3(n1370), .A4(n1368), .ZN(n1384)
         );
  XOR2_X1 U7652 ( .A(Trgpw6[8]), .B(\eq_3147/A[6] ), .Z(n1382) );
  XOR2_X1 U7653 ( .A(Trgpw6[6]), .B(\eq_3147/A[4] ), .Z(n1381) );
  XOR2_X1 U7654 ( .A(Trgpw6[7]), .B(\eq_3147/A[5] ), .Z(n1380) );
  NOR4_X1 U7655 ( .A1(n1384), .A2(n1382), .A3(n1381), .A4(n1380), .ZN(n1386)
         );
  XNOR2_X1 U7656 ( .A(Gtgpw6[24]), .B(\eq_3147/A[22] ), .ZN(n1405) );
  XNOR2_X1 U7657 ( .A(Gtgpw6[23]), .B(\eq_3147/A[21] ), .ZN(n1402) );
  XNOR2_X1 U7658 ( .A(Gtgpw6[25]), .B(\eq_3147/A[23] ), .ZN(n1401) );
  NAND3_X1 U7659 ( .A1(n1405), .A2(n1402), .A3(n1401), .ZN(n1416) );
  XOR2_X1 U7660 ( .A(Gtgpw6[28]), .B(\eq_3147/A[26] ), .Z(n1415) );
  XOR2_X1 U7661 ( .A(Gtgpw6[26]), .B(\eq_3147/A[24] ), .Z(n1409) );
  XOR2_X1 U7662 ( .A(Gtgpw6[27]), .B(\eq_3147/A[25] ), .Z(n1406) );
  NOR4_X1 U7663 ( .A1(n1416), .A2(n1415), .A3(n1409), .A4(n1406), .ZN(n1514)
         );
  XNOR2_X1 U7664 ( .A(Gtgpw6[19]), .B(\eq_3147/A[17] ), .ZN(n1427) );
  XNOR2_X1 U7665 ( .A(Gtgpw6[18]), .B(\eq_3147/A[16] ), .ZN(n1423) );
  XNOR2_X1 U7666 ( .A(Gtgpw6[17]), .B(\eq_3147/A[15] ), .ZN(n1421) );
  XNOR2_X1 U7667 ( .A(Gtgpw6[16]), .B(\eq_3147/A[14] ), .ZN(n1420) );
  NAND4_X1 U7668 ( .A1(n1427), .A2(n1423), .A3(n1421), .A4(n1420), .ZN(n1446)
         );
  XOR2_X1 U7669 ( .A(Gtgpw6[22]), .B(\eq_3147/A[20] ), .Z(n1434) );
  XOR2_X1 U7670 ( .A(Gtgpw6[20]), .B(\eq_3147/A[18] ), .Z(n1432) );
  XOR2_X1 U7671 ( .A(Gtgpw6[21]), .B(\eq_3147/A[19] ), .Z(n1429) );
  NOR4_X1 U7672 ( .A1(n1446), .A2(n1434), .A3(n1432), .A4(n1429), .ZN(n1510)
         );
  XNOR2_X1 U7673 ( .A(Gtgpw6[12]), .B(\eq_3147/A[10] ), .ZN(n1450) );
  XNOR2_X1 U7674 ( .A(Gtgpw6[11]), .B(\eq_3147/A[9] ), .ZN(n1449) );
  XNOR2_X1 U7675 ( .A(Gtgpw6[10]), .B(\eq_3147/A[8] ), .ZN(n1448) );
  XNOR2_X1 U7676 ( .A(Gtgpw6[9]), .B(\eq_3147/A[7] ), .ZN(n1447) );
  NAND4_X1 U7677 ( .A1(n1450), .A2(n1449), .A3(n1448), .A4(n1447), .ZN(n1472)
         );
  XOR2_X1 U7678 ( .A(Gtgpw6[15]), .B(\eq_3147/A[13] ), .Z(n1469) );
  XOR2_X1 U7679 ( .A(Gtgpw6[13]), .B(\eq_3147/A[11] ), .Z(n1467) );
  XOR2_X1 U7680 ( .A(Gtgpw6[14]), .B(\eq_3147/A[12] ), .Z(n1460) );
  NOR4_X1 U7681 ( .A1(n1472), .A2(n1469), .A3(n1467), .A4(n1460), .ZN(n1509)
         );
  XNOR2_X1 U7682 ( .A(Gtgpw6[5]), .B(\eq_3147/A[3] ), .ZN(n1491) );
  XNOR2_X1 U7683 ( .A(Gtgpw6[4]), .B(\eq_3147/A[2] ), .ZN(n1490) );
  NOR2_X1 U7684 ( .A1(n1516), .A2(\eq_3147/A[0] ), .ZN(n1476) );
  OAI22_X1 U7685 ( .A1(n1476), .A2(n1798), .B1(Gtgpw6[3]), .B2(n1476), .ZN(
        n1485) );
  AND2_X1 U7686 ( .A1(\eq_3147/A[0] ), .A2(n1516), .ZN(n1481) );
  OAI22_X1 U7687 ( .A1(\eq_3147/A[1] ), .A2(n1481), .B1(n1481), .B2(n1515), 
        .ZN(n1484) );
  NAND4_X1 U7688 ( .A1(n1491), .A2(n1490), .A3(n1485), .A4(n1484), .ZN(n1507)
         );
  XOR2_X1 U7689 ( .A(Gtgpw6[8]), .B(\eq_3147/A[6] ), .Z(n1506) );
  XOR2_X1 U7690 ( .A(Gtgpw6[6]), .B(\eq_3147/A[4] ), .Z(n1500) );
  XOR2_X1 U7691 ( .A(Gtgpw6[7]), .B(\eq_3147/A[5] ), .Z(n1492) );
  NOR4_X1 U7692 ( .A1(n1507), .A2(n1506), .A3(n1500), .A4(n1492), .ZN(n1508)
         );
endmodule


module CORTEXM0INTEGRATION ( FCLK, SCLK, HCLK, DCLK, PORESETn, DBGRESETn, 
        HRESETn, SWCLKTCK, nTRST, HADDR, HBURST, HMASTLOCK, HPROT, HSIZE, 
        HTRANS, HWDATA, HWRITE, HRDATA, HREADY, HRESP, HMASTER, CODENSEQ, 
        CODEHINTDE, SPECHTRANS, SWDITMS, TDI, SWDO, SWDOEN, TDO, nTDOEN, 
        DBGRESTART, DBGRESTARTED, EDBGRQ, HALTED, NMI, IRQ, TXEV, RXEV, LOCKUP, 
        SYSRESETREQ, STCALIB, STCLKEN, IRQLATENCY, ECOREVNUM, GATEHCLK, 
        SLEEPING, SLEEPDEEP, WAKEUP, WICSENSE, SLEEPHOLDREQn, SLEEPHOLDACKn, 
        WICENREQ, WICENACK, CDBGPWRUPREQ, CDBGPWRUPACK, SE, RSTBYPASS );
  output [31:0] HADDR;
  output [2:0] HBURST;
  output [3:0] HPROT;
  output [2:0] HSIZE;
  output [1:0] HTRANS;
  output [31:0] HWDATA;
  input [31:0] HRDATA;
  output [2:0] CODEHINTDE;
  input [31:0] IRQ;
  input [25:0] STCALIB;
  input [7:0] IRQLATENCY;
  input [27:0] ECOREVNUM;
  output [33:0] WICSENSE;
  input FCLK, SCLK, HCLK, DCLK, PORESETn, DBGRESETn, HRESETn, SWCLKTCK, nTRST,
         HREADY, HRESP, SWDITMS, TDI, DBGRESTART, EDBGRQ, NMI, RXEV, STCLKEN,
         SLEEPHOLDREQn, WICENREQ, CDBGPWRUPACK, SE, RSTBYPASS;
  output HMASTLOCK, HWRITE, HMASTER, CODENSEQ, SPECHTRANS, SWDO, SWDOEN, TDO,
         nTDOEN, DBGRESTARTED, HALTED, TXEV, LOCKUP, SYSRESETREQ, GATEHCLK,
         SLEEPING, SLEEPDEEP, WAKEUP, SLEEPHOLDACKn, WICENACK, CDBGPWRUPREQ;

  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2;

  cortexm0ds_logic u_logic ( .FCLK(FCLK), .SCLK(SCLK), .HCLK(HCLK), .DCLK(DCLK), .PORESETn(PORESETn), .DBGRESETn(DBGRESETn), .HRESETn(HRESETn), .SWCLKTCK(
        SWCLKTCK), .nTRST(nTRST), .HADDR(HADDR), .HPROT({HPROT[3:2], 
        SYNOPSYS_UNCONNECTED__0, HPROT[0]}), .HSIZE({SYNOPSYS_UNCONNECTED__1, 
        HSIZE[1:0]}), .HTRANS({HTRANS[1], SYNOPSYS_UNCONNECTED__2}), .HWDATA(
        HWDATA), .HWRITE(HWRITE), .HRDATA(HRDATA), .HREADY(HREADY), .HRESP(
        HRESP), .HMASTER(HMASTER), .CODENSEQ(CODENSEQ), .CODEHINTDE(CODEHINTDE), .SPECHTRANS(SPECHTRANS), .SWDITMS(SWDITMS), .TDI(TDI), .SWDO(SWDO), .SWDOEN(
        SWDOEN), .DBGRESTART(DBGRESTART), .DBGRESTARTED(DBGRESTARTED), 
        .EDBGRQ(EDBGRQ), .HALTED(HALTED), .NMI(NMI), .IRQ(IRQ), .TXEV(TXEV), 
        .RXEV(RXEV), .LOCKUP(LOCKUP), .SYSRESETREQ(SYSRESETREQ), .STCALIB(
        STCALIB), .STCLKEN(STCLKEN), .IRQLATENCY(IRQLATENCY), .ECOREVNUM(
        ECOREVNUM), .GATEHCLK(GATEHCLK), .SLEEPING(SLEEPING), .SLEEPDEEP(
        SLEEPDEEP), .SLEEPHOLDREQn(SLEEPHOLDREQn), .SLEEPHOLDACKn(
        SLEEPHOLDACKn), .WICENREQ(WICENREQ), .CDBGPWRUPREQ(CDBGPWRUPREQ), 
        .CDBGPWRUPACK(CDBGPWRUPACK), .SE(SE), .RSTBYPASS(RSTBYPASS) );
  INV_X1 U1 ( .A(1'b1), .ZN(WICENACK) );
  INV_X1 U3 ( .A(1'b1), .ZN(WICSENSE[0]) );
  INV_X1 U5 ( .A(1'b1), .ZN(WICSENSE[1]) );
  INV_X1 U7 ( .A(1'b1), .ZN(WICSENSE[2]) );
  INV_X1 U9 ( .A(1'b1), .ZN(WICSENSE[3]) );
  INV_X1 U11 ( .A(1'b1), .ZN(WICSENSE[4]) );
  INV_X1 U13 ( .A(1'b1), .ZN(WICSENSE[5]) );
  INV_X1 U15 ( .A(1'b1), .ZN(WICSENSE[6]) );
  INV_X1 U17 ( .A(1'b1), .ZN(WICSENSE[7]) );
  INV_X1 U19 ( .A(1'b1), .ZN(WICSENSE[8]) );
  INV_X1 U21 ( .A(1'b1), .ZN(WICSENSE[9]) );
  INV_X1 U23 ( .A(1'b1), .ZN(WICSENSE[10]) );
  INV_X1 U25 ( .A(1'b1), .ZN(WICSENSE[11]) );
  INV_X1 U27 ( .A(1'b1), .ZN(WICSENSE[12]) );
  INV_X1 U29 ( .A(1'b1), .ZN(WICSENSE[13]) );
  INV_X1 U31 ( .A(1'b1), .ZN(WICSENSE[14]) );
  INV_X1 U33 ( .A(1'b1), .ZN(WICSENSE[15]) );
  INV_X1 U35 ( .A(1'b1), .ZN(WICSENSE[16]) );
  INV_X1 U37 ( .A(1'b1), .ZN(WICSENSE[17]) );
  INV_X1 U39 ( .A(1'b1), .ZN(WICSENSE[18]) );
  INV_X1 U41 ( .A(1'b1), .ZN(WICSENSE[19]) );
  INV_X1 U43 ( .A(1'b1), .ZN(WICSENSE[20]) );
  INV_X1 U45 ( .A(1'b1), .ZN(WICSENSE[21]) );
  INV_X1 U47 ( .A(1'b1), .ZN(WICSENSE[22]) );
  INV_X1 U49 ( .A(1'b1), .ZN(WICSENSE[23]) );
  INV_X1 U51 ( .A(1'b1), .ZN(WICSENSE[24]) );
  INV_X1 U53 ( .A(1'b1), .ZN(WICSENSE[25]) );
  INV_X1 U55 ( .A(1'b1), .ZN(WICSENSE[26]) );
  INV_X1 U57 ( .A(1'b1), .ZN(WICSENSE[27]) );
  INV_X1 U59 ( .A(1'b1), .ZN(WICSENSE[28]) );
  INV_X1 U61 ( .A(1'b1), .ZN(WICSENSE[29]) );
  INV_X1 U63 ( .A(1'b1), .ZN(WICSENSE[30]) );
  INV_X1 U65 ( .A(1'b1), .ZN(WICSENSE[31]) );
  INV_X1 U67 ( .A(1'b1), .ZN(WICSENSE[32]) );
  INV_X1 U69 ( .A(1'b1), .ZN(WICSENSE[33]) );
  INV_X1 U71 ( .A(1'b1), .ZN(WAKEUP) );
  INV_X1 U73 ( .A(1'b1), .ZN(nTDOEN) );
  INV_X1 U75 ( .A(1'b1), .ZN(TDO) );
  INV_X1 U77 ( .A(1'b1), .ZN(HTRANS[0]) );
  INV_X1 U79 ( .A(1'b1), .ZN(HSIZE[2]) );
  INV_X1 U81 ( .A(1'b0), .ZN(HPROT[1]) );
  INV_X1 U83 ( .A(1'b1), .ZN(HMASTLOCK) );
  INV_X1 U85 ( .A(1'b1), .ZN(HBURST[0]) );
  INV_X1 U87 ( .A(1'b1), .ZN(HBURST[1]) );
  INV_X1 U89 ( .A(1'b1), .ZN(HBURST[2]) );
endmodule

